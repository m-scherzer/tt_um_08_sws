MACRO digital_top
  CLASS BLOCK ;
  FOREIGN digital_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 124.280 BY 135.000 ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 114.520 10.640 116.520 122.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 84.520 10.640 86.520 122.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.520 10.640 56.520 122.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 24.520 10.640 26.520 122.640 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 99.520 10.640 101.520 122.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 69.520 10.640 71.520 122.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 39.520 10.640 41.520 122.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.520 10.640 11.520 122.640 ;
    END
  END VPWR
  PIN i_dem_dis
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 2.000 116.240 ;
    END
  END i_dem_dis
  PIN i_reset
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 2.000 50.960 ;
    END
  END i_reset
  PIN i_sys_clk
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 2.000 83.600 ;
    END
  END i_sys_clk
  PIN o_cs_cell_hi[0]
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 5.150 133.000 5.430 135.000 ;
    END
  END o_cs_cell_hi[0]
  PIN o_cs_cell_hi[1]
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 11.130 133.000 11.410 135.000 ;
    END
  END o_cs_cell_hi[1]
  PIN o_cs_cell_hi[2]
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 17.110 133.000 17.390 135.000 ;
    END
  END o_cs_cell_hi[2]
  PIN o_cs_cell_hi[3]
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 23.090 133.000 23.370 135.000 ;
    END
  END o_cs_cell_hi[3]
  PIN o_cs_cell_hi[4]
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 29.070 133.000 29.350 135.000 ;
    END
  END o_cs_cell_hi[4]
  PIN o_cs_cell_hi[5]
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 35.050 133.000 35.330 135.000 ;
    END
  END o_cs_cell_hi[5]
  PIN o_cs_cell_hi[6]
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 41.030 133.000 41.310 135.000 ;
    END
  END o_cs_cell_hi[6]
  PIN o_cs_cell_hi[7]
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 47.010 133.000 47.290 135.000 ;
    END
  END o_cs_cell_hi[7]
  PIN o_cs_cell_hi[8]
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 52.990 133.000 53.270 135.000 ;
    END
  END o_cs_cell_hi[8]
  PIN o_cs_cell_hi[9]
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 58.970 133.000 59.250 135.000 ;
    END
  END o_cs_cell_hi[9]
  PIN o_cs_cell_lo[0]
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 64.950 133.000 65.230 135.000 ;
    END
  END o_cs_cell_lo[0]
  PIN o_cs_cell_lo[1]
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 70.930 133.000 71.210 135.000 ;
    END
  END o_cs_cell_lo[1]
  PIN o_cs_cell_lo[2]
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 76.910 133.000 77.190 135.000 ;
    END
  END o_cs_cell_lo[2]
  PIN o_cs_cell_lo[3]
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 82.890 133.000 83.170 135.000 ;
    END
  END o_cs_cell_lo[3]
  PIN o_cs_cell_lo[4]
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 88.870 133.000 89.150 135.000 ;
    END
  END o_cs_cell_lo[4]
  PIN o_cs_cell_lo[5]
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 94.850 133.000 95.130 135.000 ;
    END
  END o_cs_cell_lo[5]
  PIN o_cs_cell_lo[6]
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 100.830 133.000 101.110 135.000 ;
    END
  END o_cs_cell_lo[6]
  PIN o_cs_cell_lo[7]
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 106.810 133.000 107.090 135.000 ;
    END
  END o_cs_cell_lo[7]
  PIN o_cs_cell_lo[8]
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 112.790 133.000 113.070 135.000 ;
    END
  END o_cs_cell_lo[8]
  PIN o_cs_cell_lo[9]
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 118.770 133.000 119.050 135.000 ;
    END
  END o_cs_cell_lo[9]
  OBS
      LAYER nwell ;
        RECT 5.330 120.985 118.870 122.590 ;
      LAYER pwell ;
        RECT 5.525 119.785 6.895 120.595 ;
        RECT 6.905 119.785 12.415 120.595 ;
        RECT 12.435 119.785 13.785 120.695 ;
        RECT 13.805 119.785 17.475 120.595 ;
        RECT 18.415 119.870 18.845 120.655 ;
        RECT 18.865 119.785 24.375 120.595 ;
        RECT 24.385 119.785 29.895 120.595 ;
        RECT 29.905 119.785 31.275 120.595 ;
        RECT 31.295 119.870 31.725 120.655 ;
        RECT 36.255 120.465 37.185 120.685 ;
        RECT 39.905 120.465 42.115 120.695 ;
        RECT 31.745 119.785 42.115 120.465 ;
        RECT 42.325 119.785 44.155 120.595 ;
        RECT 44.175 119.870 44.605 120.655 ;
        RECT 44.625 119.785 50.135 120.595 ;
        RECT 50.145 119.785 55.655 120.595 ;
        RECT 55.665 119.785 57.035 120.595 ;
        RECT 57.055 119.870 57.485 120.655 ;
        RECT 57.505 119.785 63.015 120.595 ;
        RECT 63.025 119.785 68.535 120.595 ;
        RECT 68.545 119.785 69.915 120.595 ;
        RECT 69.935 119.870 70.365 120.655 ;
        RECT 70.385 119.785 75.895 120.595 ;
        RECT 75.905 119.785 81.415 120.595 ;
        RECT 81.425 119.785 82.795 120.595 ;
        RECT 82.815 119.870 83.245 120.655 ;
        RECT 83.265 119.785 88.775 120.595 ;
        RECT 88.785 119.785 94.295 120.595 ;
        RECT 94.305 119.785 95.675 120.595 ;
        RECT 95.695 119.870 96.125 120.655 ;
        RECT 96.145 119.785 97.975 120.595 ;
        RECT 102.495 120.465 103.425 120.685 ;
        RECT 106.145 120.465 108.355 120.695 ;
        RECT 97.985 119.785 108.355 120.465 ;
        RECT 108.575 119.870 109.005 120.655 ;
        RECT 109.025 119.785 114.535 120.595 ;
        RECT 114.545 119.785 117.295 120.595 ;
        RECT 117.305 119.785 118.675 120.595 ;
        RECT 5.665 119.575 5.835 119.785 ;
        RECT 7.045 119.765 7.215 119.785 ;
        RECT 7.045 119.595 7.225 119.765 ;
        RECT 7.055 119.575 7.225 119.595 ;
        RECT 8.425 119.575 8.595 119.765 ;
        RECT 13.485 119.595 13.655 119.785 ;
        RECT 13.945 119.595 14.115 119.785 ;
        RECT 17.635 119.630 17.795 119.740 ;
        RECT 19.005 119.595 19.175 119.785 ;
        RECT 20.385 119.575 20.555 119.765 ;
        RECT 20.845 119.575 21.015 119.765 ;
        RECT 24.525 119.595 24.695 119.785 ;
        RECT 30.045 119.595 30.215 119.785 ;
        RECT 31.885 119.575 32.055 119.785 ;
        RECT 35.560 119.625 35.680 119.735 ;
        RECT 36.025 119.575 36.195 119.765 ;
        RECT 42.465 119.595 42.635 119.785 ;
        RECT 44.765 119.595 44.935 119.785 ;
        RECT 46.605 119.575 46.775 119.765 ;
        RECT 50.285 119.595 50.455 119.785 ;
        RECT 55.805 119.595 55.975 119.785 ;
        RECT 57.645 119.575 57.815 119.785 ;
        RECT 59.485 119.575 59.655 119.765 ;
        RECT 63.165 119.595 63.335 119.785 ;
        RECT 68.685 119.595 68.855 119.785 ;
        RECT 70.065 119.575 70.235 119.765 ;
        RECT 70.525 119.595 70.695 119.785 ;
        RECT 76.045 119.595 76.215 119.785 ;
        RECT 80.645 119.575 80.815 119.765 ;
        RECT 81.565 119.595 81.735 119.785 ;
        RECT 82.035 119.620 82.195 119.730 ;
        RECT 83.405 119.575 83.575 119.785 ;
        RECT 88.925 119.595 89.095 119.785 ;
        RECT 94.445 119.595 94.615 119.785 ;
        RECT 96.285 119.595 96.455 119.785 ;
        RECT 98.125 119.595 98.295 119.785 ;
        RECT 104.105 119.575 104.275 119.765 ;
        RECT 105.485 119.575 105.655 119.765 ;
        RECT 105.945 119.575 106.115 119.765 ;
        RECT 109.165 119.575 109.335 119.785 ;
        RECT 114.685 119.575 114.855 119.785 ;
        RECT 118.365 119.575 118.535 119.785 ;
        RECT 5.525 118.765 6.895 119.575 ;
        RECT 6.905 118.795 8.275 119.575 ;
        RECT 8.285 118.765 10.115 119.575 ;
        RECT 10.325 118.895 20.695 119.575 ;
        RECT 20.705 118.895 31.075 119.575 ;
        RECT 10.325 118.665 12.535 118.895 ;
        RECT 15.255 118.675 16.185 118.895 ;
        RECT 25.215 118.675 26.145 118.895 ;
        RECT 28.865 118.665 31.075 118.895 ;
        RECT 31.295 118.705 31.725 119.490 ;
        RECT 31.745 118.765 35.415 119.575 ;
        RECT 35.885 118.895 46.255 119.575 ;
        RECT 46.465 118.895 56.835 119.575 ;
        RECT 40.395 118.675 41.325 118.895 ;
        RECT 44.045 118.665 46.255 118.895 ;
        RECT 50.975 118.675 51.905 118.895 ;
        RECT 54.625 118.665 56.835 118.895 ;
        RECT 57.055 118.705 57.485 119.490 ;
        RECT 57.505 118.765 59.335 119.575 ;
        RECT 59.345 118.895 69.715 119.575 ;
        RECT 69.925 118.895 80.295 119.575 ;
        RECT 63.855 118.675 64.785 118.895 ;
        RECT 67.505 118.665 69.715 118.895 ;
        RECT 74.435 118.675 75.365 118.895 ;
        RECT 78.085 118.665 80.295 118.895 ;
        RECT 80.515 118.665 81.865 119.575 ;
        RECT 82.815 118.705 83.245 119.490 ;
        RECT 83.265 118.895 93.635 119.575 ;
        RECT 87.775 118.675 88.705 118.895 ;
        RECT 91.425 118.665 93.635 118.895 ;
        RECT 94.045 118.895 104.415 119.575 ;
        RECT 94.045 118.665 96.255 118.895 ;
        RECT 98.975 118.675 99.905 118.895 ;
        RECT 104.435 118.665 105.785 119.575 ;
        RECT 105.805 118.765 108.555 119.575 ;
        RECT 108.575 118.705 109.005 119.490 ;
        RECT 109.025 118.765 114.535 119.575 ;
        RECT 114.545 118.765 117.295 119.575 ;
        RECT 117.305 118.765 118.675 119.575 ;
      LAYER nwell ;
        RECT 5.330 115.545 118.870 118.375 ;
      LAYER pwell ;
        RECT 5.525 114.345 6.895 115.155 ;
        RECT 7.105 115.025 9.315 115.255 ;
        RECT 12.035 115.025 12.965 115.245 ;
        RECT 7.105 114.345 17.475 115.025 ;
        RECT 18.415 114.430 18.845 115.215 ;
        RECT 23.375 115.025 24.305 115.245 ;
        RECT 27.025 115.025 29.235 115.255 ;
        RECT 18.865 114.345 29.235 115.025 ;
        RECT 29.455 114.345 30.805 115.255 ;
        RECT 30.825 114.345 32.195 115.155 ;
        RECT 32.215 114.345 33.565 115.255 ;
        RECT 38.095 115.025 39.025 115.245 ;
        RECT 41.745 115.025 43.955 115.255 ;
        RECT 33.585 114.345 43.955 115.025 ;
        RECT 44.175 114.430 44.605 115.215 ;
        RECT 44.625 114.345 45.995 115.125 ;
        RECT 50.975 115.025 51.905 115.245 ;
        RECT 54.625 115.025 56.835 115.255 ;
        RECT 46.465 114.345 56.835 115.025 ;
        RECT 57.045 114.345 58.415 115.125 ;
        RECT 63.855 115.025 64.785 115.245 ;
        RECT 67.505 115.025 69.715 115.255 ;
        RECT 59.345 114.345 69.715 115.025 ;
        RECT 69.935 114.430 70.365 115.215 ;
        RECT 70.385 114.345 71.755 115.125 ;
        RECT 71.775 114.345 73.125 115.255 ;
        RECT 73.145 114.345 74.515 115.155 ;
        RECT 74.535 114.345 75.885 115.255 ;
        RECT 80.415 115.025 81.345 115.245 ;
        RECT 84.065 115.025 86.275 115.255 ;
        RECT 75.905 114.345 86.275 115.025 ;
        RECT 86.485 114.345 87.855 115.125 ;
        RECT 87.875 114.345 89.225 115.255 ;
        RECT 89.705 114.345 91.075 115.125 ;
        RECT 91.085 114.345 92.455 115.155 ;
        RECT 92.475 114.345 93.825 115.255 ;
        RECT 94.305 114.345 95.675 115.125 ;
        RECT 95.695 114.430 96.125 115.215 ;
        RECT 100.655 115.025 101.585 115.245 ;
        RECT 104.305 115.025 106.515 115.255 ;
        RECT 111.235 115.025 112.165 115.245 ;
        RECT 114.885 115.025 117.095 115.255 ;
        RECT 96.145 114.345 106.515 115.025 ;
        RECT 106.725 114.345 117.095 115.025 ;
        RECT 117.305 114.345 118.675 115.155 ;
        RECT 5.665 114.135 5.835 114.345 ;
        RECT 17.165 114.135 17.335 114.345 ;
        RECT 17.635 114.190 17.795 114.300 ;
        RECT 18.545 114.135 18.715 114.325 ;
        RECT 19.005 114.135 19.175 114.345 ;
        RECT 21.305 114.135 21.475 114.325 ;
        RECT 22.685 114.135 22.855 114.325 ;
        RECT 23.145 114.135 23.315 114.325 ;
        RECT 24.525 114.135 24.695 114.325 ;
        RECT 26.825 114.135 26.995 114.325 ;
        RECT 27.285 114.135 27.455 114.325 ;
        RECT 30.505 114.155 30.675 114.345 ;
        RECT 30.965 114.295 31.135 114.345 ;
        RECT 30.960 114.185 31.135 114.295 ;
        RECT 30.965 114.155 31.135 114.185 ;
        RECT 31.885 114.135 32.055 114.325 ;
        RECT 32.345 114.155 32.515 114.345 ;
        RECT 33.265 114.135 33.435 114.325 ;
        RECT 33.725 114.155 33.895 114.345 ;
        RECT 36.945 114.135 37.115 114.325 ;
        RECT 39.245 114.135 39.415 114.325 ;
        RECT 40.625 114.135 40.795 114.325 ;
        RECT 41.085 114.135 41.255 114.325 ;
        RECT 45.685 114.135 45.855 114.345 ;
        RECT 46.145 114.295 46.315 114.325 ;
        RECT 46.140 114.185 46.315 114.295 ;
        RECT 46.145 114.135 46.315 114.185 ;
        RECT 46.605 114.155 46.775 114.345 ;
        RECT 48.900 114.185 49.020 114.295 ;
        RECT 50.285 114.135 50.455 114.325 ;
        RECT 53.040 114.135 53.210 114.325 ;
        RECT 53.515 114.180 53.675 114.290 ;
        RECT 54.425 114.135 54.595 114.325 ;
        RECT 55.805 114.135 55.975 114.325 ;
        RECT 57.645 114.135 57.815 114.325 ;
        RECT 58.105 114.155 58.275 114.345 ;
        RECT 58.575 114.190 58.735 114.300 ;
        RECT 59.485 114.155 59.655 114.345 ;
        RECT 63.160 114.185 63.280 114.295 ;
        RECT 64.545 114.135 64.715 114.325 ;
        RECT 65.005 114.135 65.175 114.325 ;
        RECT 66.840 114.185 66.960 114.295 ;
        RECT 68.225 114.135 68.395 114.325 ;
        RECT 68.685 114.135 68.855 114.325 ;
        RECT 70.520 114.185 70.640 114.295 ;
        RECT 71.445 114.155 71.615 114.345 ;
        RECT 72.825 114.155 72.995 114.345 ;
        RECT 73.285 114.325 73.455 114.345 ;
        RECT 73.280 114.155 73.455 114.325 ;
        RECT 73.280 114.135 73.450 114.155 ;
        RECT 73.745 114.135 73.915 114.325 ;
        RECT 74.665 114.155 74.835 114.345 ;
        RECT 76.045 114.135 76.215 114.345 ;
        RECT 76.505 114.135 76.675 114.325 ;
        RECT 80.195 114.180 80.355 114.290 ;
        RECT 82.025 114.135 82.195 114.325 ;
        RECT 82.480 114.185 82.600 114.295 ;
        RECT 83.405 114.135 83.575 114.325 ;
        RECT 87.545 114.155 87.715 114.345 ;
        RECT 88.005 114.155 88.175 114.345 ;
        RECT 88.925 114.135 89.095 114.325 ;
        RECT 89.380 114.185 89.500 114.295 ;
        RECT 89.845 114.155 90.015 114.345 ;
        RECT 91.225 114.155 91.395 114.345 ;
        RECT 92.605 114.155 92.775 114.345 ;
        RECT 93.980 114.185 94.100 114.295 ;
        RECT 94.445 114.135 94.615 114.345 ;
        RECT 96.285 114.155 96.455 114.345 ;
        RECT 97.200 114.185 97.320 114.295 ;
        RECT 97.665 114.135 97.835 114.325 ;
        RECT 99.055 114.180 99.215 114.290 ;
        RECT 99.965 114.135 100.135 114.325 ;
        RECT 101.345 114.135 101.515 114.325 ;
        RECT 102.725 114.135 102.895 114.325 ;
        RECT 104.565 114.135 104.735 114.325 ;
        RECT 105.945 114.135 106.115 114.325 ;
        RECT 106.865 114.155 107.035 114.345 ;
        RECT 109.165 114.135 109.335 114.325 ;
        RECT 110.555 114.180 110.715 114.290 ;
        RECT 111.465 114.135 111.635 114.325 ;
        RECT 112.845 114.135 113.015 114.325 ;
        RECT 116.535 114.180 116.695 114.290 ;
        RECT 118.365 114.135 118.535 114.345 ;
        RECT 5.525 113.325 6.895 114.135 ;
        RECT 7.105 113.455 17.475 114.135 ;
        RECT 7.105 113.225 9.315 113.455 ;
        RECT 12.035 113.235 12.965 113.455 ;
        RECT 17.495 113.225 18.845 114.135 ;
        RECT 18.865 113.325 20.235 114.135 ;
        RECT 20.245 113.355 21.615 114.135 ;
        RECT 21.625 113.355 22.995 114.135 ;
        RECT 23.015 113.225 24.365 114.135 ;
        RECT 24.385 113.325 25.755 114.135 ;
        RECT 25.765 113.355 27.135 114.135 ;
        RECT 27.145 113.325 30.815 114.135 ;
        RECT 31.295 113.265 31.725 114.050 ;
        RECT 31.745 113.355 33.115 114.135 ;
        RECT 33.125 113.325 36.795 114.135 ;
        RECT 36.805 113.325 38.175 114.135 ;
        RECT 38.185 113.355 39.555 114.135 ;
        RECT 39.575 113.225 40.925 114.135 ;
        RECT 40.945 113.325 44.615 114.135 ;
        RECT 44.635 113.225 45.985 114.135 ;
        RECT 46.005 113.325 48.755 114.135 ;
        RECT 49.225 113.355 50.595 114.135 ;
        RECT 50.745 113.225 53.355 114.135 ;
        RECT 54.295 113.225 55.645 114.135 ;
        RECT 55.675 113.225 57.025 114.135 ;
        RECT 57.055 113.265 57.485 114.050 ;
        RECT 57.505 113.325 63.015 114.135 ;
        RECT 63.485 113.355 64.855 114.135 ;
        RECT 64.865 113.325 66.695 114.135 ;
        RECT 67.175 113.225 68.525 114.135 ;
        RECT 68.545 113.325 70.375 114.135 ;
        RECT 70.985 113.225 73.595 114.135 ;
        RECT 73.605 113.325 74.975 114.135 ;
        RECT 74.985 113.355 76.355 114.135 ;
        RECT 76.365 113.325 80.035 114.135 ;
        RECT 80.965 113.355 82.335 114.135 ;
        RECT 82.815 113.265 83.245 114.050 ;
        RECT 83.265 113.325 88.775 114.135 ;
        RECT 88.785 113.325 94.295 114.135 ;
        RECT 94.305 113.325 97.055 114.135 ;
        RECT 97.525 113.355 98.895 114.135 ;
        RECT 99.825 113.355 101.195 114.135 ;
        RECT 101.215 113.225 102.565 114.135 ;
        RECT 102.585 113.325 104.415 114.135 ;
        RECT 104.425 113.355 105.795 114.135 ;
        RECT 105.805 113.325 108.555 114.135 ;
        RECT 108.575 113.265 109.005 114.050 ;
        RECT 109.035 113.225 110.385 114.135 ;
        RECT 111.335 113.225 112.685 114.135 ;
        RECT 112.705 113.325 116.375 114.135 ;
        RECT 117.305 113.325 118.675 114.135 ;
      LAYER nwell ;
        RECT 5.330 110.105 118.870 112.935 ;
      LAYER pwell ;
        RECT 5.525 108.905 6.895 109.715 ;
        RECT 6.905 108.905 9.655 109.715 ;
        RECT 9.665 108.905 11.035 109.685 ;
        RECT 11.045 108.905 12.415 109.685 ;
        RECT 12.435 108.905 13.785 109.815 ;
        RECT 13.805 108.905 17.475 109.715 ;
        RECT 18.415 108.990 18.845 109.775 ;
        RECT 18.865 108.905 24.375 109.715 ;
        RECT 24.385 108.905 29.895 109.715 ;
        RECT 30.320 108.905 31.275 109.585 ;
        RECT 31.370 108.905 40.475 109.585 ;
        RECT 40.485 108.905 44.155 109.715 ;
        RECT 44.175 108.990 44.605 109.775 ;
        RECT 44.625 108.905 50.135 109.715 ;
        RECT 50.145 108.905 51.515 109.715 ;
        RECT 51.535 108.905 52.885 109.815 ;
        RECT 52.905 108.905 58.415 109.715 ;
        RECT 58.425 108.905 63.935 109.715 ;
        RECT 63.945 108.905 69.455 109.715 ;
        RECT 69.935 108.990 70.365 109.775 ;
        RECT 70.385 108.905 75.895 109.715 ;
        RECT 75.905 108.905 81.415 109.715 ;
        RECT 81.425 108.905 85.095 109.715 ;
        RECT 86.025 108.905 95.130 109.585 ;
        RECT 95.695 108.990 96.125 109.775 ;
        RECT 96.145 108.905 97.975 109.715 ;
        RECT 97.995 108.905 99.345 109.815 ;
        RECT 99.365 108.905 104.875 109.715 ;
        RECT 104.885 108.905 106.715 109.715 ;
        RECT 111.235 109.585 112.165 109.805 ;
        RECT 114.885 109.585 117.095 109.815 ;
        RECT 106.725 108.905 117.095 109.585 ;
        RECT 117.305 108.905 118.675 109.715 ;
        RECT 5.665 108.695 5.835 108.905 ;
        RECT 7.045 108.695 7.215 108.905 ;
        RECT 9.805 108.715 9.975 108.905 ;
        RECT 11.185 108.715 11.355 108.905 ;
        RECT 12.565 108.695 12.735 108.885 ;
        RECT 13.485 108.715 13.655 108.905 ;
        RECT 13.945 108.715 14.115 108.905 ;
        RECT 17.635 108.750 17.795 108.860 ;
        RECT 18.360 108.695 18.530 108.885 ;
        RECT 19.005 108.715 19.175 108.905 ;
        RECT 22.225 108.695 22.395 108.885 ;
        RECT 24.525 108.715 24.695 108.905 ;
        RECT 24.985 108.695 25.155 108.885 ;
        RECT 25.445 108.695 25.615 108.885 ;
        RECT 30.045 108.715 30.215 108.885 ;
        RECT 30.960 108.745 31.080 108.855 ;
        RECT 31.885 108.695 32.055 108.885 ;
        RECT 33.265 108.695 33.435 108.885 ;
        RECT 36.020 108.745 36.140 108.855 ;
        RECT 40.165 108.715 40.335 108.905 ;
        RECT 40.625 108.715 40.795 108.905 ;
        RECT 44.765 108.715 44.935 108.905 ;
        RECT 45.685 108.695 45.855 108.885 ;
        RECT 46.140 108.745 46.260 108.855 ;
        RECT 46.605 108.695 46.775 108.885 ;
        RECT 50.285 108.715 50.455 108.905 ;
        RECT 51.665 108.715 51.835 108.905 ;
        RECT 53.045 108.715 53.215 108.905 ;
        RECT 56.275 108.740 56.435 108.850 ;
        RECT 57.645 108.695 57.815 108.885 ;
        RECT 58.565 108.715 58.735 108.905 ;
        RECT 63.175 108.740 63.335 108.850 ;
        RECT 64.085 108.715 64.255 108.905 ;
        RECT 65.005 108.695 65.175 108.885 ;
        RECT 65.460 108.745 65.580 108.855 ;
        RECT 66.845 108.695 67.015 108.885 ;
        RECT 67.305 108.695 67.475 108.885 ;
        RECT 69.600 108.745 69.720 108.855 ;
        RECT 70.525 108.715 70.695 108.905 ;
        RECT 72.825 108.695 72.995 108.885 ;
        RECT 76.045 108.715 76.215 108.905 ;
        RECT 78.345 108.695 78.515 108.885 ;
        RECT 80.645 108.695 80.815 108.885 ;
        RECT 81.105 108.695 81.275 108.885 ;
        RECT 81.565 108.715 81.735 108.905 ;
        RECT 83.400 108.745 83.520 108.855 ;
        RECT 85.255 108.750 85.415 108.860 ;
        RECT 86.165 108.715 86.335 108.905 ;
        RECT 87.270 108.695 87.440 108.885 ;
        RECT 88.005 108.695 88.175 108.885 ;
        RECT 89.385 108.695 89.555 108.885 ;
        RECT 93.065 108.695 93.235 108.885 ;
        RECT 94.455 108.740 94.615 108.850 ;
        RECT 95.360 108.745 95.480 108.855 ;
        RECT 96.285 108.695 96.455 108.905 ;
        RECT 96.740 108.745 96.860 108.855 ;
        RECT 97.205 108.695 97.375 108.885 ;
        RECT 98.125 108.715 98.295 108.905 ;
        RECT 98.580 108.745 98.700 108.855 ;
        RECT 99.505 108.715 99.675 108.905 ;
        RECT 105.025 108.715 105.195 108.905 ;
        RECT 106.865 108.715 107.035 108.905 ;
        RECT 108.245 108.695 108.415 108.885 ;
        RECT 109.160 108.745 109.280 108.855 ;
        RECT 109.625 108.695 109.795 108.885 ;
        RECT 111.925 108.695 112.095 108.885 ;
        RECT 112.385 108.695 112.555 108.885 ;
        RECT 116.065 108.695 116.235 108.885 ;
        RECT 118.365 108.695 118.535 108.905 ;
        RECT 5.525 107.885 6.895 108.695 ;
        RECT 6.905 107.885 12.415 108.695 ;
        RECT 12.425 107.885 17.935 108.695 ;
        RECT 17.945 108.015 21.845 108.695 ;
        RECT 17.945 107.785 18.875 108.015 ;
        RECT 22.085 107.885 23.915 108.695 ;
        RECT 23.925 107.915 25.295 108.695 ;
        RECT 25.305 107.885 30.815 108.695 ;
        RECT 31.295 107.825 31.725 108.610 ;
        RECT 31.745 107.915 33.115 108.695 ;
        RECT 33.125 107.885 35.875 108.695 ;
        RECT 36.715 108.015 45.995 108.695 ;
        RECT 46.465 108.015 55.745 108.695 ;
        RECT 36.715 107.895 39.050 108.015 ;
        RECT 36.715 107.785 37.635 107.895 ;
        RECT 43.715 107.795 44.635 108.015 ;
        RECT 47.825 107.795 48.745 108.015 ;
        RECT 53.410 107.895 55.745 108.015 ;
        RECT 54.825 107.785 55.745 107.895 ;
        RECT 57.055 107.825 57.485 108.610 ;
        RECT 57.505 107.885 63.015 108.695 ;
        RECT 63.945 107.915 65.315 108.695 ;
        RECT 65.795 107.785 67.145 108.695 ;
        RECT 67.165 107.885 72.675 108.695 ;
        RECT 72.685 107.885 78.195 108.695 ;
        RECT 78.205 107.885 79.575 108.695 ;
        RECT 79.585 107.915 80.955 108.695 ;
        RECT 80.965 107.885 82.795 108.695 ;
        RECT 82.815 107.825 83.245 108.610 ;
        RECT 83.955 108.015 87.855 108.695 ;
        RECT 86.925 107.785 87.855 108.015 ;
        RECT 87.875 107.785 89.225 108.695 ;
        RECT 89.245 107.885 92.915 108.695 ;
        RECT 92.925 107.915 94.295 108.695 ;
        RECT 95.225 107.915 96.595 108.695 ;
        RECT 97.075 107.785 98.425 108.695 ;
        RECT 99.275 108.015 108.555 108.695 ;
        RECT 99.275 107.895 101.610 108.015 ;
        RECT 99.275 107.785 100.195 107.895 ;
        RECT 106.275 107.795 107.195 108.015 ;
        RECT 108.575 107.825 109.005 108.610 ;
        RECT 109.495 107.785 110.845 108.695 ;
        RECT 110.865 107.915 112.235 108.695 ;
        RECT 112.245 107.885 115.915 108.695 ;
        RECT 115.925 107.885 117.295 108.695 ;
        RECT 117.305 107.885 118.675 108.695 ;
      LAYER nwell ;
        RECT 5.330 104.665 118.870 107.495 ;
      LAYER pwell ;
        RECT 5.525 103.465 6.895 104.275 ;
        RECT 6.905 103.465 12.415 104.275 ;
        RECT 12.425 103.465 16.095 104.275 ;
        RECT 16.565 103.465 17.935 104.245 ;
        RECT 18.415 103.550 18.845 104.335 ;
        RECT 18.875 103.465 20.225 104.375 ;
        RECT 22.525 104.145 23.445 104.365 ;
        RECT 29.525 104.265 30.445 104.375 ;
        RECT 28.110 104.145 30.445 104.265 ;
        RECT 32.185 104.145 33.105 104.365 ;
        RECT 39.185 104.265 40.105 104.375 ;
        RECT 37.770 104.145 40.105 104.265 ;
        RECT 21.165 103.465 30.445 104.145 ;
        RECT 30.825 103.465 40.105 104.145 ;
        RECT 41.415 103.465 42.765 104.375 ;
        RECT 42.795 103.465 44.145 104.375 ;
        RECT 44.175 103.550 44.605 104.335 ;
        RECT 44.625 103.465 45.995 104.245 ;
        RECT 49.665 104.145 50.595 104.375 ;
        RECT 51.965 104.145 52.885 104.365 ;
        RECT 58.965 104.265 59.885 104.375 ;
        RECT 57.550 104.145 59.885 104.265 ;
        RECT 61.625 104.145 62.545 104.365 ;
        RECT 68.625 104.265 69.545 104.375 ;
        RECT 67.210 104.145 69.545 104.265 ;
        RECT 46.695 103.465 50.595 104.145 ;
        RECT 50.605 103.465 59.885 104.145 ;
        RECT 60.265 103.465 69.545 104.145 ;
        RECT 69.935 103.550 70.365 104.335 ;
        RECT 70.395 103.465 71.745 104.375 ;
        RECT 71.765 103.465 75.435 104.275 ;
        RECT 77.725 104.145 78.645 104.365 ;
        RECT 84.725 104.265 85.645 104.375 ;
        RECT 83.310 104.145 85.645 104.265 ;
        RECT 87.385 104.145 88.305 104.365 ;
        RECT 94.385 104.265 95.305 104.375 ;
        RECT 92.970 104.145 95.305 104.265 ;
        RECT 76.365 103.465 85.645 104.145 ;
        RECT 86.025 103.465 95.305 104.145 ;
        RECT 95.695 103.550 96.125 104.335 ;
        RECT 96.515 104.265 97.435 104.375 ;
        RECT 96.515 104.145 98.850 104.265 ;
        RECT 103.515 104.145 104.435 104.365 ;
        RECT 107.165 104.145 108.085 104.365 ;
        RECT 114.165 104.265 115.085 104.375 ;
        RECT 112.750 104.145 115.085 104.265 ;
        RECT 96.515 103.465 105.795 104.145 ;
        RECT 105.805 103.465 115.085 104.145 ;
        RECT 115.475 103.465 116.825 104.375 ;
        RECT 117.305 103.465 118.675 104.275 ;
        RECT 5.665 103.255 5.835 103.465 ;
        RECT 7.045 103.255 7.215 103.465 ;
        RECT 10.735 103.300 10.895 103.410 ;
        RECT 12.565 103.255 12.735 103.465 ;
        RECT 13.020 103.305 13.140 103.415 ;
        RECT 14.405 103.255 14.575 103.445 ;
        RECT 14.865 103.255 15.035 103.445 ;
        RECT 16.240 103.305 16.360 103.415 ;
        RECT 17.625 103.275 17.795 103.465 ;
        RECT 18.080 103.305 18.200 103.415 ;
        RECT 19.005 103.275 19.175 103.465 ;
        RECT 20.395 103.310 20.555 103.420 ;
        RECT 21.305 103.275 21.475 103.465 ;
        RECT 24.800 103.255 24.970 103.445 ;
        RECT 29.585 103.255 29.755 103.445 ;
        RECT 30.045 103.255 30.215 103.445 ;
        RECT 30.965 103.275 31.135 103.465 ;
        RECT 32.160 103.255 32.330 103.445 ;
        RECT 36.025 103.255 36.195 103.445 ;
        RECT 37.860 103.305 37.980 103.415 ;
        RECT 40.635 103.310 40.795 103.420 ;
        RECT 41.730 103.255 41.900 103.445 ;
        RECT 42.465 103.255 42.635 103.465 ;
        RECT 43.845 103.275 44.015 103.465 ;
        RECT 45.685 103.275 45.855 103.465 ;
        RECT 46.140 103.305 46.260 103.415 ;
        RECT 48.905 103.255 49.075 103.445 ;
        RECT 49.360 103.305 49.480 103.415 ;
        RECT 49.825 103.255 49.995 103.445 ;
        RECT 50.010 103.275 50.180 103.465 ;
        RECT 50.745 103.275 50.915 103.465 ;
        RECT 51.205 103.255 51.375 103.445 ;
        RECT 52.860 103.255 53.030 103.445 ;
        RECT 56.720 103.305 56.840 103.415 ;
        RECT 58.565 103.255 58.735 103.445 ;
        RECT 59.025 103.255 59.195 103.445 ;
        RECT 60.405 103.275 60.575 103.465 ;
        RECT 62.700 103.305 62.820 103.415 ;
        RECT 63.165 103.255 63.335 103.445 ;
        RECT 64.545 103.255 64.715 103.445 ;
        RECT 71.445 103.275 71.615 103.465 ;
        RECT 71.905 103.275 72.075 103.465 ;
        RECT 74.215 103.300 74.375 103.410 ;
        RECT 75.125 103.255 75.295 103.445 ;
        RECT 75.595 103.310 75.755 103.420 ;
        RECT 76.505 103.275 76.675 103.465 ;
        RECT 77.430 103.255 77.600 103.445 ;
        RECT 80.185 103.255 80.355 103.445 ;
        RECT 82.485 103.255 82.655 103.445 ;
        RECT 83.680 103.255 83.850 103.445 ;
        RECT 86.165 103.275 86.335 103.465 ;
        RECT 87.545 103.255 87.715 103.445 ;
        RECT 88.920 103.305 89.040 103.415 ;
        RECT 92.790 103.255 92.960 103.445 ;
        RECT 93.525 103.255 93.695 103.445 ;
        RECT 103.185 103.255 103.355 103.445 ;
        RECT 105.485 103.275 105.655 103.465 ;
        RECT 105.945 103.255 106.115 103.465 ;
        RECT 107.325 103.255 107.495 103.445 ;
        RECT 112.570 103.255 112.740 103.445 ;
        RECT 113.305 103.255 113.475 103.445 ;
        RECT 115.605 103.275 115.775 103.465 ;
        RECT 116.980 103.305 117.100 103.415 ;
        RECT 118.365 103.255 118.535 103.465 ;
        RECT 5.525 102.445 6.895 103.255 ;
        RECT 6.905 102.445 10.575 103.255 ;
        RECT 11.505 102.475 12.875 103.255 ;
        RECT 13.355 102.345 14.705 103.255 ;
        RECT 14.725 102.575 24.005 103.255 ;
        RECT 16.085 102.355 17.005 102.575 ;
        RECT 21.670 102.455 24.005 102.575 ;
        RECT 23.085 102.345 24.005 102.455 ;
        RECT 24.385 102.575 28.285 103.255 ;
        RECT 24.385 102.345 25.315 102.575 ;
        RECT 28.535 102.345 29.885 103.255 ;
        RECT 29.905 102.445 31.275 103.255 ;
        RECT 31.295 102.385 31.725 103.170 ;
        RECT 31.745 102.575 35.645 103.255 ;
        RECT 31.745 102.345 32.675 102.575 ;
        RECT 35.885 102.445 37.715 103.255 ;
        RECT 38.415 102.575 42.315 103.255 ;
        RECT 41.385 102.345 42.315 102.575 ;
        RECT 42.325 102.445 47.835 103.255 ;
        RECT 47.845 102.475 49.215 103.255 ;
        RECT 49.695 102.345 51.045 103.255 ;
        RECT 51.065 102.475 52.435 103.255 ;
        RECT 52.445 102.575 56.345 103.255 ;
        RECT 52.445 102.345 53.375 102.575 ;
        RECT 57.055 102.385 57.485 103.170 ;
        RECT 57.515 102.345 58.865 103.255 ;
        RECT 58.885 102.445 62.555 103.255 ;
        RECT 63.025 102.475 64.395 103.255 ;
        RECT 64.405 102.575 73.685 103.255 ;
        RECT 65.765 102.355 66.685 102.575 ;
        RECT 71.350 102.455 73.685 102.575 ;
        RECT 72.765 102.345 73.685 102.455 ;
        RECT 74.995 102.345 76.345 103.255 ;
        RECT 77.285 102.345 79.895 103.255 ;
        RECT 80.045 102.445 81.415 103.255 ;
        RECT 81.435 102.345 82.785 103.255 ;
        RECT 82.815 102.385 83.245 103.170 ;
        RECT 83.265 102.575 87.165 103.255 ;
        RECT 83.265 102.345 84.195 102.575 ;
        RECT 87.405 102.475 88.775 103.255 ;
        RECT 89.475 102.575 93.375 103.255 ;
        RECT 93.385 102.575 102.665 103.255 ;
        RECT 92.445 102.345 93.375 102.575 ;
        RECT 94.745 102.355 95.665 102.575 ;
        RECT 100.330 102.455 102.665 102.575 ;
        RECT 101.745 102.345 102.665 102.455 ;
        RECT 103.045 102.445 105.795 103.255 ;
        RECT 105.805 102.475 107.175 103.255 ;
        RECT 107.185 102.445 108.555 103.255 ;
        RECT 108.575 102.385 109.005 103.170 ;
        RECT 109.255 102.575 113.155 103.255 ;
        RECT 112.225 102.345 113.155 102.575 ;
        RECT 113.165 102.445 116.835 103.255 ;
        RECT 117.305 102.445 118.675 103.255 ;
      LAYER nwell ;
        RECT 5.330 99.225 118.870 102.055 ;
      LAYER pwell ;
        RECT 5.525 98.025 6.895 98.835 ;
        RECT 6.905 98.025 8.275 98.835 ;
        RECT 9.645 98.705 10.565 98.925 ;
        RECT 16.645 98.825 17.565 98.935 ;
        RECT 15.230 98.705 17.565 98.825 ;
        RECT 8.285 98.025 17.565 98.705 ;
        RECT 18.415 98.110 18.845 98.895 ;
        RECT 18.865 98.705 19.795 98.935 ;
        RECT 18.865 98.025 22.765 98.705 ;
        RECT 23.005 98.025 28.515 98.835 ;
        RECT 28.525 98.025 34.035 98.835 ;
        RECT 34.045 98.025 37.715 98.835 ;
        RECT 37.725 98.025 39.095 98.835 ;
        RECT 39.115 98.025 40.465 98.935 ;
        RECT 40.485 98.025 44.155 98.835 ;
        RECT 44.175 98.110 44.605 98.895 ;
        RECT 44.625 98.025 48.295 98.835 ;
        RECT 48.305 98.025 49.675 98.805 ;
        RECT 50.155 98.025 51.505 98.935 ;
        RECT 51.525 98.025 57.035 98.835 ;
        RECT 57.045 98.025 62.555 98.835 ;
        RECT 62.565 98.025 65.315 98.835 ;
        RECT 65.325 98.705 66.255 98.935 ;
        RECT 65.325 98.025 69.225 98.705 ;
        RECT 69.935 98.110 70.365 98.895 ;
        RECT 72.205 98.705 73.125 98.925 ;
        RECT 79.205 98.825 80.125 98.935 ;
        RECT 77.790 98.705 80.125 98.825 ;
        RECT 70.845 98.025 80.125 98.705 ;
        RECT 80.505 98.025 86.015 98.835 ;
        RECT 86.025 98.025 91.535 98.835 ;
        RECT 91.545 98.025 95.215 98.835 ;
        RECT 95.695 98.110 96.125 98.895 ;
        RECT 96.145 98.705 97.075 98.935 ;
        RECT 96.145 98.025 100.045 98.705 ;
        RECT 100.285 98.025 105.795 98.835 ;
        RECT 106.265 98.705 107.195 98.935 ;
        RECT 106.265 98.025 110.165 98.705 ;
        RECT 110.405 98.025 115.915 98.835 ;
        RECT 115.925 98.025 117.295 98.835 ;
        RECT 117.305 98.025 118.675 98.835 ;
        RECT 5.665 97.815 5.835 98.025 ;
        RECT 7.045 97.815 7.215 98.025 ;
        RECT 8.425 97.815 8.595 98.025 ;
        RECT 18.080 97.865 18.200 97.975 ;
        RECT 18.360 97.815 18.530 98.005 ;
        RECT 19.280 97.835 19.450 98.025 ;
        RECT 22.225 97.815 22.395 98.005 ;
        RECT 23.145 97.835 23.315 98.025 ;
        RECT 27.745 97.815 27.915 98.005 ;
        RECT 28.665 97.835 28.835 98.025 ;
        RECT 33.725 97.835 33.895 98.005 ;
        RECT 34.185 97.835 34.355 98.025 ;
        RECT 37.865 97.835 38.035 98.025 ;
        RECT 40.165 97.835 40.335 98.025 ;
        RECT 40.625 97.835 40.795 98.025 ;
        RECT 33.725 97.815 33.875 97.835 ;
        RECT 43.385 97.815 43.555 98.005 ;
        RECT 43.845 97.815 44.015 98.005 ;
        RECT 44.765 97.835 44.935 98.025 ;
        RECT 45.685 97.815 45.855 98.005 ;
        RECT 49.365 97.835 49.535 98.025 ;
        RECT 49.820 97.865 49.940 97.975 ;
        RECT 50.285 97.835 50.455 98.025 ;
        RECT 51.665 97.835 51.835 98.025 ;
        RECT 55.345 97.815 55.515 98.005 ;
        RECT 57.185 97.835 57.355 98.025 ;
        RECT 57.640 97.865 57.760 97.975 ;
        RECT 60.405 97.815 60.575 98.005 ;
        RECT 60.875 97.860 61.035 97.970 ;
        RECT 62.705 97.815 62.875 98.025 ;
        RECT 63.160 97.865 63.280 97.975 ;
        RECT 63.625 97.815 63.795 98.005 ;
        RECT 65.005 97.815 65.175 98.005 ;
        RECT 65.740 97.835 65.910 98.025 ;
        RECT 68.685 97.815 68.855 98.005 ;
        RECT 69.600 97.865 69.720 97.975 ;
        RECT 70.340 97.815 70.510 98.005 ;
        RECT 70.520 97.865 70.640 97.975 ;
        RECT 70.985 97.835 71.155 98.025 ;
        RECT 75.125 97.815 75.295 98.005 ;
        RECT 75.585 97.815 75.755 98.005 ;
        RECT 80.645 97.835 80.815 98.025 ;
        RECT 81.105 97.815 81.275 98.005 ;
        RECT 83.405 97.815 83.575 98.005 ;
        RECT 86.165 97.835 86.335 98.025 ;
        RECT 86.185 97.815 86.335 97.835 ;
        RECT 90.305 97.835 90.475 98.005 ;
        RECT 90.765 97.835 90.935 98.005 ;
        RECT 91.685 97.835 91.855 98.025 ;
        RECT 90.305 97.815 90.455 97.835 ;
        RECT 5.525 97.005 6.895 97.815 ;
        RECT 6.905 97.005 8.275 97.815 ;
        RECT 8.285 97.135 17.565 97.815 ;
        RECT 9.645 96.915 10.565 97.135 ;
        RECT 15.230 97.015 17.565 97.135 ;
        RECT 16.645 96.905 17.565 97.015 ;
        RECT 17.945 97.135 21.845 97.815 ;
        RECT 17.945 96.905 18.875 97.135 ;
        RECT 22.085 97.005 27.595 97.815 ;
        RECT 27.605 97.005 31.275 97.815 ;
        RECT 31.295 96.945 31.725 97.730 ;
        RECT 31.945 96.995 33.875 97.815 ;
        RECT 34.415 97.135 43.695 97.815 ;
        RECT 34.415 97.015 36.750 97.135 ;
        RECT 31.945 96.905 32.895 96.995 ;
        RECT 34.415 96.905 35.335 97.015 ;
        RECT 41.415 96.915 42.335 97.135 ;
        RECT 43.705 97.005 45.535 97.815 ;
        RECT 45.545 97.135 54.825 97.815 ;
        RECT 46.905 96.915 47.825 97.135 ;
        RECT 52.490 97.015 54.825 97.135 ;
        RECT 53.905 96.905 54.825 97.015 ;
        RECT 55.205 97.005 57.035 97.815 ;
        RECT 57.055 96.945 57.485 97.730 ;
        RECT 57.975 97.135 60.715 97.815 ;
        RECT 61.645 97.035 63.015 97.815 ;
        RECT 63.495 96.905 64.845 97.815 ;
        RECT 64.865 97.005 68.535 97.815 ;
        RECT 68.545 97.005 69.915 97.815 ;
        RECT 69.925 97.135 73.825 97.815 ;
        RECT 69.925 96.905 70.855 97.135 ;
        RECT 74.065 97.035 75.435 97.815 ;
        RECT 75.445 97.005 80.955 97.815 ;
        RECT 80.965 97.005 82.795 97.815 ;
        RECT 82.815 96.945 83.245 97.730 ;
        RECT 83.265 97.135 86.005 97.815 ;
        RECT 86.185 96.995 88.115 97.815 ;
        RECT 87.165 96.905 88.115 96.995 ;
        RECT 88.525 96.995 90.455 97.815 ;
        RECT 90.785 97.815 90.935 97.835 ;
        RECT 93.065 97.815 93.235 98.005 ;
        RECT 95.360 97.865 95.480 97.975 ;
        RECT 96.285 97.835 96.455 98.005 ;
        RECT 96.560 97.835 96.730 98.025 ;
        RECT 96.285 97.815 96.435 97.835 ;
        RECT 96.745 97.815 96.915 98.005 ;
        RECT 100.425 97.835 100.595 98.025 ;
        RECT 102.265 97.815 102.435 98.005 ;
        RECT 105.940 97.865 106.060 97.975 ;
        RECT 106.680 97.835 106.850 98.025 ;
        RECT 107.795 97.860 107.955 97.970 ;
        RECT 110.085 97.815 110.255 98.005 ;
        RECT 110.545 97.975 110.715 98.025 ;
        RECT 110.540 97.865 110.715 97.975 ;
        RECT 110.545 97.835 110.715 97.865 ;
        RECT 111.005 97.815 111.175 98.005 ;
        RECT 112.385 97.815 112.555 98.005 ;
        RECT 116.065 97.815 116.235 98.025 ;
        RECT 118.365 97.815 118.535 98.025 ;
        RECT 90.785 96.995 92.715 97.815 ;
        RECT 92.925 97.005 94.295 97.815 ;
        RECT 88.525 96.905 89.475 96.995 ;
        RECT 91.765 96.905 92.715 96.995 ;
        RECT 94.505 96.995 96.435 97.815 ;
        RECT 96.605 97.005 102.115 97.815 ;
        RECT 102.125 97.005 107.635 97.815 ;
        RECT 94.505 96.905 95.455 96.995 ;
        RECT 108.575 96.945 109.005 97.730 ;
        RECT 109.025 97.035 110.395 97.815 ;
        RECT 110.875 96.905 112.225 97.815 ;
        RECT 112.245 97.005 115.915 97.815 ;
        RECT 115.925 97.005 117.295 97.815 ;
        RECT 117.305 97.005 118.675 97.815 ;
      LAYER nwell ;
        RECT 5.330 93.785 118.870 96.615 ;
      LAYER pwell ;
        RECT 5.525 92.585 6.895 93.395 ;
        RECT 6.905 92.585 12.415 93.395 ;
        RECT 12.425 92.585 13.795 93.365 ;
        RECT 13.815 92.585 15.165 93.495 ;
        RECT 15.185 92.585 17.935 93.395 ;
        RECT 18.415 92.670 18.845 93.455 ;
        RECT 20.465 93.405 21.415 93.495 ;
        RECT 19.485 92.585 21.415 93.405 ;
        RECT 21.825 93.405 22.775 93.495 ;
        RECT 25.065 93.405 26.015 93.495 ;
        RECT 27.365 93.405 28.315 93.495 ;
        RECT 21.825 92.585 23.755 93.405 ;
        RECT 5.665 92.375 5.835 92.585 ;
        RECT 7.045 92.375 7.215 92.585 ;
        RECT 12.565 92.375 12.735 92.565 ;
        RECT 13.485 92.395 13.655 92.585 ;
        RECT 14.865 92.395 15.035 92.585 ;
        RECT 15.325 92.395 15.495 92.585 ;
        RECT 19.485 92.565 19.635 92.585 ;
        RECT 23.605 92.565 23.755 92.585 ;
        RECT 24.085 92.585 26.015 93.405 ;
        RECT 26.385 92.585 28.315 93.405 ;
        RECT 28.610 92.585 37.715 93.265 ;
        RECT 37.725 92.585 39.095 93.365 ;
        RECT 42.765 93.265 43.695 93.495 ;
        RECT 39.795 92.585 43.695 93.265 ;
        RECT 44.175 92.670 44.605 93.455 ;
        RECT 48.985 93.405 49.935 93.495 ;
        RECT 44.625 92.585 45.995 93.365 ;
        RECT 46.005 92.585 47.835 93.395 ;
        RECT 48.005 92.585 49.935 93.405 ;
        RECT 50.145 93.265 51.075 93.495 ;
        RECT 54.485 93.405 55.435 93.495 ;
        RECT 56.785 93.405 57.735 93.495 ;
        RECT 50.145 92.585 54.045 93.265 ;
        RECT 54.485 92.585 56.415 93.405 ;
        RECT 56.785 92.585 58.715 93.405 ;
        RECT 60.245 93.265 61.165 93.485 ;
        RECT 67.245 93.385 68.165 93.495 ;
        RECT 65.830 93.265 68.165 93.385 ;
        RECT 58.885 92.585 68.165 93.265 ;
        RECT 68.545 92.585 69.915 93.395 ;
        RECT 69.935 92.670 70.365 93.455 ;
        RECT 70.385 92.585 74.055 93.395 ;
        RECT 74.525 93.265 75.455 93.495 ;
        RECT 83.925 93.405 84.875 93.495 ;
        RECT 88.985 93.405 89.935 93.495 ;
        RECT 91.285 93.405 92.235 93.495 ;
        RECT 74.525 92.585 78.425 93.265 ;
        RECT 78.665 92.585 82.335 93.395 ;
        RECT 82.345 92.585 83.715 93.395 ;
        RECT 83.925 92.585 85.855 93.405 ;
        RECT 86.025 92.585 88.115 93.395 ;
        RECT 88.985 92.585 90.915 93.405 ;
        RECT 91.285 92.585 93.215 93.405 ;
        RECT 93.385 92.585 94.755 93.365 ;
        RECT 95.695 92.670 96.125 93.455 ;
        RECT 96.145 92.585 97.975 93.395 ;
        RECT 98.455 92.585 99.805 93.495 ;
        RECT 99.825 92.585 105.335 93.395 ;
        RECT 107.625 93.265 108.545 93.485 ;
        RECT 114.625 93.385 115.545 93.495 ;
        RECT 113.210 93.265 115.545 93.385 ;
        RECT 106.265 92.585 115.545 93.265 ;
        RECT 115.925 92.585 117.295 93.395 ;
        RECT 117.305 92.585 118.675 93.395 ;
        RECT 24.085 92.565 24.235 92.585 ;
        RECT 26.385 92.565 26.535 92.585 ;
        RECT 18.085 92.535 18.255 92.565 ;
        RECT 18.080 92.425 18.255 92.535 ;
        RECT 19.000 92.425 19.120 92.535 ;
        RECT 18.085 92.375 18.255 92.425 ;
        RECT 19.465 92.395 19.635 92.565 ;
        RECT 20.840 92.425 20.960 92.535 ;
        RECT 21.305 92.395 21.475 92.565 ;
        RECT 21.325 92.375 21.475 92.395 ;
        RECT 23.605 92.375 23.775 92.565 ;
        RECT 24.065 92.395 24.235 92.565 ;
        RECT 26.365 92.395 26.535 92.565 ;
        RECT 29.125 92.375 29.295 92.565 ;
        RECT 30.960 92.425 31.080 92.535 ;
        RECT 31.890 92.375 32.060 92.565 ;
        RECT 37.405 92.395 37.575 92.585 ;
        RECT 38.785 92.395 38.955 92.585 ;
        RECT 39.240 92.425 39.360 92.535 ;
        RECT 43.110 92.395 43.280 92.585 ;
        RECT 43.845 92.535 44.015 92.565 ;
        RECT 43.840 92.425 44.015 92.535 ;
        RECT 43.845 92.375 44.015 92.425 ;
        RECT 44.305 92.375 44.475 92.565 ;
        RECT 45.685 92.395 45.855 92.585 ;
        RECT 46.145 92.395 46.315 92.585 ;
        RECT 48.005 92.565 48.155 92.585 ;
        RECT 47.985 92.395 48.155 92.565 ;
        RECT 49.825 92.375 49.995 92.565 ;
        RECT 50.560 92.395 50.730 92.585 ;
        RECT 56.265 92.565 56.415 92.585 ;
        RECT 58.565 92.565 58.715 92.585 ;
        RECT 52.585 92.395 52.755 92.565 ;
        RECT 52.605 92.375 52.755 92.395 ;
        RECT 54.885 92.375 55.055 92.565 ;
        RECT 56.265 92.395 56.435 92.565 ;
        RECT 56.720 92.425 56.840 92.535 ;
        RECT 58.565 92.395 58.735 92.565 ;
        RECT 59.025 92.375 59.195 92.585 ;
        RECT 59.485 92.395 59.655 92.565 ;
        RECT 59.505 92.375 59.655 92.395 ;
        RECT 61.785 92.375 61.955 92.565 ;
        RECT 63.900 92.375 64.070 92.565 ;
        RECT 67.765 92.375 67.935 92.565 ;
        RECT 68.685 92.395 68.855 92.585 ;
        RECT 70.525 92.395 70.695 92.585 ;
        RECT 73.285 92.375 73.455 92.565 ;
        RECT 74.200 92.425 74.320 92.535 ;
        RECT 74.940 92.395 75.110 92.585 ;
        RECT 78.805 92.375 78.975 92.585 ;
        RECT 82.485 92.535 82.655 92.585 ;
        RECT 85.705 92.565 85.855 92.585 ;
        RECT 82.480 92.425 82.655 92.535 ;
        RECT 82.485 92.395 82.655 92.425 ;
        RECT 83.415 92.420 83.575 92.530 ;
        RECT 84.325 92.375 84.495 92.565 ;
        RECT 85.705 92.395 85.875 92.565 ;
        RECT 86.165 92.395 86.335 92.585 ;
        RECT 90.765 92.565 90.915 92.585 ;
        RECT 93.065 92.565 93.215 92.585 ;
        RECT 90.765 92.395 90.935 92.565 ;
        RECT 93.065 92.395 93.235 92.565 ;
        RECT 93.525 92.375 93.695 92.585 ;
        RECT 94.915 92.430 95.075 92.540 ;
        RECT 96.285 92.395 96.455 92.585 ;
        RECT 98.120 92.425 98.240 92.535 ;
        RECT 99.505 92.395 99.675 92.585 ;
        RECT 99.965 92.395 100.135 92.585 ;
        RECT 103.185 92.375 103.355 92.565 ;
        RECT 104.565 92.375 104.735 92.565 ;
        RECT 105.495 92.430 105.655 92.540 ;
        RECT 106.405 92.395 106.575 92.585 ;
        RECT 108.240 92.425 108.360 92.535 ;
        RECT 109.440 92.375 109.610 92.565 ;
        RECT 113.305 92.375 113.475 92.565 ;
        RECT 116.065 92.395 116.235 92.585 ;
        RECT 116.980 92.425 117.100 92.535 ;
        RECT 118.365 92.375 118.535 92.585 ;
        RECT 5.525 91.565 6.895 92.375 ;
        RECT 6.905 91.565 12.415 92.375 ;
        RECT 12.425 91.565 17.935 92.375 ;
        RECT 17.945 91.565 20.695 92.375 ;
        RECT 21.325 91.555 23.255 92.375 ;
        RECT 23.465 91.565 28.975 92.375 ;
        RECT 28.985 91.565 30.815 92.375 ;
        RECT 22.305 91.465 23.255 91.555 ;
        RECT 31.295 91.505 31.725 92.290 ;
        RECT 31.745 91.465 42.755 92.375 ;
        RECT 42.795 91.465 44.145 92.375 ;
        RECT 44.165 91.565 49.675 92.375 ;
        RECT 49.685 91.565 52.435 92.375 ;
        RECT 52.605 91.555 54.535 92.375 ;
        RECT 54.745 91.565 56.575 92.375 ;
        RECT 53.585 91.465 54.535 91.555 ;
        RECT 57.055 91.505 57.485 92.290 ;
        RECT 57.505 91.695 59.335 92.375 ;
        RECT 59.505 91.555 61.435 92.375 ;
        RECT 61.645 91.695 63.475 92.375 ;
        RECT 63.485 91.695 67.385 92.375 ;
        RECT 60.485 91.465 61.435 91.555 ;
        RECT 63.485 91.465 64.415 91.695 ;
        RECT 67.625 91.565 73.135 92.375 ;
        RECT 73.145 91.565 78.655 92.375 ;
        RECT 78.665 91.565 82.335 92.375 ;
        RECT 82.815 91.505 83.245 92.290 ;
        RECT 84.185 91.695 93.290 92.375 ;
        RECT 93.385 91.695 102.665 92.375 ;
        RECT 94.745 91.475 95.665 91.695 ;
        RECT 100.330 91.575 102.665 91.695 ;
        RECT 103.045 91.595 104.415 92.375 ;
        RECT 101.745 91.465 102.665 91.575 ;
        RECT 104.425 91.565 108.095 92.375 ;
        RECT 108.575 91.505 109.005 92.290 ;
        RECT 109.025 91.695 112.925 92.375 ;
        RECT 109.025 91.465 109.955 91.695 ;
        RECT 113.165 91.565 116.835 92.375 ;
        RECT 117.305 91.565 118.675 92.375 ;
      LAYER nwell ;
        RECT 5.330 88.345 118.870 91.175 ;
      LAYER pwell ;
        RECT 5.525 87.145 6.895 87.955 ;
        RECT 6.905 87.145 12.415 87.955 ;
        RECT 12.885 87.145 14.255 87.925 ;
        RECT 14.265 87.145 17.935 87.955 ;
        RECT 18.415 87.230 18.845 88.015 ;
        RECT 18.865 87.145 20.695 87.955 ;
        RECT 22.510 87.855 23.455 88.055 ;
        RECT 20.705 87.175 23.455 87.855 ;
        RECT 5.665 86.935 5.835 87.145 ;
        RECT 7.045 86.935 7.215 87.145 ;
        RECT 9.805 86.935 9.975 87.125 ;
        RECT 10.265 86.935 10.435 87.125 ;
        RECT 12.560 86.985 12.680 87.095 ;
        RECT 13.945 86.955 14.115 87.145 ;
        RECT 14.405 86.955 14.575 87.145 ;
        RECT 18.080 86.985 18.200 87.095 ;
        RECT 19.005 86.955 19.175 87.145 ;
        RECT 20.200 86.935 20.370 87.125 ;
        RECT 20.850 86.955 21.020 87.175 ;
        RECT 22.510 87.145 23.455 87.175 ;
        RECT 23.660 87.145 27.135 88.055 ;
        RECT 28.950 87.855 29.895 88.055 ;
        RECT 27.145 87.175 29.895 87.855 ;
        RECT 24.075 86.980 24.235 87.090 ;
        RECT 24.985 86.935 25.155 87.125 ;
        RECT 26.640 86.935 26.810 87.125 ;
        RECT 26.820 86.955 26.990 87.145 ;
        RECT 27.290 86.955 27.460 87.175 ;
        RECT 28.950 87.145 29.895 87.175 ;
        RECT 30.375 87.145 31.725 88.055 ;
        RECT 33.550 87.855 34.495 88.055 ;
        RECT 31.745 87.175 34.495 87.855 ;
        RECT 35.865 87.825 36.785 88.045 ;
        RECT 42.865 87.945 43.785 88.055 ;
        RECT 41.450 87.825 43.785 87.945 ;
        RECT 30.040 86.985 30.160 87.095 ;
        RECT 30.505 86.955 30.675 87.145 ;
        RECT 31.890 86.935 32.060 87.175 ;
        RECT 33.550 87.145 34.495 87.175 ;
        RECT 34.505 87.145 43.785 87.825 ;
        RECT 44.175 87.230 44.605 88.015 ;
        RECT 44.635 87.145 45.985 88.055 ;
        RECT 46.005 87.145 51.515 87.955 ;
        RECT 51.525 87.855 52.470 88.055 ;
        RECT 51.525 87.175 54.275 87.855 ;
        RECT 51.525 87.145 52.470 87.175 ;
        RECT 34.645 86.955 34.815 87.145 ;
        RECT 35.560 86.985 35.680 87.095 ;
        RECT 39.430 86.935 39.600 87.125 ;
        RECT 40.165 86.935 40.335 87.125 ;
        RECT 44.765 86.955 44.935 87.145 ;
        RECT 46.145 86.955 46.315 87.145 ;
        RECT 53.040 86.935 53.210 87.125 ;
        RECT 5.525 86.125 6.895 86.935 ;
        RECT 6.905 86.125 8.735 86.935 ;
        RECT 8.745 86.155 10.115 86.935 ;
        RECT 10.125 86.255 19.405 86.935 ;
        RECT 11.485 86.035 12.405 86.255 ;
        RECT 17.070 86.135 19.405 86.255 ;
        RECT 18.485 86.025 19.405 86.135 ;
        RECT 19.785 86.255 23.685 86.935 ;
        RECT 19.785 86.025 20.715 86.255 ;
        RECT 24.845 86.155 26.215 86.935 ;
        RECT 26.225 86.255 30.125 86.935 ;
        RECT 26.225 86.025 27.155 86.255 ;
        RECT 31.295 86.065 31.725 86.850 ;
        RECT 31.745 86.025 35.220 86.935 ;
        RECT 36.115 86.255 40.015 86.935 ;
        RECT 40.025 86.255 49.305 86.935 ;
        RECT 39.085 86.025 40.015 86.255 ;
        RECT 41.385 86.035 42.305 86.255 ;
        RECT 46.970 86.135 49.305 86.255 ;
        RECT 48.385 86.025 49.305 86.135 ;
        RECT 49.880 86.025 53.355 86.935 ;
        RECT 53.510 86.905 53.680 87.125 ;
        RECT 53.960 86.955 54.130 87.175 ;
        RECT 54.285 87.145 59.795 87.955 ;
        RECT 59.805 87.145 65.315 87.955 ;
        RECT 66.440 87.145 69.915 88.055 ;
        RECT 69.935 87.230 70.365 88.015 ;
        RECT 72.665 87.825 73.585 88.045 ;
        RECT 79.665 87.945 80.585 88.055 ;
        RECT 78.250 87.825 80.585 87.945 ;
        RECT 71.305 87.145 80.585 87.825 ;
        RECT 81.160 87.145 84.635 88.055 ;
        RECT 84.840 87.145 88.315 88.055 ;
        RECT 88.325 87.855 89.270 88.055 ;
        RECT 91.085 87.855 92.030 88.055 ;
        RECT 88.325 87.175 91.075 87.855 ;
        RECT 91.085 87.175 93.835 87.855 ;
        RECT 88.325 87.145 89.270 87.175 ;
        RECT 54.425 86.955 54.595 87.145 ;
        RECT 56.275 86.980 56.435 87.090 ;
        RECT 57.645 86.935 57.815 87.125 ;
        RECT 59.945 86.955 60.115 87.145 ;
        RECT 61.320 86.985 61.440 87.095 ;
        RECT 64.545 86.935 64.715 87.125 ;
        RECT 65.475 86.990 65.635 87.100 ;
        RECT 68.225 86.935 68.395 87.125 ;
        RECT 69.600 86.955 69.770 87.145 ;
        RECT 70.535 86.990 70.695 87.100 ;
        RECT 71.445 86.955 71.615 87.145 ;
        RECT 71.900 86.935 72.070 87.125 ;
        RECT 72.365 86.935 72.535 87.125 ;
        RECT 75.125 86.935 75.295 87.125 ;
        RECT 75.580 86.985 75.700 87.095 ;
        RECT 76.320 86.935 76.490 87.125 ;
        RECT 80.185 86.935 80.355 87.125 ;
        RECT 84.320 86.955 84.490 87.145 ;
        RECT 86.620 86.935 86.790 87.125 ;
        RECT 55.170 86.905 56.115 86.935 ;
        RECT 53.365 86.225 56.115 86.905 ;
        RECT 55.170 86.025 56.115 86.225 ;
        RECT 57.055 86.065 57.485 86.850 ;
        RECT 57.505 86.125 61.175 86.935 ;
        RECT 61.645 86.025 64.855 86.935 ;
        RECT 64.960 86.255 68.425 86.935 ;
        RECT 64.960 86.025 65.880 86.255 ;
        RECT 68.740 86.025 72.215 86.935 ;
        RECT 72.225 86.125 74.055 86.935 ;
        RECT 74.065 86.155 75.435 86.935 ;
        RECT 75.905 86.255 79.805 86.935 ;
        RECT 75.905 86.025 76.835 86.255 ;
        RECT 80.045 86.125 82.795 86.935 ;
        RECT 82.815 86.065 83.245 86.850 ;
        RECT 83.460 86.025 86.935 86.935 ;
        RECT 87.090 86.905 87.260 87.125 ;
        RECT 88.000 86.955 88.170 87.145 ;
        RECT 89.845 86.935 90.015 87.125 ;
        RECT 90.760 86.955 90.930 87.175 ;
        RECT 91.085 87.145 92.030 87.175 ;
        RECT 92.600 86.985 92.720 87.095 ;
        RECT 88.750 86.905 89.695 86.935 ;
        RECT 86.945 86.225 89.695 86.905 ;
        RECT 88.750 86.025 89.695 86.225 ;
        RECT 89.705 86.125 92.455 86.935 ;
        RECT 93.070 86.905 93.240 87.125 ;
        RECT 93.520 86.955 93.690 87.175 ;
        RECT 93.845 87.145 95.675 87.955 ;
        RECT 95.695 87.230 96.125 88.015 ;
        RECT 96.145 87.825 97.075 88.055 ;
        RECT 100.485 87.965 101.435 88.055 ;
        RECT 96.145 87.145 100.045 87.825 ;
        RECT 100.485 87.145 102.415 87.965 ;
        RECT 104.405 87.825 105.325 88.045 ;
        RECT 111.405 87.945 112.325 88.055 ;
        RECT 109.990 87.825 112.325 87.945 ;
        RECT 103.045 87.145 112.325 87.825 ;
        RECT 112.715 87.145 114.065 88.055 ;
        RECT 114.085 87.145 115.455 87.925 ;
        RECT 115.475 87.145 116.825 88.055 ;
        RECT 117.305 87.145 118.675 87.955 ;
        RECT 93.985 86.955 94.155 87.145 ;
        RECT 94.730 86.905 95.675 86.935 ;
        RECT 95.830 86.905 96.000 87.125 ;
        RECT 96.560 86.955 96.730 87.145 ;
        RECT 102.265 87.125 102.415 87.145 ;
        RECT 100.425 86.955 100.595 87.125 ;
        RECT 102.265 86.955 102.435 87.125 ;
        RECT 102.720 86.985 102.840 87.095 ;
        RECT 103.185 86.955 103.355 87.145 ;
        RECT 100.425 86.935 100.575 86.955 ;
        RECT 104.290 86.935 104.460 87.125 ;
        RECT 105.025 86.935 105.195 87.125 ;
        RECT 112.570 86.935 112.740 87.125 ;
        RECT 113.305 86.935 113.475 87.125 ;
        RECT 113.765 86.955 113.935 87.145 ;
        RECT 115.145 86.955 115.315 87.145 ;
        RECT 115.605 86.955 115.775 87.145 ;
        RECT 116.980 86.985 117.100 87.095 ;
        RECT 118.365 86.935 118.535 87.145 ;
        RECT 97.490 86.905 98.435 86.935 ;
        RECT 92.925 86.225 95.675 86.905 ;
        RECT 95.685 86.225 98.435 86.905 ;
        RECT 94.730 86.025 95.675 86.225 ;
        RECT 97.490 86.025 98.435 86.225 ;
        RECT 98.645 86.115 100.575 86.935 ;
        RECT 100.975 86.255 104.875 86.935 ;
        RECT 98.645 86.025 99.595 86.115 ;
        RECT 103.945 86.025 104.875 86.255 ;
        RECT 104.885 86.125 108.555 86.935 ;
        RECT 108.575 86.065 109.005 86.850 ;
        RECT 109.255 86.255 113.155 86.935 ;
        RECT 112.225 86.025 113.155 86.255 ;
        RECT 113.165 86.125 116.835 86.935 ;
        RECT 117.305 86.125 118.675 86.935 ;
      LAYER nwell ;
        RECT 5.330 82.905 118.870 85.735 ;
      LAYER pwell ;
        RECT 5.525 81.705 6.895 82.515 ;
        RECT 8.265 82.385 9.185 82.605 ;
        RECT 15.265 82.505 16.185 82.615 ;
        RECT 13.850 82.385 16.185 82.505 ;
        RECT 6.905 81.705 16.185 82.385 ;
        RECT 16.575 81.705 17.925 82.615 ;
        RECT 18.415 81.790 18.845 82.575 ;
        RECT 19.785 81.705 23.260 82.615 ;
        RECT 23.465 81.705 25.295 82.515 ;
        RECT 27.125 82.385 28.045 82.605 ;
        RECT 34.125 82.505 35.045 82.615 ;
        RECT 32.710 82.385 35.045 82.505 ;
        RECT 25.765 81.705 35.045 82.385 ;
        RECT 35.425 81.705 40.935 82.515 ;
        RECT 40.945 81.705 42.775 82.515 ;
        RECT 42.785 81.705 44.155 82.485 ;
        RECT 44.175 81.790 44.605 82.575 ;
        RECT 44.625 82.385 45.555 82.615 ;
        RECT 44.625 81.705 48.525 82.385 ;
        RECT 48.765 81.705 50.135 82.515 ;
        RECT 50.340 81.705 53.815 82.615 ;
        RECT 53.825 81.705 55.655 82.515 ;
        RECT 57.485 82.385 58.405 82.605 ;
        RECT 64.485 82.505 65.405 82.615 ;
        RECT 63.070 82.385 65.405 82.505 ;
        RECT 56.125 81.705 65.405 82.385 ;
        RECT 65.980 81.705 69.455 82.615 ;
        RECT 69.935 81.790 70.365 82.575 ;
        RECT 70.580 81.705 74.055 82.615 ;
        RECT 74.065 81.705 75.895 82.515 ;
        RECT 76.375 81.705 77.725 82.615 ;
        RECT 77.745 81.705 83.255 82.515 ;
        RECT 83.265 81.705 88.775 82.515 ;
        RECT 88.785 81.705 91.535 82.515 ;
        RECT 93.810 82.415 94.755 82.615 ;
        RECT 92.005 81.735 94.755 82.415 ;
        RECT 95.695 81.790 96.125 82.575 ;
        RECT 97.265 82.525 98.215 82.615 ;
        RECT 5.665 81.495 5.835 81.705 ;
        RECT 7.045 81.495 7.215 81.705 ;
        RECT 10.725 81.495 10.895 81.685 ;
        RECT 13.025 81.495 13.195 81.685 ;
        RECT 13.760 81.495 13.930 81.685 ;
        RECT 17.625 81.495 17.795 81.705 ;
        RECT 18.080 81.545 18.200 81.655 ;
        RECT 19.015 81.550 19.175 81.660 ;
        RECT 19.930 81.515 20.100 81.705 ;
        RECT 23.145 81.495 23.315 81.685 ;
        RECT 23.605 81.515 23.775 81.705 ;
        RECT 25.440 81.545 25.560 81.655 ;
        RECT 25.905 81.515 26.075 81.705 ;
        RECT 28.665 81.495 28.835 81.685 ;
        RECT 31.885 81.495 32.055 81.685 ;
        RECT 35.565 81.515 35.735 81.705 ;
        RECT 37.405 81.495 37.575 81.685 ;
        RECT 41.085 81.515 41.255 81.705 ;
        RECT 42.925 81.495 43.095 81.685 ;
        RECT 43.845 81.515 44.015 81.705 ;
        RECT 45.040 81.515 45.210 81.705 ;
        RECT 48.445 81.495 48.615 81.685 ;
        RECT 48.905 81.515 49.075 81.705 ;
        RECT 53.500 81.515 53.670 81.705 ;
        RECT 53.965 81.495 54.135 81.705 ;
        RECT 55.800 81.545 55.920 81.655 ;
        RECT 56.265 81.515 56.435 81.705 ;
        RECT 56.720 81.545 56.840 81.655 ;
        RECT 57.645 81.495 57.815 81.685 ;
        RECT 60.405 81.495 60.575 81.685 ;
        RECT 61.785 81.495 61.955 81.685 ;
        RECT 63.165 81.495 63.335 81.685 ;
        RECT 64.545 81.495 64.715 81.685 ;
        RECT 69.140 81.515 69.310 81.705 ;
        RECT 69.600 81.545 69.720 81.655 ;
        RECT 73.740 81.515 73.910 81.705 ;
        RECT 74.205 81.515 74.375 81.705 ;
        RECT 76.040 81.545 76.160 81.655 ;
        RECT 76.965 81.495 77.135 81.685 ;
        RECT 77.425 81.515 77.595 81.705 ;
        RECT 77.885 81.515 78.055 81.705 ;
        RECT 83.405 81.685 83.575 81.705 ;
        RECT 80.640 81.495 80.810 81.685 ;
        RECT 81.105 81.495 81.275 81.685 ;
        RECT 83.405 81.515 83.580 81.685 ;
        RECT 5.525 80.685 6.895 81.495 ;
        RECT 6.905 80.685 10.575 81.495 ;
        RECT 10.585 80.685 11.955 81.495 ;
        RECT 11.975 80.585 13.325 81.495 ;
        RECT 13.345 80.815 17.245 81.495 ;
        RECT 13.345 80.585 14.275 80.815 ;
        RECT 17.485 80.685 22.995 81.495 ;
        RECT 23.005 80.685 28.515 81.495 ;
        RECT 28.525 80.685 31.275 81.495 ;
        RECT 31.295 80.625 31.725 81.410 ;
        RECT 31.745 80.685 37.255 81.495 ;
        RECT 37.265 80.685 42.775 81.495 ;
        RECT 42.785 80.685 48.295 81.495 ;
        RECT 48.305 80.685 53.815 81.495 ;
        RECT 53.825 80.685 56.575 81.495 ;
        RECT 57.055 80.625 57.485 81.410 ;
        RECT 57.505 80.685 60.255 81.495 ;
        RECT 60.275 80.585 61.625 81.495 ;
        RECT 61.645 80.685 63.015 81.495 ;
        RECT 63.025 80.715 64.395 81.495 ;
        RECT 64.405 80.815 73.595 81.495 ;
        RECT 68.915 80.595 69.845 80.815 ;
        RECT 72.675 80.585 73.595 80.815 ;
        RECT 73.700 80.815 77.165 81.495 ;
        RECT 73.700 80.585 74.620 80.815 ;
        RECT 77.480 80.585 80.955 81.495 ;
        RECT 80.965 80.685 82.795 81.495 ;
        RECT 83.410 81.465 83.580 81.515 ;
        RECT 86.165 81.495 86.335 81.685 ;
        RECT 88.925 81.515 89.095 81.705 ;
        RECT 91.685 81.655 91.855 81.685 ;
        RECT 91.680 81.545 91.855 81.655 ;
        RECT 91.685 81.495 91.855 81.545 ;
        RECT 92.150 81.515 92.320 81.735 ;
        RECT 93.810 81.705 94.755 81.735 ;
        RECT 97.265 81.705 99.195 82.525 ;
        RECT 99.365 81.705 104.875 82.515 ;
        RECT 104.885 81.705 107.635 82.515 ;
        RECT 109.005 82.385 109.925 82.605 ;
        RECT 116.005 82.505 116.925 82.615 ;
        RECT 114.590 82.385 116.925 82.505 ;
        RECT 107.645 81.705 116.925 82.385 ;
        RECT 117.305 81.705 118.675 82.515 ;
        RECT 99.045 81.685 99.195 81.705 ;
        RECT 94.915 81.550 95.075 81.660 ;
        RECT 95.375 81.540 95.535 81.650 ;
        RECT 85.070 81.465 86.015 81.495 ;
        RECT 82.815 80.625 83.245 81.410 ;
        RECT 83.265 80.785 86.015 81.465 ;
        RECT 85.070 80.585 86.015 80.785 ;
        RECT 86.025 80.685 91.535 81.495 ;
        RECT 91.545 80.685 95.215 81.495 ;
        RECT 96.290 81.465 96.460 81.685 ;
        RECT 99.045 81.495 99.215 81.685 ;
        RECT 99.505 81.515 99.675 81.705 ;
        RECT 104.565 81.495 104.735 81.685 ;
        RECT 105.025 81.515 105.195 81.705 ;
        RECT 107.785 81.515 107.955 81.705 ;
        RECT 108.240 81.545 108.360 81.655 ;
        RECT 109.165 81.495 109.335 81.685 ;
        RECT 114.685 81.495 114.855 81.685 ;
        RECT 118.365 81.495 118.535 81.705 ;
        RECT 97.950 81.465 98.895 81.495 ;
        RECT 96.145 80.785 98.895 81.465 ;
        RECT 97.950 80.585 98.895 80.785 ;
        RECT 98.905 80.685 104.415 81.495 ;
        RECT 104.425 80.685 108.095 81.495 ;
        RECT 108.575 80.625 109.005 81.410 ;
        RECT 109.025 80.685 114.535 81.495 ;
        RECT 114.545 80.685 117.295 81.495 ;
        RECT 117.305 80.685 118.675 81.495 ;
      LAYER nwell ;
        RECT 5.330 77.465 118.870 80.295 ;
      LAYER pwell ;
        RECT 5.525 76.265 6.895 77.075 ;
        RECT 6.905 76.265 10.575 77.075 ;
        RECT 10.585 76.265 11.955 77.045 ;
        RECT 12.435 76.265 13.785 77.175 ;
        RECT 13.805 76.945 14.735 77.175 ;
        RECT 13.805 76.265 17.705 76.945 ;
        RECT 18.415 76.350 18.845 77.135 ;
        RECT 19.980 76.265 23.455 77.175 ;
        RECT 23.465 76.975 24.410 77.175 ;
        RECT 23.465 76.295 26.215 76.975 ;
        RECT 23.465 76.265 24.410 76.295 ;
        RECT 5.665 76.055 5.835 76.265 ;
        RECT 7.045 76.215 7.215 76.265 ;
        RECT 7.040 76.105 7.215 76.215 ;
        RECT 7.045 76.075 7.215 76.105 ;
        RECT 7.505 76.055 7.675 76.245 ;
        RECT 11.645 76.075 11.815 76.265 ;
        RECT 12.100 76.105 12.220 76.215 ;
        RECT 13.485 76.075 13.655 76.265 ;
        RECT 14.220 76.075 14.390 76.265 ;
        RECT 17.440 76.055 17.610 76.245 ;
        RECT 18.080 76.105 18.200 76.215 ;
        RECT 19.015 76.110 19.175 76.220 ;
        RECT 21.305 76.055 21.475 76.245 ;
        RECT 23.140 76.075 23.310 76.265 ;
        RECT 25.900 76.075 26.070 76.295 ;
        RECT 26.225 76.265 31.735 77.075 ;
        RECT 31.745 76.265 35.415 77.075 ;
        RECT 35.980 76.945 36.900 77.175 ;
        RECT 35.980 76.265 39.445 76.945 ;
        RECT 39.565 76.265 41.395 77.075 ;
        RECT 41.865 76.265 43.235 77.045 ;
        RECT 44.175 76.350 44.605 77.135 ;
        RECT 44.625 76.945 45.555 77.175 ;
        RECT 44.625 76.265 48.525 76.945 ;
        RECT 48.765 76.265 50.595 77.075 ;
        RECT 51.065 76.975 52.010 77.175 ;
        RECT 51.065 76.295 53.815 76.975 ;
        RECT 51.065 76.265 52.010 76.295 ;
        RECT 26.365 76.245 26.535 76.265 ;
        RECT 26.360 76.075 26.535 76.245 ;
        RECT 26.360 76.055 26.530 76.075 ;
        RECT 5.525 75.245 6.895 76.055 ;
        RECT 7.365 75.375 16.645 76.055 ;
        RECT 8.725 75.155 9.645 75.375 ;
        RECT 14.310 75.255 16.645 75.375 ;
        RECT 15.725 75.145 16.645 75.255 ;
        RECT 17.025 75.375 20.925 76.055 ;
        RECT 17.025 75.145 17.955 75.375 ;
        RECT 21.165 75.245 22.995 76.055 ;
        RECT 23.200 75.145 26.675 76.055 ;
        RECT 26.830 76.025 27.000 76.245 ;
        RECT 29.580 76.105 29.700 76.215 ;
        RECT 30.965 76.055 31.135 76.245 ;
        RECT 31.885 76.075 32.055 76.265 ;
        RECT 33.080 76.055 33.250 76.245 ;
        RECT 35.560 76.105 35.680 76.215 ;
        RECT 37.865 76.055 38.035 76.245 ;
        RECT 38.320 76.105 38.440 76.215 ;
        RECT 38.785 76.055 38.955 76.245 ;
        RECT 39.245 76.075 39.415 76.265 ;
        RECT 39.705 76.075 39.875 76.265 ;
        RECT 41.540 76.105 41.660 76.215 ;
        RECT 42.925 76.075 43.095 76.265 ;
        RECT 43.395 76.110 43.555 76.220 ;
        RECT 45.040 76.075 45.210 76.265 ;
        RECT 48.445 76.055 48.615 76.245 ;
        RECT 48.905 76.075 49.075 76.265 ;
        RECT 53.500 76.245 53.670 76.295 ;
        RECT 53.825 76.265 59.335 77.075 ;
        RECT 59.345 76.265 64.855 77.075 ;
        RECT 65.325 76.945 66.255 77.175 ;
        RECT 65.325 76.265 69.225 76.945 ;
        RECT 69.935 76.350 70.365 77.135 ;
        RECT 70.385 76.265 73.135 77.075 ;
        RECT 73.615 76.265 74.965 77.175 ;
        RECT 74.985 76.265 76.815 77.075 ;
        RECT 80.485 76.945 81.415 77.175 ;
        RECT 82.785 76.945 83.705 77.165 ;
        RECT 89.785 77.065 90.705 77.175 ;
        RECT 88.370 76.945 90.705 77.065 ;
        RECT 77.515 76.265 81.415 76.945 ;
        RECT 81.425 76.265 90.705 76.945 ;
        RECT 91.095 76.265 92.445 77.175 ;
        RECT 92.465 76.265 95.215 77.075 ;
        RECT 95.695 76.350 96.125 77.135 ;
        RECT 96.145 76.265 99.815 77.075 ;
        RECT 99.825 76.265 101.195 77.075 ;
        RECT 102.565 76.945 103.485 77.165 ;
        RECT 109.565 77.065 110.485 77.175 ;
        RECT 108.150 76.945 110.485 77.065 ;
        RECT 101.205 76.265 110.485 76.945 ;
        RECT 110.875 76.265 112.225 77.175 ;
        RECT 112.255 76.265 113.605 77.175 ;
        RECT 113.625 76.265 117.295 77.075 ;
        RECT 117.305 76.265 118.675 77.075 ;
        RECT 50.740 76.105 50.860 76.215 ;
        RECT 53.040 76.055 53.210 76.245 ;
        RECT 53.500 76.075 53.680 76.245 ;
        RECT 53.965 76.075 54.135 76.265 ;
        RECT 53.510 76.055 53.680 76.075 ;
        RECT 57.645 76.055 57.815 76.245 ;
        RECT 59.485 76.075 59.655 76.265 ;
        RECT 60.405 76.055 60.575 76.245 ;
        RECT 60.865 76.055 61.035 76.245 ;
        RECT 62.705 76.055 62.875 76.245 ;
        RECT 65.000 76.105 65.120 76.215 ;
        RECT 65.740 76.075 65.910 76.265 ;
        RECT 68.225 76.055 68.395 76.245 ;
        RECT 69.600 76.105 69.720 76.215 ;
        RECT 69.880 76.055 70.050 76.245 ;
        RECT 70.525 76.075 70.695 76.265 ;
        RECT 73.280 76.105 73.400 76.215 ;
        RECT 73.745 76.055 73.915 76.245 ;
        RECT 74.665 76.075 74.835 76.265 ;
        RECT 75.125 76.075 75.295 76.265 ;
        RECT 76.960 76.105 77.080 76.215 ;
        RECT 79.720 76.055 79.890 76.245 ;
        RECT 80.195 76.100 80.355 76.210 ;
        RECT 80.830 76.075 81.000 76.265 ;
        RECT 81.105 76.055 81.275 76.245 ;
        RECT 81.565 76.075 81.735 76.265 ;
        RECT 82.480 76.105 82.600 76.215 ;
        RECT 28.490 76.025 29.435 76.055 ;
        RECT 26.685 75.345 29.435 76.025 ;
        RECT 28.490 75.145 29.435 75.345 ;
        RECT 29.905 75.275 31.275 76.055 ;
        RECT 31.295 75.185 31.725 75.970 ;
        RECT 32.665 75.375 36.565 76.055 ;
        RECT 32.665 75.145 33.595 75.375 ;
        RECT 36.815 75.145 38.165 76.055 ;
        RECT 38.645 75.375 47.925 76.055 ;
        RECT 40.005 75.155 40.925 75.375 ;
        RECT 45.590 75.255 47.925 75.375 ;
        RECT 47.005 75.145 47.925 75.255 ;
        RECT 48.305 75.245 49.675 76.055 ;
        RECT 49.880 75.145 53.355 76.055 ;
        RECT 53.365 75.145 56.840 76.055 ;
        RECT 57.055 75.185 57.485 75.970 ;
        RECT 57.505 75.245 58.875 76.055 ;
        RECT 58.885 75.375 60.715 76.055 ;
        RECT 60.725 75.375 62.555 76.055 ;
        RECT 58.885 75.145 60.230 75.375 ;
        RECT 61.210 75.145 62.555 75.375 ;
        RECT 62.565 75.245 68.075 76.055 ;
        RECT 68.085 75.245 69.455 76.055 ;
        RECT 69.465 75.375 73.365 76.055 ;
        RECT 69.465 75.145 70.395 75.375 ;
        RECT 73.605 75.245 76.355 76.055 ;
        RECT 76.560 75.145 80.035 76.055 ;
        RECT 80.965 75.275 82.335 76.055 ;
        RECT 83.265 76.025 84.210 76.055 ;
        RECT 85.700 76.025 85.870 76.245 ;
        RECT 86.165 76.055 86.335 76.245 ;
        RECT 89.840 76.105 89.960 76.215 ;
        RECT 92.145 76.075 92.315 76.265 ;
        RECT 92.605 76.075 92.775 76.265 ;
        RECT 93.520 76.055 93.690 76.245 ;
        RECT 93.990 76.055 94.160 76.245 ;
        RECT 95.360 76.105 95.480 76.215 ;
        RECT 96.285 76.075 96.455 76.265 ;
        RECT 97.665 76.055 97.835 76.245 ;
        RECT 99.500 76.105 99.620 76.215 ;
        RECT 99.965 76.075 100.135 76.265 ;
        RECT 101.345 76.075 101.515 76.265 ;
        RECT 103.370 76.055 103.540 76.245 ;
        RECT 105.025 76.055 105.195 76.245 ;
        RECT 105.485 76.055 105.655 76.245 ;
        RECT 107.325 76.055 107.495 76.245 ;
        RECT 109.440 76.055 109.610 76.245 ;
        RECT 111.925 76.075 112.095 76.265 ;
        RECT 113.305 76.055 113.475 76.265 ;
        RECT 113.765 76.075 113.935 76.265 ;
        RECT 116.980 76.105 117.100 76.215 ;
        RECT 118.365 76.055 118.535 76.265 ;
        RECT 82.815 75.185 83.245 75.970 ;
        RECT 83.265 75.345 86.015 76.025 ;
        RECT 83.265 75.145 84.210 75.345 ;
        RECT 86.025 75.245 89.695 76.055 ;
        RECT 90.360 75.145 93.835 76.055 ;
        RECT 93.845 75.145 97.320 76.055 ;
        RECT 97.525 75.245 99.355 76.055 ;
        RECT 100.055 75.375 103.955 76.055 ;
        RECT 103.025 75.145 103.955 75.375 ;
        RECT 103.965 75.275 105.335 76.055 ;
        RECT 105.345 75.245 107.175 76.055 ;
        RECT 107.185 75.275 108.555 76.055 ;
        RECT 108.575 75.185 109.005 75.970 ;
        RECT 109.025 75.375 112.925 76.055 ;
        RECT 109.025 75.145 109.955 75.375 ;
        RECT 113.165 75.245 116.835 76.055 ;
        RECT 117.305 75.245 118.675 76.055 ;
      LAYER nwell ;
        RECT 5.330 72.025 118.870 74.855 ;
      LAYER pwell ;
        RECT 5.525 70.825 6.895 71.635 ;
        RECT 6.905 70.825 8.275 71.635 ;
        RECT 12.795 71.505 13.725 71.725 ;
        RECT 16.555 71.505 17.475 71.735 ;
        RECT 8.285 70.825 17.475 71.505 ;
        RECT 18.415 70.910 18.845 71.695 ;
        RECT 18.960 71.505 19.880 71.735 ;
        RECT 18.960 70.825 22.425 71.505 ;
        RECT 22.740 70.825 26.215 71.735 ;
        RECT 26.225 70.825 27.595 71.635 ;
        RECT 32.115 71.505 33.045 71.725 ;
        RECT 35.875 71.505 36.795 71.735 ;
        RECT 27.605 70.825 36.795 71.505 ;
        RECT 36.805 70.825 38.635 71.635 ;
        RECT 38.655 70.825 40.005 71.735 ;
        RECT 40.025 70.825 41.395 71.605 ;
        RECT 42.335 70.825 43.685 71.735 ;
        RECT 44.175 70.910 44.605 71.695 ;
        RECT 44.625 71.505 45.555 71.735 ;
        RECT 44.625 70.825 48.525 71.505 ;
        RECT 48.765 70.825 52.435 71.635 ;
        RECT 54.710 71.535 55.655 71.735 ;
        RECT 52.905 70.855 55.655 71.535 ;
        RECT 62.590 71.505 63.935 71.735 ;
        RECT 5.665 70.615 5.835 70.825 ;
        RECT 7.045 70.615 7.215 70.825 ;
        RECT 8.425 70.635 8.595 70.825 ;
        RECT 10.735 70.660 10.895 70.770 ;
        RECT 12.565 70.615 12.735 70.805 ;
        RECT 13.020 70.665 13.140 70.775 ;
        RECT 13.485 70.615 13.655 70.805 ;
        RECT 14.865 70.615 15.035 70.805 ;
        RECT 17.635 70.670 17.795 70.780 ;
        RECT 20.380 70.665 20.500 70.775 ;
        RECT 22.225 70.635 22.395 70.825 ;
        RECT 24.060 70.615 24.230 70.805 ;
        RECT 25.900 70.635 26.070 70.825 ;
        RECT 26.365 70.635 26.535 70.825 ;
        RECT 27.745 70.805 27.915 70.825 ;
        RECT 27.740 70.635 27.915 70.805 ;
        RECT 27.740 70.615 27.910 70.635 ;
        RECT 5.525 69.805 6.895 70.615 ;
        RECT 6.905 69.805 10.575 70.615 ;
        RECT 11.505 69.835 12.875 70.615 ;
        RECT 13.355 69.705 14.705 70.615 ;
        RECT 14.725 69.805 20.235 70.615 ;
        RECT 20.900 69.705 24.375 70.615 ;
        RECT 24.580 69.705 28.055 70.615 ;
        RECT 28.210 70.585 28.380 70.805 ;
        RECT 30.960 70.665 31.080 70.775 ;
        RECT 31.885 70.615 32.055 70.805 ;
        RECT 36.945 70.635 37.115 70.825 ;
        RECT 37.405 70.615 37.575 70.805 ;
        RECT 38.785 70.635 38.955 70.825 ;
        RECT 41.085 70.635 41.255 70.825 ;
        RECT 41.555 70.670 41.715 70.780 ;
        RECT 42.465 70.635 42.635 70.825 ;
        RECT 43.840 70.665 43.960 70.775 ;
        RECT 45.040 70.635 45.210 70.825 ;
        RECT 47.065 70.615 47.235 70.805 ;
        RECT 48.905 70.635 49.075 70.825 ;
        RECT 52.585 70.775 52.755 70.805 ;
        RECT 52.580 70.665 52.755 70.775 ;
        RECT 52.585 70.615 52.755 70.665 ;
        RECT 53.050 70.635 53.220 70.855 ;
        RECT 54.710 70.825 55.655 70.855 ;
        RECT 55.675 70.825 58.415 71.505 ;
        RECT 59.345 70.825 62.085 71.505 ;
        RECT 62.105 70.825 63.935 71.505 ;
        RECT 63.945 71.505 65.290 71.735 ;
        RECT 63.945 70.825 65.775 71.505 ;
        RECT 65.785 70.825 67.615 71.635 ;
        RECT 68.085 70.825 69.455 71.605 ;
        RECT 69.935 70.910 70.365 71.695 ;
        RECT 70.385 70.825 71.755 71.605 ;
        RECT 72.225 71.505 73.155 71.735 ;
        RECT 72.225 70.825 76.125 71.505 ;
        RECT 76.365 70.825 78.195 71.635 ;
        RECT 78.400 70.825 81.875 71.735 ;
        RECT 81.885 71.535 82.830 71.735 ;
        RECT 81.885 70.855 84.635 71.535 ;
        RECT 81.885 70.825 82.830 70.855 ;
        RECT 56.275 70.660 56.435 70.770 ;
        RECT 58.105 70.635 58.275 70.825 ;
        RECT 58.575 70.670 58.735 70.780 ;
        RECT 59.485 70.635 59.655 70.825 ;
        RECT 59.945 70.615 60.115 70.805 ;
        RECT 61.785 70.615 61.955 70.805 ;
        RECT 62.245 70.615 62.415 70.825 ;
        RECT 65.000 70.665 65.120 70.775 ;
        RECT 65.465 70.615 65.635 70.825 ;
        RECT 65.925 70.635 66.095 70.825 ;
        RECT 67.760 70.665 67.880 70.775 ;
        RECT 69.145 70.635 69.315 70.825 ;
        RECT 69.600 70.665 69.720 70.775 ;
        RECT 70.525 70.635 70.695 70.825 ;
        RECT 71.900 70.665 72.020 70.775 ;
        RECT 72.640 70.635 72.810 70.825 ;
        RECT 76.045 70.615 76.215 70.805 ;
        RECT 76.505 70.615 76.675 70.825 ;
        RECT 81.560 70.635 81.730 70.825 ;
        RECT 82.035 70.660 82.195 70.770 ;
        RECT 83.405 70.615 83.575 70.805 ;
        RECT 84.320 70.635 84.490 70.855 ;
        RECT 84.645 70.825 88.315 71.635 ;
        RECT 88.520 70.825 91.995 71.735 ;
        RECT 92.005 70.825 95.675 71.635 ;
        RECT 95.695 70.910 96.125 71.695 ;
        RECT 96.145 70.825 97.515 71.605 ;
        RECT 97.525 70.825 98.895 71.635 ;
        RECT 98.915 70.825 100.265 71.735 ;
        RECT 100.285 70.825 105.795 71.635 ;
        RECT 105.805 70.825 107.175 71.635 ;
        RECT 108.545 71.505 109.465 71.725 ;
        RECT 115.545 71.625 116.465 71.735 ;
        RECT 114.130 71.505 116.465 71.625 ;
        RECT 107.185 70.825 116.465 71.505 ;
        RECT 117.305 70.825 118.675 71.635 ;
        RECT 84.785 70.635 84.955 70.825 ;
        RECT 88.925 70.615 89.095 70.805 ;
        RECT 91.680 70.635 91.850 70.825 ;
        RECT 92.145 70.635 92.315 70.825 ;
        RECT 93.520 70.615 93.690 70.805 ;
        RECT 93.985 70.615 94.155 70.805 ;
        RECT 97.205 70.635 97.375 70.825 ;
        RECT 97.665 70.635 97.835 70.825 ;
        RECT 99.965 70.635 100.135 70.825 ;
        RECT 100.425 70.635 100.595 70.825 ;
        RECT 103.645 70.615 103.815 70.805 ;
        RECT 105.945 70.635 106.115 70.825 ;
        RECT 107.325 70.615 107.495 70.825 ;
        RECT 109.440 70.615 109.610 70.805 ;
        RECT 113.305 70.615 113.475 70.805 ;
        RECT 116.980 70.665 117.100 70.775 ;
        RECT 118.365 70.615 118.535 70.825 ;
        RECT 29.870 70.585 30.815 70.615 ;
        RECT 28.065 69.905 30.815 70.585 ;
        RECT 29.870 69.705 30.815 69.905 ;
        RECT 31.295 69.745 31.725 70.530 ;
        RECT 31.745 69.805 37.255 70.615 ;
        RECT 37.265 69.935 46.545 70.615 ;
        RECT 38.625 69.715 39.545 69.935 ;
        RECT 44.210 69.815 46.545 69.935 ;
        RECT 45.625 69.705 46.545 69.815 ;
        RECT 46.925 69.805 52.435 70.615 ;
        RECT 52.445 69.805 56.115 70.615 ;
        RECT 57.055 69.745 57.485 70.530 ;
        RECT 57.535 69.705 60.255 70.615 ;
        RECT 60.265 69.935 62.095 70.615 ;
        RECT 60.265 69.705 61.610 69.935 ;
        RECT 62.105 69.805 64.855 70.615 ;
        RECT 65.325 69.935 74.605 70.615 ;
        RECT 66.685 69.715 67.605 69.935 ;
        RECT 72.270 69.815 74.605 69.935 ;
        RECT 73.685 69.705 74.605 69.815 ;
        RECT 74.995 69.705 76.345 70.615 ;
        RECT 76.365 69.805 81.875 70.615 ;
        RECT 82.815 69.745 83.245 70.530 ;
        RECT 83.265 69.805 88.775 70.615 ;
        RECT 88.785 69.805 90.155 70.615 ;
        RECT 90.360 69.705 93.835 70.615 ;
        RECT 93.845 69.935 103.125 70.615 ;
        RECT 95.205 69.715 96.125 69.935 ;
        RECT 100.790 69.815 103.125 69.935 ;
        RECT 102.205 69.705 103.125 69.815 ;
        RECT 103.505 69.805 107.175 70.615 ;
        RECT 107.185 69.805 108.555 70.615 ;
        RECT 108.575 69.745 109.005 70.530 ;
        RECT 109.025 69.935 112.925 70.615 ;
        RECT 109.025 69.705 109.955 69.935 ;
        RECT 113.165 69.805 116.835 70.615 ;
        RECT 117.305 69.805 118.675 70.615 ;
      LAYER nwell ;
        RECT 5.330 66.585 118.870 69.415 ;
      LAYER pwell ;
        RECT 5.525 65.385 6.895 66.195 ;
        RECT 6.905 65.385 12.415 66.195 ;
        RECT 12.425 65.385 14.255 66.195 ;
        RECT 14.405 65.385 17.015 66.295 ;
        RECT 17.025 65.385 18.395 66.195 ;
        RECT 18.415 65.470 18.845 66.255 ;
        RECT 18.865 65.385 22.535 66.195 ;
        RECT 22.545 65.385 26.020 66.295 ;
        RECT 26.420 65.385 29.895 66.295 ;
        RECT 29.905 65.385 31.735 66.195 ;
        RECT 32.205 65.385 35.680 66.295 ;
        RECT 35.885 65.385 41.395 66.195 ;
        RECT 41.405 65.385 44.155 66.195 ;
        RECT 44.175 65.470 44.605 66.255 ;
        RECT 44.625 65.385 48.295 66.195 ;
        RECT 49.420 65.385 52.895 66.295 ;
        RECT 53.100 65.385 56.575 66.295 ;
        RECT 56.585 65.385 58.415 66.195 ;
        RECT 58.425 65.385 67.530 66.065 ;
        RECT 67.625 65.385 69.455 66.195 ;
        RECT 69.935 65.470 70.365 66.255 ;
        RECT 71.745 66.065 72.665 66.285 ;
        RECT 78.745 66.185 79.665 66.295 ;
        RECT 77.330 66.065 79.665 66.185 ;
        RECT 70.385 65.385 79.665 66.065 ;
        RECT 80.045 65.385 81.875 66.195 ;
        RECT 82.540 65.385 86.015 66.295 ;
        RECT 86.220 65.385 89.695 66.295 ;
        RECT 89.900 65.385 93.375 66.295 ;
        RECT 93.385 65.385 95.215 66.195 ;
        RECT 95.695 65.470 96.125 66.255 ;
        RECT 96.145 66.065 97.075 66.295 ;
        RECT 96.145 65.385 100.045 66.065 ;
        RECT 100.285 65.385 103.955 66.195 ;
        RECT 103.965 65.385 105.335 66.195 ;
        RECT 105.345 65.385 106.715 66.165 ;
        RECT 108.085 66.065 109.005 66.285 ;
        RECT 115.085 66.185 116.005 66.295 ;
        RECT 113.670 66.065 116.005 66.185 ;
        RECT 106.725 65.385 116.005 66.065 ;
        RECT 117.305 65.385 118.675 66.195 ;
        RECT 5.665 65.175 5.835 65.385 ;
        RECT 7.045 65.175 7.215 65.385 ;
        RECT 12.565 65.195 12.735 65.385 ;
        RECT 16.700 65.365 16.870 65.385 ;
        RECT 16.700 65.195 16.875 65.365 ;
        RECT 16.705 65.175 16.875 65.195 ;
        RECT 17.165 65.175 17.335 65.385 ;
        RECT 19.005 65.195 19.175 65.385 ;
        RECT 20.855 65.220 21.015 65.330 ;
        RECT 22.690 65.195 22.860 65.385 ;
        RECT 24.980 65.175 25.150 65.365 ;
        RECT 25.455 65.220 25.615 65.330 ;
        RECT 27.285 65.175 27.455 65.365 ;
        RECT 27.745 65.175 27.915 65.365 ;
        RECT 29.125 65.175 29.295 65.365 ;
        RECT 29.580 65.195 29.750 65.385 ;
        RECT 30.045 65.195 30.215 65.385 ;
        RECT 30.960 65.225 31.080 65.335 ;
        RECT 31.880 65.225 32.000 65.335 ;
        RECT 32.350 65.195 32.520 65.385 ;
        RECT 33.265 65.175 33.435 65.365 ;
        RECT 33.725 65.175 33.895 65.365 ;
        RECT 36.025 65.195 36.195 65.385 ;
        RECT 36.485 65.175 36.655 65.365 ;
        RECT 36.945 65.175 37.115 65.365 ;
        RECT 38.780 65.225 38.900 65.335 ;
        RECT 40.165 65.175 40.335 65.365 ;
        RECT 40.625 65.175 40.795 65.365 ;
        RECT 41.545 65.195 41.715 65.385 ;
        RECT 42.460 65.225 42.580 65.335 ;
        RECT 42.925 65.175 43.095 65.365 ;
        RECT 44.765 65.195 44.935 65.385 ;
        RECT 48.455 65.230 48.615 65.340 ;
        RECT 52.580 65.195 52.750 65.385 ;
        RECT 53.050 65.175 53.220 65.365 ;
        RECT 56.260 65.195 56.430 65.385 ;
        RECT 56.725 65.335 56.895 65.385 ;
        RECT 56.720 65.225 56.895 65.335 ;
        RECT 56.725 65.195 56.895 65.225 ;
        RECT 57.650 65.175 57.820 65.365 ;
        RECT 58.565 65.195 58.735 65.385 ;
        RECT 62.705 65.175 62.875 65.365 ;
        RECT 64.545 65.175 64.715 65.365 ;
        RECT 65.005 65.175 65.175 65.365 ;
        RECT 67.765 65.195 67.935 65.385 ;
        RECT 68.680 65.225 68.800 65.335 ;
        RECT 69.150 65.175 69.320 65.365 ;
        RECT 69.600 65.225 69.720 65.335 ;
        RECT 70.525 65.195 70.695 65.385 ;
        RECT 71.905 65.175 72.075 65.365 ;
        RECT 73.285 65.175 73.455 65.365 ;
        RECT 78.800 65.225 78.920 65.335 ;
        RECT 80.185 65.195 80.355 65.385 ;
        RECT 82.020 65.225 82.140 65.335 ;
        RECT 82.480 65.175 82.650 65.365 ;
        RECT 85.700 65.195 85.870 65.385 ;
        RECT 86.625 65.175 86.795 65.365 ;
        RECT 87.090 65.175 87.260 65.365 ;
        RECT 89.380 65.195 89.550 65.385 ;
        RECT 90.770 65.175 90.940 65.365 ;
        RECT 93.060 65.195 93.230 65.385 ;
        RECT 93.525 65.195 93.695 65.385 ;
        RECT 94.445 65.175 94.615 65.365 ;
        RECT 95.360 65.225 95.480 65.335 ;
        RECT 96.560 65.195 96.730 65.385 ;
        RECT 100.425 65.195 100.595 65.385 ;
        RECT 101.345 65.175 101.515 65.365 ;
        RECT 104.105 65.195 104.275 65.385 ;
        RECT 105.025 65.175 105.195 65.365 ;
        RECT 105.485 65.175 105.655 65.385 ;
        RECT 106.865 65.195 107.035 65.385 ;
        RECT 108.245 65.175 108.415 65.365 ;
        RECT 109.440 65.175 109.610 65.365 ;
        RECT 114.225 65.175 114.395 65.365 ;
        RECT 114.685 65.175 114.855 65.365 ;
        RECT 116.065 65.175 116.235 65.365 ;
        RECT 116.535 65.230 116.695 65.340 ;
        RECT 118.365 65.175 118.535 65.385 ;
        RECT 5.525 64.365 6.895 65.175 ;
        RECT 6.905 64.365 12.415 65.175 ;
        RECT 13.440 64.495 16.905 65.175 ;
        RECT 13.440 64.265 14.360 64.495 ;
        RECT 17.025 64.365 20.695 65.175 ;
        RECT 21.820 64.265 25.295 65.175 ;
        RECT 26.225 64.395 27.595 65.175 ;
        RECT 27.605 64.395 28.975 65.175 ;
        RECT 28.985 64.365 30.815 65.175 ;
        RECT 31.295 64.305 31.725 65.090 ;
        RECT 32.215 64.265 33.565 65.175 ;
        RECT 33.585 64.365 35.415 65.175 ;
        RECT 35.425 64.395 36.795 65.175 ;
        RECT 36.805 64.365 38.635 65.175 ;
        RECT 39.115 64.265 40.465 65.175 ;
        RECT 40.485 64.365 42.315 65.175 ;
        RECT 42.785 64.495 52.065 65.175 ;
        RECT 44.145 64.275 45.065 64.495 ;
        RECT 49.730 64.375 52.065 64.495 ;
        RECT 51.145 64.265 52.065 64.375 ;
        RECT 52.905 64.265 56.380 65.175 ;
        RECT 57.055 64.305 57.485 65.090 ;
        RECT 57.505 64.265 60.980 65.175 ;
        RECT 61.185 64.495 63.015 65.175 ;
        RECT 63.025 64.495 64.855 65.175 ;
        RECT 61.185 64.265 62.530 64.495 ;
        RECT 63.025 64.265 64.370 64.495 ;
        RECT 64.865 64.365 68.535 65.175 ;
        RECT 69.005 64.265 71.615 65.175 ;
        RECT 71.775 64.265 73.125 65.175 ;
        RECT 73.145 64.365 78.655 65.175 ;
        RECT 79.320 64.265 82.795 65.175 ;
        RECT 82.815 64.305 83.245 65.090 ;
        RECT 83.360 64.495 86.825 65.175 ;
        RECT 83.360 64.265 84.280 64.495 ;
        RECT 86.945 64.265 90.420 65.175 ;
        RECT 90.625 64.265 94.100 65.175 ;
        RECT 94.305 64.365 97.975 65.175 ;
        RECT 98.080 64.495 101.545 65.175 ;
        RECT 101.760 64.495 105.225 65.175 ;
        RECT 98.080 64.265 99.000 64.495 ;
        RECT 101.760 64.265 102.680 64.495 ;
        RECT 105.345 64.365 107.175 65.175 ;
        RECT 107.185 64.395 108.555 65.175 ;
        RECT 108.575 64.305 109.005 65.090 ;
        RECT 109.025 64.495 112.925 65.175 ;
        RECT 109.025 64.265 109.955 64.495 ;
        RECT 113.175 64.265 114.525 65.175 ;
        RECT 114.555 64.265 115.905 65.175 ;
        RECT 115.925 64.365 117.295 65.175 ;
        RECT 117.305 64.365 118.675 65.175 ;
      LAYER nwell ;
        RECT 5.330 61.145 118.870 63.975 ;
      LAYER pwell ;
        RECT 5.525 59.945 6.895 60.755 ;
        RECT 6.905 59.945 10.575 60.755 ;
        RECT 11.045 59.945 12.415 60.725 ;
        RECT 12.895 59.945 14.245 60.855 ;
        RECT 14.265 60.625 15.195 60.855 ;
        RECT 14.265 59.945 18.165 60.625 ;
        RECT 18.415 60.030 18.845 60.815 ;
        RECT 18.865 60.625 19.795 60.855 ;
        RECT 23.100 60.625 24.020 60.855 ;
        RECT 27.240 60.625 28.160 60.855 ;
        RECT 18.865 59.945 22.765 60.625 ;
        RECT 23.100 59.945 26.565 60.625 ;
        RECT 27.240 59.945 30.705 60.625 ;
        RECT 30.875 59.945 34.035 60.855 ;
        RECT 35.405 60.625 36.325 60.845 ;
        RECT 42.405 60.745 43.325 60.855 ;
        RECT 40.990 60.625 43.325 60.745 ;
        RECT 34.045 59.945 43.325 60.625 ;
        RECT 44.175 60.030 44.605 60.815 ;
        RECT 45.545 59.945 46.915 60.725 ;
        RECT 46.925 60.625 47.855 60.855 ;
        RECT 46.925 59.945 50.825 60.625 ;
        RECT 51.075 59.945 52.425 60.855 ;
        RECT 52.445 59.945 57.955 60.755 ;
        RECT 57.965 59.945 60.715 60.755 ;
        RECT 61.185 60.625 62.530 60.855 ;
        RECT 63.025 60.625 64.370 60.855 ;
        RECT 65.350 60.625 66.695 60.855 ;
        RECT 67.190 60.625 68.535 60.855 ;
        RECT 61.185 59.945 63.015 60.625 ;
        RECT 63.025 59.945 64.855 60.625 ;
        RECT 64.865 59.945 66.695 60.625 ;
        RECT 66.705 59.945 68.535 60.625 ;
        RECT 68.545 59.945 69.915 60.755 ;
        RECT 69.935 60.030 70.365 60.815 ;
        RECT 70.385 59.945 72.215 60.755 ;
        RECT 72.225 59.945 73.595 60.725 ;
        RECT 73.605 59.945 75.435 60.755 ;
        RECT 75.905 60.625 76.835 60.855 ;
        RECT 83.245 60.625 84.175 60.855 ;
        RECT 75.905 59.945 79.805 60.625 ;
        RECT 80.275 59.945 84.175 60.625 ;
        RECT 84.185 59.945 85.555 60.725 ;
        RECT 88.765 60.625 89.695 60.855 ;
        RECT 85.795 59.945 89.695 60.625 ;
        RECT 89.800 60.625 90.720 60.855 ;
        RECT 89.800 59.945 93.265 60.625 ;
        RECT 93.385 59.945 95.215 60.755 ;
        RECT 95.695 60.030 96.125 60.815 ;
        RECT 99.345 60.625 100.275 60.855 ;
        RECT 96.375 59.945 100.275 60.625 ;
        RECT 100.285 59.945 101.655 60.755 ;
        RECT 104.865 60.625 105.795 60.855 ;
        RECT 107.165 60.625 108.085 60.845 ;
        RECT 114.165 60.745 115.085 60.855 ;
        RECT 112.750 60.625 115.085 60.745 ;
        RECT 101.895 59.945 105.795 60.625 ;
        RECT 105.805 59.945 115.085 60.625 ;
        RECT 115.465 59.945 117.295 60.755 ;
        RECT 117.305 59.945 118.675 60.755 ;
        RECT 5.665 59.735 5.835 59.945 ;
        RECT 7.045 59.735 7.215 59.945 ;
        RECT 8.880 59.785 9.000 59.895 ;
        RECT 9.345 59.735 9.515 59.925 ;
        RECT 10.725 59.895 10.895 59.925 ;
        RECT 10.720 59.785 10.895 59.895 ;
        RECT 10.725 59.735 10.895 59.785 ;
        RECT 12.105 59.755 12.275 59.945 ;
        RECT 12.560 59.785 12.680 59.895 ;
        RECT 13.945 59.755 14.115 59.945 ;
        RECT 14.680 59.755 14.850 59.945 ;
        RECT 19.280 59.755 19.450 59.945 ;
        RECT 19.930 59.735 20.100 59.925 ;
        RECT 26.090 59.735 26.260 59.925 ;
        RECT 26.365 59.755 26.535 59.945 ;
        RECT 26.820 59.785 26.940 59.895 ;
        RECT 27.560 59.735 27.730 59.925 ;
        RECT 30.505 59.755 30.675 59.945 ;
        RECT 30.965 59.755 31.135 59.945 ;
        RECT 31.885 59.735 32.055 59.925 ;
        RECT 34.185 59.755 34.355 59.945 ;
        RECT 41.085 59.735 41.255 59.925 ;
        RECT 43.840 59.785 43.960 59.895 ;
        RECT 44.775 59.790 44.935 59.900 ;
        RECT 46.605 59.755 46.775 59.945 ;
        RECT 47.340 59.755 47.510 59.945 ;
        RECT 47.525 59.735 47.695 59.925 ;
        RECT 47.985 59.735 48.155 59.925 ;
        RECT 50.745 59.735 50.915 59.925 ;
        RECT 51.205 59.755 51.375 59.945 ;
        RECT 51.480 59.735 51.650 59.925 ;
        RECT 52.585 59.755 52.755 59.945 ;
        RECT 55.345 59.735 55.515 59.925 ;
        RECT 57.645 59.735 57.815 59.925 ;
        RECT 58.105 59.755 58.275 59.945 ;
        RECT 60.860 59.785 60.980 59.895 ;
        RECT 62.705 59.755 62.875 59.945 ;
        RECT 63.160 59.785 63.280 59.895 ;
        RECT 63.625 59.735 63.795 59.925 ;
        RECT 64.545 59.755 64.715 59.945 ;
        RECT 65.005 59.755 65.175 59.945 ;
        RECT 66.390 59.735 66.560 59.925 ;
        RECT 66.845 59.755 67.015 59.945 ;
        RECT 68.685 59.755 68.855 59.945 ;
        RECT 69.145 59.735 69.315 59.925 ;
        RECT 70.525 59.755 70.695 59.945 ;
        RECT 73.285 59.755 73.455 59.945 ;
        RECT 73.745 59.755 73.915 59.945 ;
        RECT 75.580 59.785 75.700 59.895 ;
        RECT 76.320 59.755 76.490 59.945 ;
        RECT 79.265 59.735 79.435 59.925 ;
        RECT 79.725 59.735 79.895 59.925 ;
        RECT 81.565 59.735 81.735 59.925 ;
        RECT 83.590 59.755 83.760 59.945 ;
        RECT 84.325 59.755 84.495 59.945 ;
        RECT 86.625 59.735 86.795 59.925 ;
        RECT 87.095 59.780 87.255 59.890 ;
        RECT 88.005 59.735 88.175 59.925 ;
        RECT 89.110 59.755 89.280 59.945 ;
        RECT 93.065 59.755 93.235 59.945 ;
        RECT 93.525 59.755 93.695 59.945 ;
        RECT 95.360 59.785 95.480 59.895 ;
        RECT 99.690 59.755 99.860 59.945 ;
        RECT 100.425 59.755 100.595 59.945 ;
        RECT 105.210 59.755 105.380 59.945 ;
        RECT 105.945 59.735 106.115 59.945 ;
        RECT 106.405 59.735 106.575 59.925 ;
        RECT 107.795 59.780 107.955 59.890 ;
        RECT 109.165 59.735 109.335 59.925 ;
        RECT 114.685 59.735 114.855 59.925 ;
        RECT 115.605 59.755 115.775 59.945 ;
        RECT 118.365 59.735 118.535 59.945 ;
        RECT 5.525 58.925 6.895 59.735 ;
        RECT 6.905 58.925 8.735 59.735 ;
        RECT 9.205 58.955 10.575 59.735 ;
        RECT 10.585 59.055 19.775 59.735 ;
        RECT 15.095 58.835 16.025 59.055 ;
        RECT 18.855 58.825 19.775 59.055 ;
        RECT 19.785 58.825 22.395 59.735 ;
        RECT 22.775 59.055 26.675 59.735 ;
        RECT 25.745 58.825 26.675 59.055 ;
        RECT 27.145 59.055 31.045 59.735 ;
        RECT 27.145 58.825 28.075 59.055 ;
        RECT 31.295 58.865 31.725 59.650 ;
        RECT 31.745 59.055 40.850 59.735 ;
        RECT 40.945 58.925 46.455 59.735 ;
        RECT 46.465 58.955 47.835 59.735 ;
        RECT 47.845 58.925 49.675 59.735 ;
        RECT 49.685 58.955 51.055 59.735 ;
        RECT 51.065 59.055 54.965 59.735 ;
        RECT 51.065 58.825 51.995 59.055 ;
        RECT 55.205 58.925 57.035 59.735 ;
        RECT 57.055 58.865 57.485 59.650 ;
        RECT 57.505 58.925 63.015 59.735 ;
        RECT 63.485 59.055 66.225 59.735 ;
        RECT 66.245 58.825 68.855 59.735 ;
        RECT 69.005 59.055 78.195 59.735 ;
        RECT 73.515 58.835 74.445 59.055 ;
        RECT 77.275 58.825 78.195 59.055 ;
        RECT 78.205 58.955 79.575 59.735 ;
        RECT 79.585 58.925 81.415 59.735 ;
        RECT 81.435 58.825 82.785 59.735 ;
        RECT 82.815 58.865 83.245 59.650 ;
        RECT 83.360 59.055 86.825 59.735 ;
        RECT 87.865 59.055 97.055 59.735 ;
        RECT 83.360 58.825 84.280 59.055 ;
        RECT 92.375 58.835 93.305 59.055 ;
        RECT 96.135 58.825 97.055 59.055 ;
        RECT 97.065 59.055 106.255 59.735 ;
        RECT 97.065 58.825 97.985 59.055 ;
        RECT 100.815 58.835 101.745 59.055 ;
        RECT 106.265 58.955 107.635 59.735 ;
        RECT 108.575 58.865 109.005 59.650 ;
        RECT 109.025 58.925 114.535 59.735 ;
        RECT 114.545 58.925 117.295 59.735 ;
        RECT 117.305 58.925 118.675 59.735 ;
      LAYER nwell ;
        RECT 5.330 55.705 118.870 58.535 ;
      LAYER pwell ;
        RECT 5.525 54.505 6.895 55.315 ;
        RECT 6.905 54.505 8.275 55.315 ;
        RECT 12.795 55.185 13.725 55.405 ;
        RECT 16.555 55.185 17.475 55.415 ;
        RECT 8.285 54.505 17.475 55.185 ;
        RECT 18.415 54.590 18.845 55.375 ;
        RECT 18.960 55.185 19.880 55.415 ;
        RECT 22.640 55.185 23.560 55.415 ;
        RECT 27.585 55.185 28.505 55.405 ;
        RECT 34.585 55.305 35.505 55.415 ;
        RECT 33.170 55.185 35.505 55.305 ;
        RECT 18.960 54.505 22.425 55.185 ;
        RECT 22.640 54.505 26.105 55.185 ;
        RECT 26.225 54.505 35.505 55.185 ;
        RECT 35.885 55.185 36.815 55.415 ;
        RECT 35.885 54.505 39.785 55.185 ;
        RECT 40.025 54.505 43.695 55.315 ;
        RECT 44.175 54.590 44.605 55.375 ;
        RECT 45.555 54.505 46.905 55.415 ;
        RECT 46.935 54.505 48.285 55.415 ;
        RECT 49.665 55.185 50.585 55.405 ;
        RECT 56.665 55.305 57.585 55.415 ;
        RECT 55.250 55.185 57.585 55.305 ;
        RECT 48.305 54.505 57.585 55.185 ;
        RECT 57.965 54.505 59.795 55.315 ;
        RECT 59.835 54.505 62.555 55.415 ;
        RECT 62.575 54.505 65.315 55.185 ;
        RECT 65.325 54.505 68.065 55.185 ;
        RECT 68.085 54.505 69.915 55.315 ;
        RECT 69.935 54.590 70.365 55.375 ;
        RECT 70.385 54.505 72.995 55.415 ;
        RECT 73.615 54.505 74.965 55.415 ;
        RECT 74.985 54.505 76.815 55.315 ;
        RECT 81.335 55.185 82.265 55.405 ;
        RECT 85.095 55.185 86.015 55.415 ;
        RECT 89.600 55.185 90.520 55.415 ;
        RECT 76.825 54.505 86.015 55.185 ;
        RECT 87.055 54.505 90.520 55.185 ;
        RECT 90.720 55.185 91.640 55.415 ;
        RECT 90.720 54.505 94.185 55.185 ;
        RECT 94.315 54.505 95.665 55.415 ;
        RECT 95.695 54.590 96.125 55.375 ;
        RECT 96.195 54.505 99.355 55.415 ;
        RECT 99.365 54.505 100.735 55.285 ;
        RECT 100.745 55.185 101.665 55.415 ;
        RECT 104.495 55.185 105.425 55.405 ;
        RECT 100.745 54.505 109.935 55.185 ;
        RECT 109.945 54.505 115.455 55.315 ;
        RECT 115.465 54.505 117.295 55.315 ;
        RECT 117.305 54.505 118.675 55.315 ;
        RECT 5.665 54.295 5.835 54.505 ;
        RECT 7.045 54.295 7.215 54.505 ;
        RECT 8.425 54.315 8.595 54.505 ;
        RECT 9.805 54.295 9.975 54.485 ;
        RECT 12.565 54.295 12.735 54.485 ;
        RECT 13.025 54.295 13.195 54.485 ;
        RECT 17.635 54.350 17.795 54.460 ;
        RECT 20.110 54.295 20.280 54.485 ;
        RECT 20.840 54.345 20.960 54.455 ;
        RECT 21.305 54.295 21.475 54.485 ;
        RECT 22.225 54.315 22.395 54.505 ;
        RECT 25.905 54.315 26.075 54.505 ;
        RECT 26.365 54.315 26.535 54.505 ;
        RECT 30.515 54.340 30.675 54.450 ;
        RECT 31.885 54.295 32.055 54.485 ;
        RECT 35.560 54.345 35.680 54.455 ;
        RECT 36.300 54.315 36.470 54.505 ;
        RECT 36.945 54.295 37.115 54.485 ;
        RECT 37.400 54.345 37.520 54.455 ;
        RECT 38.140 54.295 38.310 54.485 ;
        RECT 40.165 54.315 40.335 54.505 ;
        RECT 42.005 54.295 42.175 54.485 ;
        RECT 43.385 54.295 43.555 54.485 ;
        RECT 43.840 54.345 43.960 54.455 ;
        RECT 44.775 54.350 44.935 54.460 ;
        RECT 45.685 54.315 45.855 54.505 ;
        RECT 47.065 54.315 47.235 54.505 ;
        RECT 48.445 54.315 48.615 54.505 ;
        RECT 53.320 54.295 53.490 54.485 ;
        RECT 57.645 54.295 57.815 54.485 ;
        RECT 58.105 54.315 58.275 54.505 ;
        RECT 61.325 54.295 61.495 54.485 ;
        RECT 62.245 54.315 62.415 54.505 ;
        RECT 63.165 54.295 63.335 54.485 ;
        RECT 65.005 54.295 65.175 54.505 ;
        RECT 65.465 54.315 65.635 54.505 ;
        RECT 68.225 54.315 68.395 54.505 ;
        RECT 70.530 54.485 70.700 54.505 ;
        RECT 70.525 54.315 70.700 54.485 ;
        RECT 73.280 54.345 73.400 54.455 ;
        RECT 73.745 54.315 73.915 54.505 ;
        RECT 75.125 54.315 75.295 54.505 ;
        RECT 70.525 54.295 70.695 54.315 ;
        RECT 76.045 54.295 76.215 54.485 ;
        RECT 76.965 54.315 77.135 54.505 ;
        RECT 81.565 54.295 81.735 54.485 ;
        RECT 83.405 54.295 83.575 54.485 ;
        RECT 86.175 54.350 86.335 54.460 ;
        RECT 87.085 54.315 87.255 54.505 ;
        RECT 88.925 54.295 89.095 54.485 ;
        RECT 93.985 54.315 94.155 54.505 ;
        RECT 95.365 54.315 95.535 54.505 ;
        RECT 96.285 54.315 96.455 54.505 ;
        RECT 98.125 54.295 98.295 54.485 ;
        RECT 99.505 54.295 99.675 54.505 ;
        RECT 100.885 54.295 101.055 54.485 ;
        RECT 104.560 54.345 104.680 54.455 ;
        RECT 105.945 54.295 106.115 54.485 ;
        RECT 106.405 54.295 106.575 54.485 ;
        RECT 108.240 54.345 108.360 54.455 ;
        RECT 109.165 54.295 109.335 54.485 ;
        RECT 109.625 54.315 109.795 54.505 ;
        RECT 110.085 54.315 110.255 54.505 ;
        RECT 114.685 54.295 114.855 54.485 ;
        RECT 115.605 54.315 115.775 54.505 ;
        RECT 118.365 54.295 118.535 54.505 ;
        RECT 5.525 53.485 6.895 54.295 ;
        RECT 6.905 53.485 9.655 54.295 ;
        RECT 9.665 53.615 11.495 54.295 ;
        RECT 11.505 53.515 12.875 54.295 ;
        RECT 12.995 53.615 16.460 54.295 ;
        RECT 16.795 53.615 20.695 54.295 ;
        RECT 21.165 53.615 30.355 54.295 ;
        RECT 15.540 53.385 16.460 53.615 ;
        RECT 19.765 53.385 20.695 53.615 ;
        RECT 25.675 53.395 26.605 53.615 ;
        RECT 29.435 53.385 30.355 53.615 ;
        RECT 31.295 53.425 31.725 54.210 ;
        RECT 31.745 53.485 35.415 54.295 ;
        RECT 35.885 53.515 37.255 54.295 ;
        RECT 37.725 53.615 41.625 54.295 ;
        RECT 37.725 53.385 38.655 53.615 ;
        RECT 41.865 53.485 43.235 54.295 ;
        RECT 43.245 53.615 52.525 54.295 ;
        RECT 44.605 53.395 45.525 53.615 ;
        RECT 50.190 53.495 52.525 53.615 ;
        RECT 51.605 53.385 52.525 53.495 ;
        RECT 52.905 53.615 56.805 54.295 ;
        RECT 52.905 53.385 53.835 53.615 ;
        RECT 57.055 53.425 57.485 54.210 ;
        RECT 57.505 53.485 61.175 54.295 ;
        RECT 61.185 53.615 63.015 54.295 ;
        RECT 63.025 53.615 64.855 54.295 ;
        RECT 61.670 53.385 63.015 53.615 ;
        RECT 63.510 53.385 64.855 53.615 ;
        RECT 64.865 53.485 70.375 54.295 ;
        RECT 70.385 53.485 75.895 54.295 ;
        RECT 75.905 53.485 81.415 54.295 ;
        RECT 81.425 53.485 82.795 54.295 ;
        RECT 82.815 53.425 83.245 54.210 ;
        RECT 83.265 53.485 88.775 54.295 ;
        RECT 88.785 53.615 97.890 54.295 ;
        RECT 97.985 53.485 99.355 54.295 ;
        RECT 99.375 53.385 100.725 54.295 ;
        RECT 100.745 53.485 104.415 54.295 ;
        RECT 104.895 53.385 106.245 54.295 ;
        RECT 106.265 53.485 108.095 54.295 ;
        RECT 108.575 53.425 109.005 54.210 ;
        RECT 109.025 53.485 114.535 54.295 ;
        RECT 114.545 53.485 117.295 54.295 ;
        RECT 117.305 53.485 118.675 54.295 ;
      LAYER nwell ;
        RECT 5.330 50.265 118.870 53.095 ;
      LAYER pwell ;
        RECT 5.525 49.065 6.895 49.875 ;
        RECT 6.905 49.065 8.275 49.875 ;
        RECT 12.795 49.745 13.725 49.965 ;
        RECT 16.555 49.745 17.475 49.975 ;
        RECT 8.285 49.065 17.475 49.745 ;
        RECT 18.415 49.150 18.845 49.935 ;
        RECT 18.875 49.065 20.225 49.975 ;
        RECT 20.245 49.065 21.615 49.875 ;
        RECT 21.625 49.065 25.100 49.975 ;
        RECT 25.315 49.065 26.665 49.975 ;
        RECT 26.685 49.065 32.195 49.875 ;
        RECT 37.635 49.745 38.565 49.965 ;
        RECT 41.395 49.745 42.315 49.975 ;
        RECT 33.125 49.065 42.315 49.745 ;
        RECT 42.335 49.065 43.685 49.975 ;
        RECT 44.175 49.150 44.605 49.935 ;
        RECT 44.720 49.745 45.640 49.975 ;
        RECT 44.720 49.065 48.185 49.745 ;
        RECT 48.445 49.065 51.055 49.975 ;
        RECT 51.065 49.065 56.575 49.875 ;
        RECT 56.585 49.065 62.095 49.875 ;
        RECT 62.105 49.065 67.615 49.875 ;
        RECT 67.625 49.065 69.455 49.875 ;
        RECT 69.935 49.150 70.365 49.935 ;
        RECT 70.385 49.065 71.755 49.845 ;
        RECT 71.775 49.065 73.125 49.975 ;
        RECT 73.145 49.065 76.815 49.875 ;
        RECT 76.825 49.065 78.195 49.875 ;
        RECT 78.400 49.065 81.875 49.975 ;
        RECT 82.080 49.065 85.555 49.975 ;
        RECT 85.760 49.065 89.235 49.975 ;
        RECT 90.165 49.065 91.535 49.845 ;
        RECT 92.200 49.065 95.675 49.975 ;
        RECT 95.695 49.150 96.125 49.935 ;
        RECT 96.145 49.065 101.655 49.875 ;
        RECT 101.665 49.065 107.175 49.875 ;
        RECT 107.185 49.065 112.695 49.875 ;
        RECT 112.705 49.065 116.375 49.875 ;
        RECT 117.305 49.065 118.675 49.875 ;
        RECT 5.665 48.855 5.835 49.065 ;
        RECT 7.045 48.855 7.215 49.065 ;
        RECT 8.425 48.875 8.595 49.065 ;
        RECT 12.565 48.855 12.735 49.045 ;
        RECT 14.865 48.855 15.035 49.045 ;
        RECT 15.325 48.855 15.495 49.045 ;
        RECT 17.635 48.910 17.795 49.020 ;
        RECT 19.925 48.875 20.095 49.065 ;
        RECT 20.385 48.875 20.555 49.065 ;
        RECT 20.845 48.855 21.015 49.045 ;
        RECT 21.770 48.875 21.940 49.065 ;
        RECT 25.445 49.045 25.615 49.065 ;
        RECT 25.440 48.875 25.615 49.045 ;
        RECT 25.440 48.855 25.610 48.875 ;
        RECT 25.910 48.855 26.080 49.045 ;
        RECT 26.825 48.875 26.995 49.065 ;
        RECT 29.585 48.855 29.755 49.045 ;
        RECT 31.885 48.855 32.055 49.045 ;
        RECT 32.355 48.910 32.515 49.020 ;
        RECT 33.265 48.875 33.435 49.065 ;
        RECT 37.405 48.855 37.575 49.045 ;
        RECT 42.925 48.855 43.095 49.045 ;
        RECT 43.385 48.875 43.555 49.065 ;
        RECT 43.840 48.905 43.960 49.015 ;
        RECT 47.985 48.875 48.155 49.065 ;
        RECT 48.440 48.905 48.560 49.015 ;
        RECT 50.740 48.875 50.910 49.065 ;
        RECT 51.205 48.875 51.375 49.065 ;
        RECT 52.120 48.855 52.290 49.045 ;
        RECT 52.585 48.855 52.755 49.045 ;
        RECT 56.275 48.900 56.435 49.010 ;
        RECT 56.725 48.875 56.895 49.065 ;
        RECT 57.645 48.855 57.815 49.045 ;
        RECT 60.405 48.855 60.575 49.045 ;
        RECT 62.245 48.875 62.415 49.065 ;
        RECT 64.540 48.855 64.710 49.045 ;
        RECT 65.005 48.855 65.175 49.045 ;
        RECT 66.845 48.855 67.015 49.045 ;
        RECT 67.765 48.875 67.935 49.065 ;
        RECT 69.600 48.905 69.720 49.015 ;
        RECT 71.445 48.875 71.615 49.065 ;
        RECT 71.905 48.875 72.075 49.065 ;
        RECT 73.285 48.875 73.455 49.065 ;
        RECT 76.320 48.855 76.490 49.045 ;
        RECT 76.965 48.875 77.135 49.065 ;
        RECT 80.185 48.855 80.355 49.045 ;
        RECT 81.560 48.875 81.730 49.065 ;
        RECT 85.240 48.875 85.410 49.065 ;
        RECT 86.625 48.855 86.795 49.045 ;
        RECT 87.090 48.855 87.260 49.045 ;
        RECT 88.920 48.875 89.090 49.065 ;
        RECT 89.395 48.910 89.555 49.020 ;
        RECT 90.305 48.875 90.475 49.065 ;
        RECT 91.680 48.905 91.800 49.015 ;
        RECT 93.980 48.855 94.150 49.045 ;
        RECT 94.450 48.855 94.620 49.045 ;
        RECT 95.360 48.875 95.530 49.065 ;
        RECT 96.285 48.875 96.455 49.065 ;
        RECT 98.120 48.905 98.240 49.015 ;
        RECT 101.805 48.875 101.975 49.065 ;
        RECT 101.990 48.855 102.160 49.045 ;
        RECT 105.945 48.855 106.115 49.045 ;
        RECT 106.405 48.855 106.575 49.045 ;
        RECT 107.325 48.875 107.495 49.065 ;
        RECT 107.795 48.900 107.955 49.010 ;
        RECT 109.165 48.855 109.335 49.045 ;
        RECT 112.845 48.875 113.015 49.065 ;
        RECT 114.685 48.855 114.855 49.045 ;
        RECT 116.535 48.910 116.695 49.020 ;
        RECT 118.365 48.855 118.535 49.065 ;
        RECT 5.525 48.045 6.895 48.855 ;
        RECT 6.905 48.045 12.415 48.855 ;
        RECT 12.425 48.045 13.795 48.855 ;
        RECT 13.815 47.945 15.165 48.855 ;
        RECT 15.185 48.045 20.695 48.855 ;
        RECT 20.705 48.045 22.075 48.855 ;
        RECT 22.280 47.945 25.755 48.855 ;
        RECT 25.765 47.945 29.240 48.855 ;
        RECT 29.445 48.045 31.275 48.855 ;
        RECT 31.295 47.985 31.725 48.770 ;
        RECT 31.745 48.045 37.255 48.855 ;
        RECT 37.265 48.045 42.775 48.855 ;
        RECT 42.785 48.045 48.295 48.855 ;
        RECT 48.960 47.945 52.435 48.855 ;
        RECT 52.445 48.045 56.115 48.855 ;
        RECT 57.055 47.985 57.485 48.770 ;
        RECT 57.505 48.045 60.255 48.855 ;
        RECT 60.265 48.175 62.095 48.855 ;
        RECT 60.750 47.945 62.095 48.175 ;
        RECT 62.245 47.945 64.855 48.855 ;
        RECT 64.865 48.045 66.695 48.855 ;
        RECT 66.705 48.175 75.895 48.855 ;
        RECT 71.215 47.955 72.145 48.175 ;
        RECT 74.975 47.945 75.895 48.175 ;
        RECT 75.905 48.175 79.805 48.855 ;
        RECT 75.905 47.945 76.835 48.175 ;
        RECT 80.045 48.045 82.795 48.855 ;
        RECT 82.815 47.985 83.245 48.770 ;
        RECT 83.360 48.175 86.825 48.855 ;
        RECT 83.360 47.945 84.280 48.175 ;
        RECT 86.945 47.945 90.420 48.855 ;
        RECT 90.820 47.945 94.295 48.855 ;
        RECT 94.305 47.945 97.780 48.855 ;
        RECT 98.675 48.175 102.575 48.855 ;
        RECT 101.645 47.945 102.575 48.175 ;
        RECT 102.680 48.175 106.145 48.855 ;
        RECT 102.680 47.945 103.600 48.175 ;
        RECT 106.265 48.075 107.635 48.855 ;
        RECT 108.575 47.985 109.005 48.770 ;
        RECT 109.025 48.045 114.535 48.855 ;
        RECT 114.545 48.045 117.295 48.855 ;
        RECT 117.305 48.045 118.675 48.855 ;
      LAYER nwell ;
        RECT 5.330 44.825 118.870 47.655 ;
      LAYER pwell ;
        RECT 5.525 43.625 6.895 44.435 ;
        RECT 6.905 43.625 12.415 44.435 ;
        RECT 12.425 43.625 15.175 44.435 ;
        RECT 15.185 43.625 16.555 44.405 ;
        RECT 16.565 43.625 18.395 44.435 ;
        RECT 18.415 43.710 18.845 44.495 ;
        RECT 18.865 44.305 19.795 44.535 ;
        RECT 18.865 43.625 22.765 44.305 ;
        RECT 23.005 43.625 24.835 44.435 ;
        RECT 25.040 43.625 28.515 44.535 ;
        RECT 28.525 43.625 29.895 44.435 ;
        RECT 29.905 43.625 31.275 44.405 ;
        RECT 31.285 43.625 34.760 44.535 ;
        RECT 34.965 43.625 40.475 44.435 ;
        RECT 40.485 43.625 44.155 44.435 ;
        RECT 44.175 43.710 44.605 44.495 ;
        RECT 44.720 44.305 45.640 44.535 ;
        RECT 44.720 43.625 48.185 44.305 ;
        RECT 48.305 43.625 49.675 44.435 ;
        RECT 49.880 43.625 53.355 44.535 ;
        RECT 53.365 43.625 56.840 44.535 ;
        RECT 57.505 43.625 60.225 44.535 ;
        RECT 60.265 44.305 61.610 44.535 ;
        RECT 62.105 44.305 63.450 44.535 ;
        RECT 64.430 44.305 65.775 44.535 ;
        RECT 60.265 43.625 62.095 44.305 ;
        RECT 62.105 43.625 63.935 44.305 ;
        RECT 63.945 43.625 65.775 44.305 ;
        RECT 65.785 43.625 68.535 44.435 ;
        RECT 68.545 43.625 69.915 44.405 ;
        RECT 69.935 43.710 70.365 44.495 ;
        RECT 74.895 44.305 75.825 44.525 ;
        RECT 78.655 44.305 79.575 44.535 ;
        RECT 70.385 43.625 79.575 44.305 ;
        RECT 79.680 44.305 80.600 44.535 ;
        RECT 79.680 43.625 83.145 44.305 ;
        RECT 83.265 43.625 86.740 44.535 ;
        RECT 87.040 44.305 87.960 44.535 ;
        RECT 91.545 44.305 92.475 44.535 ;
        RECT 87.040 43.625 90.505 44.305 ;
        RECT 91.545 43.625 95.445 44.305 ;
        RECT 95.695 43.710 96.125 44.495 ;
        RECT 100.655 44.305 101.585 44.525 ;
        RECT 104.415 44.305 105.335 44.535 ;
        RECT 96.145 43.625 105.335 44.305 ;
        RECT 105.355 43.625 106.705 44.535 ;
        RECT 106.735 43.625 108.085 44.535 ;
        RECT 108.105 43.625 113.615 44.435 ;
        RECT 113.625 43.625 117.295 44.435 ;
        RECT 117.305 43.625 118.675 44.435 ;
        RECT 5.665 43.415 5.835 43.625 ;
        RECT 7.045 43.415 7.215 43.625 ;
        RECT 9.800 43.465 9.920 43.575 ;
        RECT 11.185 43.415 11.355 43.605 ;
        RECT 12.565 43.415 12.735 43.625 ;
        RECT 13.025 43.415 13.195 43.605 ;
        RECT 16.245 43.435 16.415 43.625 ;
        RECT 16.705 43.435 16.875 43.625 ;
        RECT 19.280 43.435 19.450 43.625 ;
        RECT 23.145 43.415 23.315 43.625 ;
        RECT 23.600 43.465 23.720 43.575 ;
        RECT 24.065 43.415 24.235 43.605 ;
        RECT 27.745 43.415 27.915 43.605 ;
        RECT 28.200 43.435 28.370 43.625 ;
        RECT 28.665 43.435 28.835 43.625 ;
        RECT 30.045 43.435 30.215 43.625 ;
        RECT 31.430 43.435 31.600 43.625 ;
        RECT 31.885 43.415 32.055 43.605 ;
        RECT 35.105 43.435 35.275 43.625 ;
        RECT 40.625 43.435 40.795 43.625 ;
        RECT 42.005 43.415 42.175 43.605 ;
        RECT 42.465 43.415 42.635 43.605 ;
        RECT 44.120 43.415 44.290 43.605 ;
        RECT 47.985 43.415 48.155 43.625 ;
        RECT 48.445 43.435 48.615 43.625 ;
        RECT 49.830 43.415 50.000 43.605 ;
        RECT 53.040 43.435 53.210 43.625 ;
        RECT 53.510 43.435 53.680 43.625 ;
        RECT 56.725 43.415 56.895 43.605 ;
        RECT 57.180 43.465 57.300 43.575 ;
        RECT 57.645 43.435 57.815 43.625 ;
        RECT 61.325 43.435 61.495 43.605 ;
        RECT 61.785 43.435 61.955 43.625 ;
        RECT 63.625 43.435 63.795 43.625 ;
        RECT 61.325 43.415 61.395 43.435 ;
        RECT 64.085 43.415 64.255 43.625 ;
        RECT 64.545 43.415 64.715 43.605 ;
        RECT 65.925 43.435 66.095 43.625 ;
        RECT 67.305 43.415 67.475 43.605 ;
        RECT 67.765 43.415 67.935 43.605 ;
        RECT 68.685 43.435 68.855 43.625 ;
        RECT 70.525 43.415 70.695 43.625 ;
        RECT 76.690 43.415 76.860 43.605 ;
        RECT 77.425 43.415 77.595 43.605 ;
        RECT 82.485 43.415 82.655 43.605 ;
        RECT 82.945 43.435 83.115 43.625 ;
        RECT 83.410 43.435 83.580 43.625 ;
        RECT 83.680 43.415 83.850 43.605 ;
        RECT 90.305 43.435 90.475 43.625 ;
        RECT 90.760 43.580 90.930 43.605 ;
        RECT 90.760 43.470 90.935 43.580 ;
        RECT 90.760 43.415 90.930 43.470 ;
        RECT 91.220 43.465 91.340 43.575 ;
        RECT 91.960 43.435 92.130 43.625 ;
        RECT 94.900 43.415 95.070 43.605 ;
        RECT 95.360 43.465 95.480 43.575 ;
        RECT 95.825 43.415 95.995 43.605 ;
        RECT 96.285 43.435 96.455 43.625 ;
        RECT 106.405 43.435 106.575 43.625 ;
        RECT 106.865 43.435 107.035 43.625 ;
        RECT 108.245 43.415 108.415 43.625 ;
        RECT 109.165 43.415 109.335 43.605 ;
        RECT 113.765 43.435 113.935 43.625 ;
        RECT 114.685 43.415 114.855 43.605 ;
        RECT 118.365 43.415 118.535 43.625 ;
        RECT 5.525 42.605 6.895 43.415 ;
        RECT 6.905 42.605 9.655 43.415 ;
        RECT 10.125 42.635 11.495 43.415 ;
        RECT 11.515 42.505 12.865 43.415 ;
        RECT 12.885 42.735 22.075 43.415 ;
        RECT 17.395 42.515 18.325 42.735 ;
        RECT 21.155 42.505 22.075 42.735 ;
        RECT 22.095 42.505 23.445 43.415 ;
        RECT 24.035 42.735 27.500 43.415 ;
        RECT 27.715 42.735 31.180 43.415 ;
        RECT 26.580 42.505 27.500 42.735 ;
        RECT 30.260 42.505 31.180 42.735 ;
        RECT 31.295 42.545 31.725 43.330 ;
        RECT 31.745 42.735 40.935 43.415 ;
        RECT 36.255 42.515 37.185 42.735 ;
        RECT 40.015 42.505 40.935 42.735 ;
        RECT 40.955 42.505 42.305 43.415 ;
        RECT 42.325 42.635 43.695 43.415 ;
        RECT 43.705 42.735 47.605 43.415 ;
        RECT 43.705 42.505 44.635 42.735 ;
        RECT 47.845 42.605 49.675 43.415 ;
        RECT 49.685 42.505 53.160 43.415 ;
        RECT 53.460 42.735 56.925 43.415 ;
        RECT 53.460 42.505 54.380 42.735 ;
        RECT 57.055 42.545 57.485 43.330 ;
        RECT 59.125 43.185 61.395 43.415 ;
        RECT 58.640 42.505 61.395 43.185 ;
        RECT 61.655 42.735 64.395 43.415 ;
        RECT 64.405 42.735 66.235 43.415 ;
        RECT 64.890 42.505 66.235 42.735 ;
        RECT 66.255 42.505 67.605 43.415 ;
        RECT 67.625 42.605 70.375 43.415 ;
        RECT 70.385 42.735 73.125 43.415 ;
        RECT 73.375 42.735 77.275 43.415 ;
        RECT 76.345 42.505 77.275 42.735 ;
        RECT 77.285 42.605 79.115 43.415 ;
        RECT 79.220 42.735 82.685 43.415 ;
        RECT 79.220 42.505 80.140 42.735 ;
        RECT 82.815 42.545 83.245 43.330 ;
        RECT 83.265 42.735 87.165 43.415 ;
        RECT 83.265 42.505 84.195 42.735 ;
        RECT 87.600 42.505 91.075 43.415 ;
        RECT 91.740 42.505 95.215 43.415 ;
        RECT 95.795 42.735 99.260 43.415 ;
        RECT 98.340 42.505 99.260 42.735 ;
        RECT 99.365 42.735 108.555 43.415 ;
        RECT 99.365 42.505 100.285 42.735 ;
        RECT 103.115 42.515 104.045 42.735 ;
        RECT 108.575 42.545 109.005 43.330 ;
        RECT 109.025 42.605 114.535 43.415 ;
        RECT 114.545 42.605 117.295 43.415 ;
        RECT 117.305 42.605 118.675 43.415 ;
      LAYER nwell ;
        RECT 5.330 39.385 118.870 42.215 ;
      LAYER pwell ;
        RECT 5.525 38.185 6.895 38.995 ;
        RECT 6.905 38.185 8.275 38.995 ;
        RECT 12.795 38.865 13.725 39.085 ;
        RECT 16.555 38.865 17.475 39.095 ;
        RECT 8.285 38.185 17.475 38.865 ;
        RECT 18.415 38.270 18.845 39.055 ;
        RECT 18.865 38.865 19.795 39.095 ;
        RECT 18.865 38.185 22.765 38.865 ;
        RECT 23.200 38.185 26.675 39.095 ;
        RECT 26.685 38.865 27.615 39.095 ;
        RECT 26.685 38.185 30.585 38.865 ;
        RECT 30.825 38.185 33.575 38.995 ;
        RECT 33.585 38.865 34.515 39.095 ;
        RECT 33.585 38.185 37.485 38.865 ;
        RECT 37.725 38.185 41.395 38.995 ;
        RECT 41.405 38.185 42.775 38.995 ;
        RECT 42.795 38.185 44.145 39.095 ;
        RECT 44.175 38.270 44.605 39.055 ;
        RECT 49.135 38.865 50.065 39.085 ;
        RECT 52.895 38.865 53.815 39.095 ;
        RECT 44.625 38.185 53.815 38.865 ;
        RECT 54.985 38.415 57.740 39.095 ;
        RECT 58.110 38.415 63.475 39.095 ;
        RECT 63.700 38.415 66.455 39.095 ;
        RECT 54.985 38.185 57.255 38.415 ;
        RECT 59.050 38.185 63.475 38.415 ;
        RECT 64.185 38.185 66.455 38.415 ;
        RECT 66.705 38.185 69.455 38.995 ;
        RECT 69.935 38.270 70.365 39.055 ;
        RECT 70.385 38.185 72.215 38.995 ;
        RECT 72.695 38.185 74.045 39.095 ;
        RECT 74.065 38.185 76.815 38.995 ;
        RECT 77.335 38.185 80.495 39.095 ;
        RECT 80.505 38.185 81.875 38.965 ;
        RECT 81.885 38.185 83.255 38.965 ;
        RECT 83.265 38.185 84.635 38.965 ;
        RECT 84.740 38.865 85.660 39.095 ;
        RECT 88.420 38.865 89.340 39.095 ;
        RECT 92.100 38.865 93.020 39.095 ;
        RECT 84.740 38.185 88.205 38.865 ;
        RECT 88.420 38.185 91.885 38.865 ;
        RECT 92.100 38.185 95.565 38.865 ;
        RECT 95.695 38.270 96.125 39.055 ;
        RECT 96.145 38.185 97.975 38.995 ;
        RECT 101.645 38.865 102.575 39.095 ;
        RECT 98.675 38.185 102.575 38.865 ;
        RECT 102.680 38.865 103.600 39.095 ;
        RECT 108.920 38.865 109.840 39.095 ;
        RECT 102.680 38.185 106.145 38.865 ;
        RECT 106.375 38.185 109.840 38.865 ;
        RECT 109.945 38.185 111.315 38.965 ;
        RECT 111.325 38.185 116.835 38.995 ;
        RECT 117.305 38.185 118.675 38.995 ;
        RECT 5.665 37.975 5.835 38.185 ;
        RECT 7.045 37.975 7.215 38.185 ;
        RECT 8.425 37.995 8.595 38.185 ;
        RECT 12.565 37.975 12.735 38.165 ;
        RECT 17.635 38.030 17.795 38.140 ;
        RECT 18.085 37.975 18.255 38.165 ;
        RECT 19.280 37.995 19.450 38.185 ;
        RECT 26.360 38.165 26.530 38.185 ;
        RECT 22.685 37.975 22.855 38.165 ;
        RECT 26.360 37.995 26.535 38.165 ;
        RECT 26.820 38.025 26.940 38.135 ;
        RECT 27.100 37.995 27.270 38.185 ;
        RECT 26.365 37.975 26.535 37.995 ;
        RECT 27.285 37.975 27.455 38.165 ;
        RECT 30.965 38.135 31.135 38.185 ;
        RECT 30.960 38.025 31.135 38.135 ;
        RECT 30.965 37.995 31.135 38.025 ;
        RECT 32.805 37.975 32.975 38.165 ;
        RECT 34.000 37.995 34.170 38.185 ;
        RECT 34.185 37.975 34.355 38.165 ;
        RECT 34.655 38.020 34.815 38.130 ;
        RECT 37.865 37.995 38.035 38.185 ;
        RECT 38.785 37.975 38.955 38.165 ;
        RECT 39.245 37.975 39.415 38.165 ;
        RECT 41.545 37.995 41.715 38.185 ;
        RECT 42.925 37.995 43.095 38.185 ;
        RECT 44.765 37.995 44.935 38.185 ;
        RECT 54.985 38.165 55.055 38.185 ;
        RECT 45.040 37.975 45.210 38.165 ;
        RECT 48.905 37.975 49.075 38.165 ;
        RECT 53.975 38.030 54.135 38.140 ;
        RECT 54.425 37.975 54.595 38.165 ;
        RECT 54.885 37.995 55.055 38.165 ;
        RECT 57.645 37.975 57.815 38.165 ;
        RECT 62.245 37.975 62.415 38.165 ;
        RECT 63.165 37.995 63.335 38.185 ;
        RECT 66.385 38.165 66.455 38.185 ;
        RECT 66.385 37.995 66.555 38.165 ;
        RECT 66.845 37.995 67.015 38.185 ;
        RECT 67.765 37.975 67.935 38.165 ;
        RECT 69.600 38.025 69.720 38.135 ;
        RECT 70.525 37.995 70.695 38.185 ;
        RECT 72.360 38.025 72.480 38.135 ;
        RECT 72.825 37.995 72.995 38.185 ;
        RECT 73.280 38.025 73.400 38.135 ;
        RECT 73.745 37.975 73.915 38.165 ;
        RECT 74.205 37.995 74.375 38.185 ;
        RECT 76.960 38.025 77.080 38.135 ;
        RECT 77.425 37.995 77.595 38.185 ;
        RECT 81.565 37.995 81.735 38.185 ;
        RECT 82.025 37.995 82.195 38.185 ;
        RECT 83.405 37.995 83.575 38.185 ;
        RECT 84.325 37.975 84.495 38.165 ;
        RECT 84.780 38.025 84.900 38.135 ;
        RECT 88.005 37.995 88.175 38.185 ;
        RECT 88.650 37.975 88.820 38.165 ;
        RECT 89.660 37.975 89.830 38.165 ;
        RECT 91.685 37.995 91.855 38.185 ;
        RECT 94.445 37.975 94.615 38.165 ;
        RECT 94.905 37.975 95.075 38.165 ;
        RECT 95.365 37.995 95.535 38.185 ;
        RECT 96.285 37.995 96.455 38.185 ;
        RECT 98.125 38.135 98.295 38.165 ;
        RECT 97.660 38.025 97.780 38.135 ;
        RECT 98.120 38.025 98.295 38.135 ;
        RECT 98.125 37.975 98.295 38.025 ;
        RECT 101.990 37.995 102.160 38.185 ;
        RECT 105.945 37.995 106.115 38.185 ;
        RECT 106.405 37.995 106.575 38.185 ;
        RECT 107.325 37.975 107.495 38.165 ;
        RECT 109.165 37.975 109.335 38.165 ;
        RECT 111.005 37.995 111.175 38.185 ;
        RECT 111.465 37.995 111.635 38.185 ;
        RECT 114.685 37.975 114.855 38.165 ;
        RECT 116.980 38.025 117.100 38.135 ;
        RECT 118.365 37.975 118.535 38.185 ;
        RECT 5.525 37.165 6.895 37.975 ;
        RECT 6.905 37.165 12.415 37.975 ;
        RECT 12.425 37.165 17.935 37.975 ;
        RECT 17.945 37.165 19.315 37.975 ;
        RECT 19.420 37.295 22.885 37.975 ;
        RECT 23.100 37.295 26.565 37.975 ;
        RECT 27.255 37.295 30.720 37.975 ;
        RECT 19.420 37.065 20.340 37.295 ;
        RECT 23.100 37.065 24.020 37.295 ;
        RECT 29.800 37.065 30.720 37.295 ;
        RECT 31.295 37.105 31.725 37.890 ;
        RECT 31.755 37.065 33.105 37.975 ;
        RECT 33.125 37.195 34.495 37.975 ;
        RECT 35.520 37.295 38.985 37.975 ;
        RECT 35.520 37.065 36.440 37.295 ;
        RECT 39.105 37.165 44.615 37.975 ;
        RECT 44.625 37.295 48.525 37.975 ;
        RECT 44.625 37.065 45.555 37.295 ;
        RECT 48.765 37.165 54.275 37.975 ;
        RECT 54.285 37.165 57.035 37.975 ;
        RECT 57.055 37.105 57.485 37.890 ;
        RECT 57.505 37.745 59.075 37.975 ;
        RECT 61.165 37.935 62.085 37.975 ;
        RECT 61.165 37.745 62.095 37.935 ;
        RECT 57.505 37.385 62.095 37.745 ;
        RECT 57.505 37.295 62.085 37.385 ;
        RECT 59.085 37.065 62.085 37.295 ;
        RECT 62.105 37.165 67.615 37.975 ;
        RECT 67.625 37.165 73.135 37.975 ;
        RECT 73.605 37.295 82.795 37.975 ;
        RECT 78.115 37.075 79.045 37.295 ;
        RECT 81.875 37.065 82.795 37.295 ;
        RECT 82.815 37.105 83.245 37.890 ;
        RECT 83.275 37.065 84.625 37.975 ;
        RECT 85.335 37.295 89.235 37.975 ;
        RECT 88.305 37.065 89.235 37.295 ;
        RECT 89.245 37.295 93.145 37.975 ;
        RECT 89.245 37.065 90.175 37.295 ;
        RECT 93.395 37.065 94.745 37.975 ;
        RECT 94.765 37.165 97.515 37.975 ;
        RECT 97.985 37.295 107.175 37.975 ;
        RECT 102.495 37.075 103.425 37.295 ;
        RECT 106.255 37.065 107.175 37.295 ;
        RECT 107.185 37.165 108.555 37.975 ;
        RECT 108.575 37.105 109.005 37.890 ;
        RECT 109.025 37.165 114.535 37.975 ;
        RECT 114.545 37.165 117.295 37.975 ;
        RECT 117.305 37.165 118.675 37.975 ;
      LAYER nwell ;
        RECT 5.330 33.945 118.870 36.775 ;
      LAYER pwell ;
        RECT 5.525 32.745 6.895 33.555 ;
        RECT 6.905 32.745 12.415 33.555 ;
        RECT 12.425 32.745 17.935 33.555 ;
        RECT 18.415 32.830 18.845 33.615 ;
        RECT 18.865 32.745 20.235 33.525 ;
        RECT 20.245 32.745 22.075 33.555 ;
        RECT 25.200 33.425 26.120 33.655 ;
        RECT 30.735 33.425 31.665 33.645 ;
        RECT 34.495 33.425 35.415 33.655 ;
        RECT 22.655 32.745 26.120 33.425 ;
        RECT 26.225 32.745 35.415 33.425 ;
        RECT 35.425 32.745 40.935 33.555 ;
        RECT 40.945 32.745 42.775 33.555 ;
        RECT 42.785 32.745 44.155 33.525 ;
        RECT 44.175 32.830 44.605 33.615 ;
        RECT 45.095 32.745 46.445 33.655 ;
        RECT 46.465 32.745 51.975 33.555 ;
        RECT 51.985 32.745 57.495 33.555 ;
        RECT 57.505 32.745 63.015 33.555 ;
        RECT 63.025 32.745 65.775 33.555 ;
        RECT 65.880 33.425 66.800 33.655 ;
        RECT 65.880 32.745 69.345 33.425 ;
        RECT 69.935 32.830 70.365 33.615 ;
        RECT 70.385 32.745 71.755 33.555 ;
        RECT 71.765 32.745 73.135 33.525 ;
        RECT 73.145 33.425 74.075 33.655 ;
        RECT 90.995 33.425 91.925 33.645 ;
        RECT 94.755 33.425 95.675 33.655 ;
        RECT 73.145 32.745 77.045 33.425 ;
        RECT 77.285 32.745 86.390 33.425 ;
        RECT 86.485 32.745 95.675 33.425 ;
        RECT 95.695 32.830 96.125 33.615 ;
        RECT 96.155 32.745 97.505 33.655 ;
        RECT 97.525 32.745 101.195 33.555 ;
        RECT 101.205 32.745 102.575 33.555 ;
        RECT 102.595 32.745 103.945 33.655 ;
        RECT 103.965 32.745 109.475 33.555 ;
        RECT 109.485 32.745 114.995 33.555 ;
        RECT 115.005 32.745 116.835 33.555 ;
        RECT 117.305 32.745 118.675 33.555 ;
        RECT 5.665 32.535 5.835 32.745 ;
        RECT 7.045 32.535 7.215 32.745 ;
        RECT 12.565 32.535 12.735 32.745 ;
        RECT 13.945 32.535 14.115 32.725 ;
        RECT 15.325 32.535 15.495 32.725 ;
        RECT 18.080 32.585 18.200 32.695 ;
        RECT 19.925 32.555 20.095 32.745 ;
        RECT 20.385 32.555 20.555 32.745 ;
        RECT 22.220 32.585 22.340 32.695 ;
        RECT 22.685 32.555 22.855 32.745 ;
        RECT 24.800 32.535 24.970 32.725 ;
        RECT 26.365 32.555 26.535 32.745 ;
        RECT 28.665 32.535 28.835 32.725 ;
        RECT 30.965 32.535 31.135 32.725 ;
        RECT 32.160 32.535 32.330 32.725 ;
        RECT 35.565 32.555 35.735 32.745 ;
        RECT 36.025 32.555 36.195 32.725 ;
        RECT 40.165 32.535 40.335 32.725 ;
        RECT 40.625 32.535 40.795 32.725 ;
        RECT 41.085 32.555 41.255 32.745 ;
        RECT 43.845 32.555 44.015 32.745 ;
        RECT 44.760 32.585 44.880 32.695 ;
        RECT 45.225 32.555 45.395 32.745 ;
        RECT 46.605 32.555 46.775 32.745 ;
        RECT 50.285 32.535 50.455 32.725 ;
        RECT 52.125 32.555 52.295 32.745 ;
        RECT 53.975 32.580 54.135 32.690 ;
        RECT 56.720 32.535 56.890 32.725 ;
        RECT 57.645 32.535 57.815 32.745 ;
        RECT 59.025 32.535 59.195 32.725 ;
        RECT 62.245 32.535 62.415 32.725 ;
        RECT 63.165 32.555 63.335 32.745 ;
        RECT 69.145 32.555 69.315 32.745 ;
        RECT 69.600 32.585 69.720 32.695 ;
        RECT 70.525 32.555 70.695 32.745 ;
        RECT 71.905 32.535 72.075 32.745 ;
        RECT 73.560 32.555 73.730 32.745 ;
        RECT 77.425 32.555 77.595 32.745 ;
        RECT 81.105 32.535 81.275 32.725 ;
        RECT 82.480 32.585 82.600 32.695 ;
        RECT 83.680 32.535 83.850 32.725 ;
        RECT 86.625 32.555 86.795 32.745 ;
        RECT 87.545 32.535 87.715 32.725 ;
        RECT 97.205 32.535 97.375 32.745 ;
        RECT 97.665 32.555 97.835 32.745 ;
        RECT 101.345 32.555 101.515 32.745 ;
        RECT 102.725 32.535 102.895 32.745 ;
        RECT 104.105 32.555 104.275 32.745 ;
        RECT 108.240 32.585 108.360 32.695 ;
        RECT 109.165 32.535 109.335 32.725 ;
        RECT 109.625 32.555 109.795 32.745 ;
        RECT 114.685 32.535 114.855 32.725 ;
        RECT 115.145 32.555 115.315 32.745 ;
        RECT 116.980 32.585 117.100 32.695 ;
        RECT 118.365 32.535 118.535 32.745 ;
        RECT 5.525 31.725 6.895 32.535 ;
        RECT 6.905 31.725 12.415 32.535 ;
        RECT 12.425 31.725 13.795 32.535 ;
        RECT 13.805 31.755 15.175 32.535 ;
        RECT 15.185 31.855 24.375 32.535 ;
        RECT 19.695 31.635 20.625 31.855 ;
        RECT 23.455 31.625 24.375 31.855 ;
        RECT 24.385 31.855 28.285 32.535 ;
        RECT 24.385 31.625 25.315 31.855 ;
        RECT 28.525 31.725 29.895 32.535 ;
        RECT 29.905 31.755 31.275 32.535 ;
        RECT 31.295 31.665 31.725 32.450 ;
        RECT 31.745 31.855 35.645 32.535 ;
        RECT 36.290 31.855 38.715 32.535 ;
        RECT 31.745 31.625 32.675 31.855 ;
        RECT 39.105 31.755 40.475 32.535 ;
        RECT 40.485 31.855 49.765 32.535 ;
        RECT 41.845 31.635 42.765 31.855 ;
        RECT 47.430 31.735 49.765 31.855 ;
        RECT 48.845 31.625 49.765 31.735 ;
        RECT 50.145 31.725 53.815 32.535 ;
        RECT 54.745 31.625 57.035 32.535 ;
        RECT 57.055 31.665 57.485 32.450 ;
        RECT 57.505 31.725 58.875 32.535 ;
        RECT 58.985 31.625 62.095 32.535 ;
        RECT 62.105 31.855 71.715 32.535 ;
        RECT 71.765 31.855 80.955 32.535 ;
        RECT 66.615 31.635 67.545 31.855 ;
        RECT 70.375 31.625 71.715 31.855 ;
        RECT 76.275 31.635 77.205 31.855 ;
        RECT 80.035 31.625 80.955 31.855 ;
        RECT 80.965 31.755 82.335 32.535 ;
        RECT 82.815 31.665 83.245 32.450 ;
        RECT 83.265 31.855 87.165 32.535 ;
        RECT 87.405 31.855 96.685 32.535 ;
        RECT 83.265 31.625 84.195 31.855 ;
        RECT 88.765 31.635 89.685 31.855 ;
        RECT 94.350 31.735 96.685 31.855 ;
        RECT 95.765 31.625 96.685 31.735 ;
        RECT 97.065 31.725 102.575 32.535 ;
        RECT 102.585 31.725 108.095 32.535 ;
        RECT 108.575 31.665 109.005 32.450 ;
        RECT 109.025 31.725 114.535 32.535 ;
        RECT 114.545 31.725 117.295 32.535 ;
        RECT 117.305 31.725 118.675 32.535 ;
      LAYER nwell ;
        RECT 5.330 28.505 118.870 31.335 ;
      LAYER pwell ;
        RECT 5.525 27.305 6.895 28.115 ;
        RECT 6.905 27.305 12.415 28.115 ;
        RECT 12.425 27.305 16.095 28.115 ;
        RECT 17.035 27.305 18.385 28.215 ;
        RECT 18.415 27.390 18.845 28.175 ;
        RECT 18.865 27.985 19.795 28.215 ;
        RECT 18.865 27.305 22.765 27.985 ;
        RECT 23.015 27.305 24.365 28.215 ;
        RECT 24.385 27.305 28.055 28.115 ;
        RECT 28.065 27.305 29.435 28.115 ;
        RECT 29.530 27.305 38.635 27.985 ;
        RECT 38.655 27.305 40.005 28.215 ;
        RECT 40.025 27.305 42.775 28.115 ;
        RECT 42.795 27.305 44.145 28.215 ;
        RECT 44.175 27.390 44.605 28.175 ;
        RECT 44.625 27.985 45.555 28.215 ;
        RECT 44.625 27.305 48.525 27.985 ;
        RECT 48.765 27.305 54.275 28.115 ;
        RECT 54.285 27.305 57.955 28.115 ;
        RECT 57.965 28.015 58.895 28.215 ;
        RECT 60.230 28.015 61.175 28.215 ;
        RECT 57.965 27.535 61.175 28.015 ;
        RECT 58.105 27.335 61.175 27.535 ;
        RECT 5.665 27.095 5.835 27.305 ;
        RECT 7.045 27.095 7.215 27.305 ;
        RECT 12.565 27.095 12.735 27.305 ;
        RECT 13.945 27.095 14.115 27.285 ;
        RECT 16.255 27.150 16.415 27.260 ;
        RECT 17.165 27.115 17.335 27.305 ;
        RECT 19.280 27.115 19.450 27.305 ;
        RECT 23.145 27.095 23.315 27.285 ;
        RECT 24.065 27.115 24.235 27.305 ;
        RECT 24.525 27.115 24.695 27.305 ;
        RECT 28.205 27.115 28.375 27.305 ;
        RECT 28.665 27.095 28.835 27.285 ;
        RECT 35.105 27.095 35.275 27.285 ;
        RECT 35.565 27.095 35.735 27.285 ;
        RECT 38.325 27.095 38.495 27.305 ;
        RECT 39.705 27.115 39.875 27.305 ;
        RECT 40.165 27.115 40.335 27.305 ;
        RECT 42.925 27.115 43.095 27.305 ;
        RECT 45.040 27.115 45.210 27.305 ;
        RECT 47.985 27.095 48.155 27.285 ;
        RECT 48.905 27.115 49.075 27.305 ;
        RECT 53.505 27.095 53.675 27.285 ;
        RECT 54.425 27.115 54.595 27.305 ;
        RECT 57.645 27.095 57.815 27.285 ;
        RECT 58.105 27.115 58.275 27.335 ;
        RECT 60.230 27.305 61.175 27.335 ;
        RECT 61.185 28.015 62.130 28.215 ;
        RECT 63.465 28.015 64.395 28.215 ;
        RECT 61.185 27.535 64.395 28.015 ;
        RECT 61.185 27.335 64.255 27.535 ;
        RECT 61.185 27.305 62.130 27.335 ;
        RECT 61.780 27.095 61.950 27.285 ;
        RECT 62.245 27.095 62.415 27.285 ;
        RECT 64.085 27.115 64.255 27.335 ;
        RECT 64.405 27.305 66.235 28.115 ;
        RECT 66.715 27.305 68.065 28.215 ;
        RECT 68.085 27.305 69.915 28.115 ;
        RECT 69.935 27.390 70.365 28.175 ;
        RECT 70.385 27.305 74.055 28.115 ;
        RECT 74.985 27.985 75.905 28.215 ;
        RECT 78.735 27.985 79.665 28.205 ;
        RECT 74.985 27.305 84.175 27.985 ;
        RECT 84.195 27.305 85.545 28.215 ;
        RECT 85.565 27.305 91.075 28.115 ;
        RECT 91.085 27.305 94.755 28.115 ;
        RECT 95.695 27.390 96.125 28.175 ;
        RECT 96.145 27.305 101.655 28.115 ;
        RECT 101.665 27.305 107.175 28.115 ;
        RECT 107.185 27.305 112.695 28.115 ;
        RECT 112.705 27.305 116.375 28.115 ;
        RECT 117.305 27.305 118.675 28.115 ;
        RECT 64.545 27.095 64.715 27.305 ;
        RECT 66.380 27.145 66.500 27.255 ;
        RECT 66.845 27.115 67.015 27.305 ;
        RECT 68.225 27.115 68.395 27.305 ;
        RECT 70.065 27.095 70.235 27.285 ;
        RECT 70.525 27.115 70.695 27.305 ;
        RECT 74.215 27.150 74.375 27.260 ;
        RECT 78.805 27.095 78.975 27.285 ;
        RECT 79.265 27.095 79.435 27.285 ;
        RECT 80.645 27.095 80.815 27.285 ;
        RECT 82.480 27.145 82.600 27.255 ;
        RECT 83.405 27.095 83.575 27.285 ;
        RECT 83.865 27.115 84.035 27.305 ;
        RECT 84.325 27.115 84.495 27.305 ;
        RECT 85.705 27.115 85.875 27.305 ;
        RECT 88.925 27.095 89.095 27.285 ;
        RECT 91.225 27.115 91.395 27.305 ;
        RECT 94.445 27.095 94.615 27.285 ;
        RECT 94.915 27.150 95.075 27.260 ;
        RECT 96.285 27.115 96.455 27.305 ;
        RECT 99.965 27.095 100.135 27.285 ;
        RECT 101.805 27.115 101.975 27.305 ;
        RECT 105.485 27.095 105.655 27.285 ;
        RECT 107.325 27.115 107.495 27.305 ;
        RECT 108.240 27.145 108.360 27.255 ;
        RECT 109.165 27.095 109.335 27.285 ;
        RECT 112.845 27.115 113.015 27.305 ;
        RECT 114.685 27.095 114.855 27.285 ;
        RECT 116.535 27.150 116.695 27.260 ;
        RECT 118.365 27.095 118.535 27.305 ;
        RECT 5.525 26.285 6.895 27.095 ;
        RECT 6.905 26.285 12.415 27.095 ;
        RECT 12.425 26.285 13.795 27.095 ;
        RECT 13.805 26.415 22.995 27.095 ;
        RECT 18.315 26.195 19.245 26.415 ;
        RECT 22.075 26.185 22.995 26.415 ;
        RECT 23.005 26.285 28.515 27.095 ;
        RECT 28.525 26.285 31.275 27.095 ;
        RECT 31.295 26.225 31.725 27.010 ;
        RECT 31.840 26.415 35.305 27.095 ;
        RECT 31.840 26.185 32.760 26.415 ;
        RECT 35.425 26.285 38.175 27.095 ;
        RECT 38.185 26.415 47.465 27.095 ;
        RECT 39.545 26.195 40.465 26.415 ;
        RECT 45.130 26.295 47.465 26.415 ;
        RECT 46.545 26.185 47.465 26.295 ;
        RECT 47.845 26.285 53.355 27.095 ;
        RECT 53.365 26.285 57.035 27.095 ;
        RECT 57.055 26.225 57.485 27.010 ;
        RECT 57.505 26.285 58.875 27.095 ;
        RECT 59.175 26.185 62.095 27.095 ;
        RECT 62.105 26.415 64.395 27.095 ;
        RECT 63.475 26.185 64.395 26.415 ;
        RECT 64.405 26.285 69.915 27.095 ;
        RECT 69.925 26.285 75.435 27.095 ;
        RECT 75.540 26.415 79.005 27.095 ;
        RECT 75.540 26.185 76.460 26.415 ;
        RECT 79.135 26.185 80.485 27.095 ;
        RECT 80.505 26.285 82.335 27.095 ;
        RECT 82.815 26.225 83.245 27.010 ;
        RECT 83.265 26.285 88.775 27.095 ;
        RECT 88.785 26.285 94.295 27.095 ;
        RECT 94.305 26.285 99.815 27.095 ;
        RECT 99.825 26.285 105.335 27.095 ;
        RECT 105.345 26.285 108.095 27.095 ;
        RECT 108.575 26.225 109.005 27.010 ;
        RECT 109.025 26.285 114.535 27.095 ;
        RECT 114.545 26.285 117.295 27.095 ;
        RECT 117.305 26.285 118.675 27.095 ;
      LAYER nwell ;
        RECT 5.330 23.065 118.870 25.895 ;
      LAYER pwell ;
        RECT 5.525 21.865 6.895 22.675 ;
        RECT 6.905 21.865 12.415 22.675 ;
        RECT 12.425 21.865 17.935 22.675 ;
        RECT 18.415 21.950 18.845 22.735 ;
        RECT 18.865 21.865 24.375 22.675 ;
        RECT 24.385 21.865 27.135 22.675 ;
        RECT 31.655 22.545 32.585 22.765 ;
        RECT 35.415 22.545 36.335 22.775 ;
        RECT 27.145 21.865 36.335 22.545 ;
        RECT 36.345 21.865 41.855 22.675 ;
        RECT 41.865 21.865 43.695 22.675 ;
        RECT 44.175 21.950 44.605 22.735 ;
        RECT 44.625 21.865 46.455 22.675 ;
        RECT 46.475 21.865 47.825 22.775 ;
        RECT 47.855 21.865 49.205 22.775 ;
        RECT 49.225 21.865 50.595 22.645 ;
        RECT 50.625 21.865 51.975 22.775 ;
        RECT 53.035 22.545 53.965 22.775 ;
        RECT 56.940 22.545 57.860 22.775 ;
        RECT 59.545 22.545 62.545 22.775 ;
        RECT 52.130 21.865 53.965 22.545 ;
        RECT 54.395 21.865 57.860 22.545 ;
        RECT 57.965 22.455 62.545 22.545 ;
        RECT 57.965 22.095 62.555 22.455 ;
        RECT 57.965 21.865 59.535 22.095 ;
        RECT 61.625 21.905 62.555 22.095 ;
        RECT 61.625 21.865 62.545 21.905 ;
        RECT 62.565 21.865 64.395 22.545 ;
        RECT 64.405 21.865 65.775 22.645 ;
        RECT 65.785 21.865 69.455 22.675 ;
        RECT 69.935 21.950 70.365 22.735 ;
        RECT 70.385 21.865 75.895 22.675 ;
        RECT 75.905 21.865 81.415 22.675 ;
        RECT 81.425 21.865 86.935 22.675 ;
        RECT 86.945 21.865 92.455 22.675 ;
        RECT 92.465 21.865 95.215 22.675 ;
        RECT 95.695 21.950 96.125 22.735 ;
        RECT 96.145 21.865 101.655 22.675 ;
        RECT 101.665 21.865 107.175 22.675 ;
        RECT 107.185 21.865 112.695 22.675 ;
        RECT 112.705 21.865 116.375 22.675 ;
        RECT 117.305 21.865 118.675 22.675 ;
        RECT 5.665 21.655 5.835 21.865 ;
        RECT 7.045 21.655 7.215 21.865 ;
        RECT 12.565 21.655 12.735 21.865 ;
        RECT 18.085 21.815 18.255 21.845 ;
        RECT 18.080 21.705 18.255 21.815 ;
        RECT 18.085 21.655 18.255 21.705 ;
        RECT 19.005 21.675 19.175 21.865 ;
        RECT 23.605 21.655 23.775 21.845 ;
        RECT 24.525 21.675 24.695 21.865 ;
        RECT 27.285 21.675 27.455 21.865 ;
        RECT 29.125 21.655 29.295 21.845 ;
        RECT 30.960 21.705 31.080 21.815 ;
        RECT 31.885 21.655 32.055 21.845 ;
        RECT 36.485 21.675 36.655 21.865 ;
        RECT 37.405 21.655 37.575 21.845 ;
        RECT 42.005 21.675 42.175 21.865 ;
        RECT 42.925 21.655 43.095 21.845 ;
        RECT 43.840 21.705 43.960 21.815 ;
        RECT 44.765 21.655 44.935 21.865 ;
        RECT 46.605 21.675 46.775 21.865 ;
        RECT 48.905 21.675 49.075 21.865 ;
        RECT 50.285 21.675 50.455 21.865 ;
        RECT 50.740 21.675 50.910 21.865 ;
        RECT 52.130 21.845 52.295 21.865 ;
        RECT 52.125 21.675 52.295 21.845 ;
        RECT 53.960 21.705 54.080 21.815 ;
        RECT 54.425 21.655 54.595 21.865 ;
        RECT 56.720 21.705 56.840 21.815 ;
        RECT 57.645 21.655 57.815 21.845 ;
        RECT 58.105 21.675 58.275 21.865 ;
        RECT 59.485 21.655 59.655 21.845 ;
        RECT 62.705 21.675 62.875 21.865 ;
        RECT 64.545 21.675 64.715 21.865 ;
        RECT 65.925 21.675 66.095 21.865 ;
        RECT 69.600 21.705 69.720 21.815 ;
        RECT 70.525 21.675 70.695 21.865 ;
        RECT 73.285 21.655 73.455 21.845 ;
        RECT 73.745 21.655 73.915 21.845 ;
        RECT 76.045 21.675 76.215 21.865 ;
        RECT 79.265 21.655 79.435 21.845 ;
        RECT 81.565 21.675 81.735 21.865 ;
        RECT 83.405 21.655 83.575 21.845 ;
        RECT 87.085 21.675 87.255 21.865 ;
        RECT 88.925 21.655 89.095 21.845 ;
        RECT 92.605 21.675 92.775 21.865 ;
        RECT 94.445 21.655 94.615 21.845 ;
        RECT 95.360 21.705 95.480 21.815 ;
        RECT 96.285 21.675 96.455 21.865 ;
        RECT 99.965 21.655 100.135 21.845 ;
        RECT 101.805 21.675 101.975 21.865 ;
        RECT 105.485 21.655 105.655 21.845 ;
        RECT 107.325 21.675 107.495 21.865 ;
        RECT 108.240 21.705 108.360 21.815 ;
        RECT 109.165 21.655 109.335 21.845 ;
        RECT 112.845 21.675 113.015 21.865 ;
        RECT 114.685 21.655 114.855 21.845 ;
        RECT 116.535 21.710 116.695 21.820 ;
        RECT 118.365 21.655 118.535 21.865 ;
        RECT 5.525 20.845 6.895 21.655 ;
        RECT 6.905 20.845 12.415 21.655 ;
        RECT 12.425 20.845 17.935 21.655 ;
        RECT 17.945 20.845 23.455 21.655 ;
        RECT 23.465 20.845 28.975 21.655 ;
        RECT 28.985 20.845 30.815 21.655 ;
        RECT 31.295 20.785 31.725 21.570 ;
        RECT 31.745 20.845 37.255 21.655 ;
        RECT 37.265 20.845 42.775 21.655 ;
        RECT 42.785 20.845 44.615 21.655 ;
        RECT 44.625 20.975 53.815 21.655 ;
        RECT 54.285 20.975 56.575 21.655 ;
        RECT 49.135 20.755 50.065 20.975 ;
        RECT 52.895 20.745 53.815 20.975 ;
        RECT 55.655 20.745 56.575 20.975 ;
        RECT 57.055 20.785 57.485 21.570 ;
        RECT 57.505 20.975 59.335 21.655 ;
        RECT 59.345 20.975 63.015 21.655 ;
        RECT 62.085 20.745 63.015 20.975 ;
        RECT 63.225 20.975 73.595 21.655 ;
        RECT 63.225 20.745 65.435 20.975 ;
        RECT 68.155 20.755 69.085 20.975 ;
        RECT 73.605 20.845 79.115 21.655 ;
        RECT 79.125 20.845 82.795 21.655 ;
        RECT 82.815 20.785 83.245 21.570 ;
        RECT 83.265 20.845 88.775 21.655 ;
        RECT 88.785 20.845 94.295 21.655 ;
        RECT 94.305 20.845 99.815 21.655 ;
        RECT 99.825 20.845 105.335 21.655 ;
        RECT 105.345 20.845 108.095 21.655 ;
        RECT 108.575 20.785 109.005 21.570 ;
        RECT 109.025 20.845 114.535 21.655 ;
        RECT 114.545 20.845 117.295 21.655 ;
        RECT 117.305 20.845 118.675 21.655 ;
      LAYER nwell ;
        RECT 5.330 17.625 118.870 20.455 ;
      LAYER pwell ;
        RECT 5.525 16.425 6.895 17.235 ;
        RECT 6.905 16.425 12.415 17.235 ;
        RECT 12.425 16.425 17.935 17.235 ;
        RECT 18.415 16.510 18.845 17.295 ;
        RECT 18.865 16.425 24.375 17.235 ;
        RECT 24.385 16.425 29.895 17.235 ;
        RECT 29.905 16.425 35.415 17.235 ;
        RECT 35.425 16.425 40.935 17.235 ;
        RECT 40.945 16.425 43.695 17.235 ;
        RECT 44.175 16.510 44.605 17.295 ;
        RECT 44.625 16.425 46.455 17.235 ;
        RECT 50.975 17.105 51.905 17.325 ;
        RECT 54.735 17.105 55.655 17.335 ;
        RECT 60.175 17.105 61.105 17.325 ;
        RECT 63.935 17.105 64.855 17.335 ;
        RECT 46.465 16.425 55.655 17.105 ;
        RECT 55.665 16.425 64.855 17.105 ;
        RECT 64.875 16.425 66.225 17.335 ;
        RECT 67.175 16.425 68.525 17.335 ;
        RECT 68.545 16.425 69.915 17.235 ;
        RECT 69.935 16.510 70.365 17.295 ;
        RECT 70.385 16.425 75.895 17.235 ;
        RECT 75.905 16.425 81.415 17.235 ;
        RECT 81.425 16.425 86.935 17.235 ;
        RECT 86.945 16.425 92.455 17.235 ;
        RECT 92.465 16.425 95.215 17.235 ;
        RECT 95.695 16.510 96.125 17.295 ;
        RECT 96.145 16.425 101.655 17.235 ;
        RECT 101.665 16.425 107.175 17.235 ;
        RECT 107.185 16.425 112.695 17.235 ;
        RECT 112.705 16.425 116.375 17.235 ;
        RECT 117.305 16.425 118.675 17.235 ;
        RECT 5.665 16.215 5.835 16.425 ;
        RECT 7.045 16.215 7.215 16.425 ;
        RECT 12.565 16.215 12.735 16.425 ;
        RECT 18.085 16.375 18.255 16.405 ;
        RECT 18.080 16.265 18.255 16.375 ;
        RECT 18.085 16.215 18.255 16.265 ;
        RECT 19.005 16.235 19.175 16.425 ;
        RECT 23.605 16.215 23.775 16.405 ;
        RECT 24.525 16.235 24.695 16.425 ;
        RECT 29.125 16.215 29.295 16.405 ;
        RECT 30.045 16.235 30.215 16.425 ;
        RECT 30.960 16.265 31.080 16.375 ;
        RECT 31.885 16.215 32.055 16.405 ;
        RECT 35.565 16.235 35.735 16.425 ;
        RECT 37.405 16.215 37.575 16.405 ;
        RECT 41.085 16.235 41.255 16.425 ;
        RECT 42.925 16.215 43.095 16.405 ;
        RECT 43.840 16.265 43.960 16.375 ;
        RECT 44.765 16.235 44.935 16.425 ;
        RECT 46.605 16.235 46.775 16.425 ;
        RECT 48.445 16.215 48.615 16.405 ;
        RECT 52.135 16.260 52.295 16.370 ;
        RECT 53.045 16.215 53.215 16.405 ;
        RECT 55.805 16.235 55.975 16.425 ;
        RECT 56.275 16.260 56.435 16.370 ;
        RECT 59.025 16.215 59.195 16.405 ;
        RECT 60.405 16.215 60.575 16.405 ;
        RECT 60.865 16.215 61.035 16.405 ;
        RECT 65.925 16.235 66.095 16.425 ;
        RECT 66.385 16.215 66.555 16.405 ;
        RECT 67.305 16.235 67.475 16.425 ;
        RECT 68.685 16.235 68.855 16.425 ;
        RECT 70.525 16.235 70.695 16.425 ;
        RECT 71.905 16.215 72.075 16.405 ;
        RECT 76.045 16.235 76.215 16.425 ;
        RECT 77.425 16.215 77.595 16.405 ;
        RECT 81.565 16.235 81.735 16.425 ;
        RECT 83.405 16.215 83.575 16.405 ;
        RECT 87.085 16.235 87.255 16.425 ;
        RECT 88.925 16.215 89.095 16.405 ;
        RECT 92.605 16.235 92.775 16.425 ;
        RECT 94.445 16.215 94.615 16.405 ;
        RECT 95.360 16.265 95.480 16.375 ;
        RECT 96.285 16.235 96.455 16.425 ;
        RECT 99.965 16.215 100.135 16.405 ;
        RECT 101.805 16.235 101.975 16.425 ;
        RECT 105.485 16.215 105.655 16.405 ;
        RECT 107.325 16.235 107.495 16.425 ;
        RECT 108.240 16.265 108.360 16.375 ;
        RECT 109.165 16.215 109.335 16.405 ;
        RECT 112.845 16.235 113.015 16.425 ;
        RECT 114.685 16.215 114.855 16.405 ;
        RECT 116.535 16.270 116.695 16.380 ;
        RECT 118.365 16.215 118.535 16.425 ;
        RECT 5.525 15.405 6.895 16.215 ;
        RECT 6.905 15.405 12.415 16.215 ;
        RECT 12.425 15.405 17.935 16.215 ;
        RECT 17.945 15.405 23.455 16.215 ;
        RECT 23.465 15.405 28.975 16.215 ;
        RECT 28.985 15.405 30.815 16.215 ;
        RECT 31.295 15.345 31.725 16.130 ;
        RECT 31.745 15.405 37.255 16.215 ;
        RECT 37.265 15.405 42.775 16.215 ;
        RECT 42.785 15.405 48.295 16.215 ;
        RECT 48.305 15.405 51.975 16.215 ;
        RECT 53.005 15.305 56.115 16.215 ;
        RECT 57.055 15.345 57.485 16.130 ;
        RECT 57.505 15.535 59.335 16.215 ;
        RECT 57.505 15.305 58.850 15.535 ;
        RECT 59.355 15.305 60.705 16.215 ;
        RECT 60.725 15.405 66.235 16.215 ;
        RECT 66.245 15.405 71.755 16.215 ;
        RECT 71.765 15.405 77.275 16.215 ;
        RECT 77.285 15.405 82.795 16.215 ;
        RECT 82.815 15.345 83.245 16.130 ;
        RECT 83.265 15.405 88.775 16.215 ;
        RECT 88.785 15.405 94.295 16.215 ;
        RECT 94.305 15.405 99.815 16.215 ;
        RECT 99.825 15.405 105.335 16.215 ;
        RECT 105.345 15.405 108.095 16.215 ;
        RECT 108.575 15.345 109.005 16.130 ;
        RECT 109.025 15.405 114.535 16.215 ;
        RECT 114.545 15.405 117.295 16.215 ;
        RECT 117.305 15.405 118.675 16.215 ;
      LAYER nwell ;
        RECT 5.330 12.185 118.870 15.015 ;
      LAYER pwell ;
        RECT 5.525 10.985 6.895 11.795 ;
        RECT 6.905 10.985 12.415 11.795 ;
        RECT 12.425 10.985 17.935 11.795 ;
        RECT 18.415 11.070 18.845 11.855 ;
        RECT 18.865 10.985 24.375 11.795 ;
        RECT 24.385 10.985 29.895 11.795 ;
        RECT 29.905 10.985 31.275 11.795 ;
        RECT 31.295 11.070 31.725 11.855 ;
        RECT 31.745 10.985 37.255 11.795 ;
        RECT 37.265 10.985 42.775 11.795 ;
        RECT 42.785 10.985 44.155 11.795 ;
        RECT 44.175 11.070 44.605 11.855 ;
        RECT 44.625 10.985 50.135 11.795 ;
        RECT 50.145 10.985 55.655 11.795 ;
        RECT 55.665 10.985 57.035 11.795 ;
        RECT 57.055 11.070 57.485 11.855 ;
        RECT 57.505 10.985 63.015 11.795 ;
        RECT 63.025 10.985 68.535 11.795 ;
        RECT 68.545 10.985 69.915 11.795 ;
        RECT 69.935 11.070 70.365 11.855 ;
        RECT 70.385 10.985 75.895 11.795 ;
        RECT 75.905 10.985 81.415 11.795 ;
        RECT 81.425 10.985 82.795 11.795 ;
        RECT 82.815 11.070 83.245 11.855 ;
        RECT 83.265 10.985 88.775 11.795 ;
        RECT 88.785 10.985 94.295 11.795 ;
        RECT 94.305 10.985 95.675 11.795 ;
        RECT 95.695 11.070 96.125 11.855 ;
        RECT 96.145 10.985 101.655 11.795 ;
        RECT 101.665 10.985 107.175 11.795 ;
        RECT 107.185 10.985 108.555 11.795 ;
        RECT 108.575 11.070 109.005 11.855 ;
        RECT 109.025 10.985 114.535 11.795 ;
        RECT 114.545 10.985 117.295 11.795 ;
        RECT 117.305 10.985 118.675 11.795 ;
        RECT 5.665 10.795 5.835 10.985 ;
        RECT 7.045 10.795 7.215 10.985 ;
        RECT 12.565 10.795 12.735 10.985 ;
        RECT 18.080 10.825 18.200 10.935 ;
        RECT 19.005 10.795 19.175 10.985 ;
        RECT 24.525 10.795 24.695 10.985 ;
        RECT 30.045 10.795 30.215 10.985 ;
        RECT 31.885 10.795 32.055 10.985 ;
        RECT 37.405 10.795 37.575 10.985 ;
        RECT 42.925 10.795 43.095 10.985 ;
        RECT 44.765 10.795 44.935 10.985 ;
        RECT 50.285 10.795 50.455 10.985 ;
        RECT 55.805 10.795 55.975 10.985 ;
        RECT 57.645 10.795 57.815 10.985 ;
        RECT 63.165 10.795 63.335 10.985 ;
        RECT 68.685 10.795 68.855 10.985 ;
        RECT 70.525 10.795 70.695 10.985 ;
        RECT 76.045 10.795 76.215 10.985 ;
        RECT 81.565 10.795 81.735 10.985 ;
        RECT 83.405 10.795 83.575 10.985 ;
        RECT 88.925 10.795 89.095 10.985 ;
        RECT 94.445 10.795 94.615 10.985 ;
        RECT 96.285 10.795 96.455 10.985 ;
        RECT 101.805 10.795 101.975 10.985 ;
        RECT 107.325 10.795 107.495 10.985 ;
        RECT 109.165 10.795 109.335 10.985 ;
        RECT 114.685 10.795 114.855 10.985 ;
        RECT 118.365 10.795 118.535 10.985 ;
      LAYER li1 ;
        RECT 5.520 122.315 118.680 122.485 ;
        RECT 5.605 121.225 6.815 122.315 ;
        RECT 6.985 121.880 12.330 122.315 ;
        RECT 5.605 120.515 6.125 121.055 ;
        RECT 6.295 120.685 6.815 121.225 ;
        RECT 5.605 119.765 6.815 120.515 ;
        RECT 8.570 120.310 8.910 121.140 ;
        RECT 10.390 120.630 10.740 121.880 ;
        RECT 12.565 121.175 12.775 122.315 ;
        RECT 12.945 121.165 13.275 122.145 ;
        RECT 13.445 121.175 13.675 122.315 ;
        RECT 13.885 121.225 17.395 122.315 ;
        RECT 6.985 119.765 12.330 120.310 ;
        RECT 12.565 119.765 12.775 120.585 ;
        RECT 12.945 120.565 13.195 121.165 ;
        RECT 13.365 120.755 13.695 121.005 ;
        RECT 12.945 119.935 13.275 120.565 ;
        RECT 13.445 119.765 13.675 120.585 ;
        RECT 13.885 120.535 15.535 121.055 ;
        RECT 15.705 120.705 17.395 121.225 ;
        RECT 18.485 121.150 18.775 122.315 ;
        RECT 18.945 121.880 24.290 122.315 ;
        RECT 24.465 121.880 29.810 122.315 ;
        RECT 13.885 119.765 17.395 120.535 ;
        RECT 18.485 119.765 18.775 120.490 ;
        RECT 20.530 120.310 20.870 121.140 ;
        RECT 22.350 120.630 22.700 121.880 ;
        RECT 26.050 120.310 26.390 121.140 ;
        RECT 27.870 120.630 28.220 121.880 ;
        RECT 29.985 121.225 31.195 122.315 ;
        RECT 29.985 120.515 30.505 121.055 ;
        RECT 30.675 120.685 31.195 121.225 ;
        RECT 31.365 121.150 31.655 122.315 ;
        RECT 31.830 121.645 32.085 122.145 ;
        RECT 32.255 121.815 32.585 122.315 ;
        RECT 31.830 121.475 32.580 121.645 ;
        RECT 31.830 120.655 32.180 121.305 ;
        RECT 18.945 119.765 24.290 120.310 ;
        RECT 24.465 119.765 29.810 120.310 ;
        RECT 29.985 119.765 31.195 120.515 ;
        RECT 31.365 119.765 31.655 120.490 ;
        RECT 32.350 120.485 32.580 121.475 ;
        RECT 31.830 120.315 32.580 120.485 ;
        RECT 31.830 120.025 32.085 120.315 ;
        RECT 32.255 119.765 32.585 120.145 ;
        RECT 32.755 120.025 32.925 122.145 ;
        RECT 33.095 121.345 33.420 122.130 ;
        RECT 33.590 121.855 33.840 122.315 ;
        RECT 34.010 121.815 34.260 122.145 ;
        RECT 34.475 121.815 35.155 122.145 ;
        RECT 34.010 121.685 34.180 121.815 ;
        RECT 33.785 121.515 34.180 121.685 ;
        RECT 33.155 120.295 33.615 121.345 ;
        RECT 33.785 120.155 33.955 121.515 ;
        RECT 34.350 121.255 34.815 121.645 ;
        RECT 34.125 120.445 34.475 121.065 ;
        RECT 34.645 120.665 34.815 121.255 ;
        RECT 34.985 121.035 35.155 121.815 ;
        RECT 35.325 121.715 35.495 122.055 ;
        RECT 35.730 121.885 36.060 122.315 ;
        RECT 36.230 121.715 36.400 122.055 ;
        RECT 36.695 121.855 37.065 122.315 ;
        RECT 35.325 121.545 36.400 121.715 ;
        RECT 37.235 121.685 37.405 122.145 ;
        RECT 37.640 121.805 38.510 122.145 ;
        RECT 38.680 121.855 38.930 122.315 ;
        RECT 36.845 121.515 37.405 121.685 ;
        RECT 36.845 121.375 37.015 121.515 ;
        RECT 35.515 121.205 37.015 121.375 ;
        RECT 37.710 121.345 38.170 121.635 ;
        RECT 34.985 120.865 36.675 121.035 ;
        RECT 34.645 120.445 35.000 120.665 ;
        RECT 35.170 120.155 35.340 120.865 ;
        RECT 35.545 120.445 36.335 120.695 ;
        RECT 36.505 120.685 36.675 120.865 ;
        RECT 36.845 120.515 37.015 121.205 ;
        RECT 33.285 119.765 33.615 120.125 ;
        RECT 33.785 119.985 34.280 120.155 ;
        RECT 34.485 119.985 35.340 120.155 ;
        RECT 36.215 119.765 36.545 120.225 ;
        RECT 36.755 120.125 37.015 120.515 ;
        RECT 37.205 121.335 38.170 121.345 ;
        RECT 38.340 121.425 38.510 121.805 ;
        RECT 39.100 121.765 39.270 122.055 ;
        RECT 39.450 121.935 39.780 122.315 ;
        RECT 39.100 121.595 39.900 121.765 ;
        RECT 37.205 121.175 37.880 121.335 ;
        RECT 38.340 121.255 39.560 121.425 ;
        RECT 37.205 120.385 37.415 121.175 ;
        RECT 38.340 121.165 38.510 121.255 ;
        RECT 37.585 120.385 37.935 121.005 ;
        RECT 38.105 120.995 38.510 121.165 ;
        RECT 38.105 120.215 38.275 120.995 ;
        RECT 38.445 120.545 38.665 120.825 ;
        RECT 38.845 120.715 39.385 121.085 ;
        RECT 39.730 120.975 39.900 121.595 ;
        RECT 40.075 121.255 40.245 122.315 ;
        RECT 40.455 121.305 40.745 122.145 ;
        RECT 40.915 121.475 41.085 122.315 ;
        RECT 41.295 121.305 41.545 122.145 ;
        RECT 41.755 121.475 41.925 122.315 ;
        RECT 40.455 121.135 42.180 121.305 ;
        RECT 42.405 121.225 44.075 122.315 ;
        RECT 38.445 120.375 38.975 120.545 ;
        RECT 36.755 119.955 37.105 120.125 ;
        RECT 37.325 119.935 38.275 120.215 ;
        RECT 38.445 119.765 38.635 120.205 ;
        RECT 38.805 120.145 38.975 120.375 ;
        RECT 39.145 120.315 39.385 120.715 ;
        RECT 39.555 120.965 39.900 120.975 ;
        RECT 39.555 120.755 41.585 120.965 ;
        RECT 39.555 120.500 39.880 120.755 ;
        RECT 41.770 120.585 42.180 121.135 ;
        RECT 39.555 120.145 39.875 120.500 ;
        RECT 38.805 119.975 39.875 120.145 ;
        RECT 40.075 119.765 40.245 120.575 ;
        RECT 40.415 120.415 42.180 120.585 ;
        RECT 42.405 120.535 43.155 121.055 ;
        RECT 43.325 120.705 44.075 121.225 ;
        RECT 44.245 121.150 44.535 122.315 ;
        RECT 44.705 121.880 50.050 122.315 ;
        RECT 50.225 121.880 55.570 122.315 ;
        RECT 40.415 119.935 40.745 120.415 ;
        RECT 40.915 119.765 41.085 120.235 ;
        RECT 41.255 119.935 41.585 120.415 ;
        RECT 41.755 119.765 41.925 120.235 ;
        RECT 42.405 119.765 44.075 120.535 ;
        RECT 44.245 119.765 44.535 120.490 ;
        RECT 46.290 120.310 46.630 121.140 ;
        RECT 48.110 120.630 48.460 121.880 ;
        RECT 51.810 120.310 52.150 121.140 ;
        RECT 53.630 120.630 53.980 121.880 ;
        RECT 55.745 121.225 56.955 122.315 ;
        RECT 55.745 120.515 56.265 121.055 ;
        RECT 56.435 120.685 56.955 121.225 ;
        RECT 57.125 121.150 57.415 122.315 ;
        RECT 57.585 121.880 62.930 122.315 ;
        RECT 63.105 121.880 68.450 122.315 ;
        RECT 44.705 119.765 50.050 120.310 ;
        RECT 50.225 119.765 55.570 120.310 ;
        RECT 55.745 119.765 56.955 120.515 ;
        RECT 57.125 119.765 57.415 120.490 ;
        RECT 59.170 120.310 59.510 121.140 ;
        RECT 60.990 120.630 61.340 121.880 ;
        RECT 64.690 120.310 65.030 121.140 ;
        RECT 66.510 120.630 66.860 121.880 ;
        RECT 68.625 121.225 69.835 122.315 ;
        RECT 68.625 120.515 69.145 121.055 ;
        RECT 69.315 120.685 69.835 121.225 ;
        RECT 70.005 121.150 70.295 122.315 ;
        RECT 70.465 121.880 75.810 122.315 ;
        RECT 75.985 121.880 81.330 122.315 ;
        RECT 57.585 119.765 62.930 120.310 ;
        RECT 63.105 119.765 68.450 120.310 ;
        RECT 68.625 119.765 69.835 120.515 ;
        RECT 70.005 119.765 70.295 120.490 ;
        RECT 72.050 120.310 72.390 121.140 ;
        RECT 73.870 120.630 74.220 121.880 ;
        RECT 77.570 120.310 77.910 121.140 ;
        RECT 79.390 120.630 79.740 121.880 ;
        RECT 81.505 121.225 82.715 122.315 ;
        RECT 81.505 120.515 82.025 121.055 ;
        RECT 82.195 120.685 82.715 121.225 ;
        RECT 82.885 121.150 83.175 122.315 ;
        RECT 83.345 121.880 88.690 122.315 ;
        RECT 88.865 121.880 94.210 122.315 ;
        RECT 70.465 119.765 75.810 120.310 ;
        RECT 75.985 119.765 81.330 120.310 ;
        RECT 81.505 119.765 82.715 120.515 ;
        RECT 82.885 119.765 83.175 120.490 ;
        RECT 84.930 120.310 85.270 121.140 ;
        RECT 86.750 120.630 87.100 121.880 ;
        RECT 90.450 120.310 90.790 121.140 ;
        RECT 92.270 120.630 92.620 121.880 ;
        RECT 94.385 121.225 95.595 122.315 ;
        RECT 94.385 120.515 94.905 121.055 ;
        RECT 95.075 120.685 95.595 121.225 ;
        RECT 95.765 121.150 96.055 122.315 ;
        RECT 96.225 121.225 97.895 122.315 ;
        RECT 98.070 121.645 98.325 122.145 ;
        RECT 98.495 121.815 98.825 122.315 ;
        RECT 98.070 121.475 98.820 121.645 ;
        RECT 96.225 120.535 96.975 121.055 ;
        RECT 97.145 120.705 97.895 121.225 ;
        RECT 98.070 120.655 98.420 121.305 ;
        RECT 83.345 119.765 88.690 120.310 ;
        RECT 88.865 119.765 94.210 120.310 ;
        RECT 94.385 119.765 95.595 120.515 ;
        RECT 95.765 119.765 96.055 120.490 ;
        RECT 96.225 119.765 97.895 120.535 ;
        RECT 98.590 120.485 98.820 121.475 ;
        RECT 98.070 120.315 98.820 120.485 ;
        RECT 98.070 120.025 98.325 120.315 ;
        RECT 98.495 119.765 98.825 120.145 ;
        RECT 98.995 120.025 99.165 122.145 ;
        RECT 99.335 121.345 99.660 122.130 ;
        RECT 99.830 121.855 100.080 122.315 ;
        RECT 100.250 121.815 100.500 122.145 ;
        RECT 100.715 121.815 101.395 122.145 ;
        RECT 100.250 121.685 100.420 121.815 ;
        RECT 100.025 121.515 100.420 121.685 ;
        RECT 99.395 120.295 99.855 121.345 ;
        RECT 100.025 120.155 100.195 121.515 ;
        RECT 100.590 121.255 101.055 121.645 ;
        RECT 100.365 120.445 100.715 121.065 ;
        RECT 100.885 120.665 101.055 121.255 ;
        RECT 101.225 121.035 101.395 121.815 ;
        RECT 101.565 121.715 101.735 122.055 ;
        RECT 101.970 121.885 102.300 122.315 ;
        RECT 102.470 121.715 102.640 122.055 ;
        RECT 102.935 121.855 103.305 122.315 ;
        RECT 101.565 121.545 102.640 121.715 ;
        RECT 103.475 121.685 103.645 122.145 ;
        RECT 103.880 121.805 104.750 122.145 ;
        RECT 104.920 121.855 105.170 122.315 ;
        RECT 103.085 121.515 103.645 121.685 ;
        RECT 103.085 121.375 103.255 121.515 ;
        RECT 101.755 121.205 103.255 121.375 ;
        RECT 103.950 121.345 104.410 121.635 ;
        RECT 101.225 120.865 102.915 121.035 ;
        RECT 100.885 120.445 101.240 120.665 ;
        RECT 101.410 120.155 101.580 120.865 ;
        RECT 101.785 120.445 102.575 120.695 ;
        RECT 102.745 120.685 102.915 120.865 ;
        RECT 103.085 120.515 103.255 121.205 ;
        RECT 99.525 119.765 99.855 120.125 ;
        RECT 100.025 119.985 100.520 120.155 ;
        RECT 100.725 119.985 101.580 120.155 ;
        RECT 102.455 119.765 102.785 120.225 ;
        RECT 102.995 120.125 103.255 120.515 ;
        RECT 103.445 121.335 104.410 121.345 ;
        RECT 104.580 121.425 104.750 121.805 ;
        RECT 105.340 121.765 105.510 122.055 ;
        RECT 105.690 121.935 106.020 122.315 ;
        RECT 105.340 121.595 106.140 121.765 ;
        RECT 103.445 121.175 104.120 121.335 ;
        RECT 104.580 121.255 105.800 121.425 ;
        RECT 103.445 120.385 103.655 121.175 ;
        RECT 104.580 121.165 104.750 121.255 ;
        RECT 103.825 120.385 104.175 121.005 ;
        RECT 104.345 120.995 104.750 121.165 ;
        RECT 104.345 120.215 104.515 120.995 ;
        RECT 104.685 120.545 104.905 120.825 ;
        RECT 105.085 120.715 105.625 121.085 ;
        RECT 105.970 120.975 106.140 121.595 ;
        RECT 106.315 121.255 106.485 122.315 ;
        RECT 106.695 121.305 106.985 122.145 ;
        RECT 107.155 121.475 107.325 122.315 ;
        RECT 107.535 121.305 107.785 122.145 ;
        RECT 107.995 121.475 108.165 122.315 ;
        RECT 106.695 121.135 108.420 121.305 ;
        RECT 108.645 121.150 108.935 122.315 ;
        RECT 109.105 121.880 114.450 122.315 ;
        RECT 104.685 120.375 105.215 120.545 ;
        RECT 102.995 119.955 103.345 120.125 ;
        RECT 103.565 119.935 104.515 120.215 ;
        RECT 104.685 119.765 104.875 120.205 ;
        RECT 105.045 120.145 105.215 120.375 ;
        RECT 105.385 120.315 105.625 120.715 ;
        RECT 105.795 120.965 106.140 120.975 ;
        RECT 105.795 120.755 107.825 120.965 ;
        RECT 105.795 120.500 106.120 120.755 ;
        RECT 108.010 120.585 108.420 121.135 ;
        RECT 105.795 120.145 106.115 120.500 ;
        RECT 105.045 119.975 106.115 120.145 ;
        RECT 106.315 119.765 106.485 120.575 ;
        RECT 106.655 120.415 108.420 120.585 ;
        RECT 106.655 119.935 106.985 120.415 ;
        RECT 107.155 119.765 107.325 120.235 ;
        RECT 107.495 119.935 107.825 120.415 ;
        RECT 107.995 119.765 108.165 120.235 ;
        RECT 108.645 119.765 108.935 120.490 ;
        RECT 110.690 120.310 111.030 121.140 ;
        RECT 112.510 120.630 112.860 121.880 ;
        RECT 114.625 121.225 117.215 122.315 ;
        RECT 114.625 120.535 115.835 121.055 ;
        RECT 116.005 120.705 117.215 121.225 ;
        RECT 117.385 121.225 118.595 122.315 ;
        RECT 117.385 120.685 117.905 121.225 ;
        RECT 109.105 119.765 114.450 120.310 ;
        RECT 114.625 119.765 117.215 120.535 ;
        RECT 118.075 120.515 118.595 121.055 ;
        RECT 117.385 119.765 118.595 120.515 ;
        RECT 5.520 119.595 118.680 119.765 ;
        RECT 5.605 118.845 6.815 119.595 ;
        RECT 7.075 119.045 7.245 119.425 ;
        RECT 7.425 119.215 7.755 119.595 ;
        RECT 7.075 118.875 7.740 119.045 ;
        RECT 7.935 118.920 8.195 119.425 ;
        RECT 5.605 118.305 6.125 118.845 ;
        RECT 6.295 118.135 6.815 118.675 ;
        RECT 7.005 118.325 7.345 118.695 ;
        RECT 7.570 118.620 7.740 118.875 ;
        RECT 7.570 118.290 7.845 118.620 ;
        RECT 7.570 118.145 7.740 118.290 ;
        RECT 5.605 117.045 6.815 118.135 ;
        RECT 7.065 117.975 7.740 118.145 ;
        RECT 8.015 118.120 8.195 118.920 ;
        RECT 8.365 118.825 10.035 119.595 ;
        RECT 10.515 119.125 10.685 119.595 ;
        RECT 10.855 118.945 11.185 119.425 ;
        RECT 11.355 119.125 11.525 119.595 ;
        RECT 11.695 118.945 12.025 119.425 ;
        RECT 8.365 118.305 9.115 118.825 ;
        RECT 10.260 118.775 12.025 118.945 ;
        RECT 12.195 118.785 12.365 119.595 ;
        RECT 12.565 119.215 13.635 119.385 ;
        RECT 12.565 118.860 12.885 119.215 ;
        RECT 9.285 118.135 10.035 118.655 ;
        RECT 7.065 117.215 7.245 117.975 ;
        RECT 7.425 117.045 7.755 117.805 ;
        RECT 7.925 117.215 8.195 118.120 ;
        RECT 8.365 117.045 10.035 118.135 ;
        RECT 10.260 118.225 10.670 118.775 ;
        RECT 12.560 118.605 12.885 118.860 ;
        RECT 10.855 118.395 12.885 118.605 ;
        RECT 12.540 118.385 12.885 118.395 ;
        RECT 13.055 118.645 13.295 119.045 ;
        RECT 13.465 118.985 13.635 119.215 ;
        RECT 13.805 119.155 13.995 119.595 ;
        RECT 14.165 119.145 15.115 119.425 ;
        RECT 15.335 119.235 15.685 119.405 ;
        RECT 13.465 118.815 13.995 118.985 ;
        RECT 10.260 118.055 11.985 118.225 ;
        RECT 10.515 117.045 10.685 117.885 ;
        RECT 10.895 117.215 11.145 118.055 ;
        RECT 11.355 117.045 11.525 117.885 ;
        RECT 11.695 117.215 11.985 118.055 ;
        RECT 12.195 117.045 12.365 118.105 ;
        RECT 12.540 117.765 12.710 118.385 ;
        RECT 13.055 118.275 13.595 118.645 ;
        RECT 13.775 118.535 13.995 118.815 ;
        RECT 14.165 118.365 14.335 119.145 ;
        RECT 13.930 118.195 14.335 118.365 ;
        RECT 14.505 118.355 14.855 118.975 ;
        RECT 13.930 118.105 14.100 118.195 ;
        RECT 15.025 118.185 15.235 118.975 ;
        RECT 12.880 117.935 14.100 118.105 ;
        RECT 14.560 118.025 15.235 118.185 ;
        RECT 12.540 117.595 13.340 117.765 ;
        RECT 12.660 117.045 12.990 117.425 ;
        RECT 13.170 117.305 13.340 117.595 ;
        RECT 13.930 117.555 14.100 117.935 ;
        RECT 14.270 118.015 15.235 118.025 ;
        RECT 15.425 118.845 15.685 119.235 ;
        RECT 15.895 119.135 16.225 119.595 ;
        RECT 17.100 119.205 17.955 119.375 ;
        RECT 18.160 119.205 18.655 119.375 ;
        RECT 18.825 119.235 19.155 119.595 ;
        RECT 15.425 118.155 15.595 118.845 ;
        RECT 15.765 118.495 15.935 118.675 ;
        RECT 16.105 118.665 16.895 118.915 ;
        RECT 17.100 118.495 17.270 119.205 ;
        RECT 17.440 118.695 17.795 118.915 ;
        RECT 15.765 118.325 17.455 118.495 ;
        RECT 14.270 117.725 14.730 118.015 ;
        RECT 15.425 117.985 16.925 118.155 ;
        RECT 15.425 117.845 15.595 117.985 ;
        RECT 15.035 117.675 15.595 117.845 ;
        RECT 13.510 117.045 13.760 117.505 ;
        RECT 13.930 117.215 14.800 117.555 ;
        RECT 15.035 117.215 15.205 117.675 ;
        RECT 16.040 117.645 17.115 117.815 ;
        RECT 15.375 117.045 15.745 117.505 ;
        RECT 16.040 117.305 16.210 117.645 ;
        RECT 16.380 117.045 16.710 117.475 ;
        RECT 16.945 117.305 17.115 117.645 ;
        RECT 17.285 117.545 17.455 118.325 ;
        RECT 17.625 118.105 17.795 118.695 ;
        RECT 17.965 118.295 18.315 118.915 ;
        RECT 17.625 117.715 18.090 118.105 ;
        RECT 18.485 117.845 18.655 119.205 ;
        RECT 18.825 118.015 19.285 119.065 ;
        RECT 18.260 117.675 18.655 117.845 ;
        RECT 18.260 117.545 18.430 117.675 ;
        RECT 17.285 117.215 17.965 117.545 ;
        RECT 18.180 117.215 18.430 117.545 ;
        RECT 18.600 117.045 18.850 117.505 ;
        RECT 19.020 117.230 19.345 118.015 ;
        RECT 19.515 117.215 19.685 119.335 ;
        RECT 19.855 119.215 20.185 119.595 ;
        RECT 20.355 119.045 20.610 119.335 ;
        RECT 19.860 118.875 20.610 119.045 ;
        RECT 20.790 119.045 21.045 119.335 ;
        RECT 21.215 119.215 21.545 119.595 ;
        RECT 20.790 118.875 21.540 119.045 ;
        RECT 19.860 117.885 20.090 118.875 ;
        RECT 20.260 118.055 20.610 118.705 ;
        RECT 20.790 118.055 21.140 118.705 ;
        RECT 21.310 117.885 21.540 118.875 ;
        RECT 19.860 117.715 20.610 117.885 ;
        RECT 19.855 117.045 20.185 117.545 ;
        RECT 20.355 117.215 20.610 117.715 ;
        RECT 20.790 117.715 21.540 117.885 ;
        RECT 20.790 117.215 21.045 117.715 ;
        RECT 21.215 117.045 21.545 117.545 ;
        RECT 21.715 117.215 21.885 119.335 ;
        RECT 22.245 119.235 22.575 119.595 ;
        RECT 22.745 119.205 23.240 119.375 ;
        RECT 23.445 119.205 24.300 119.375 ;
        RECT 22.115 118.015 22.575 119.065 ;
        RECT 22.055 117.230 22.380 118.015 ;
        RECT 22.745 117.845 22.915 119.205 ;
        RECT 23.085 118.295 23.435 118.915 ;
        RECT 23.605 118.695 23.960 118.915 ;
        RECT 23.605 118.105 23.775 118.695 ;
        RECT 24.130 118.495 24.300 119.205 ;
        RECT 25.175 119.135 25.505 119.595 ;
        RECT 25.715 119.235 26.065 119.405 ;
        RECT 24.505 118.665 25.295 118.915 ;
        RECT 25.715 118.845 25.975 119.235 ;
        RECT 26.285 119.145 27.235 119.425 ;
        RECT 27.405 119.155 27.595 119.595 ;
        RECT 27.765 119.215 28.835 119.385 ;
        RECT 25.465 118.495 25.635 118.675 ;
        RECT 22.745 117.675 23.140 117.845 ;
        RECT 23.310 117.715 23.775 118.105 ;
        RECT 23.945 118.325 25.635 118.495 ;
        RECT 22.970 117.545 23.140 117.675 ;
        RECT 23.945 117.545 24.115 118.325 ;
        RECT 25.805 118.155 25.975 118.845 ;
        RECT 24.475 117.985 25.975 118.155 ;
        RECT 26.165 118.185 26.375 118.975 ;
        RECT 26.545 118.355 26.895 118.975 ;
        RECT 27.065 118.365 27.235 119.145 ;
        RECT 27.765 118.985 27.935 119.215 ;
        RECT 27.405 118.815 27.935 118.985 ;
        RECT 27.405 118.535 27.625 118.815 ;
        RECT 28.105 118.645 28.345 119.045 ;
        RECT 27.065 118.195 27.470 118.365 ;
        RECT 27.805 118.275 28.345 118.645 ;
        RECT 28.515 118.860 28.835 119.215 ;
        RECT 28.515 118.605 28.840 118.860 ;
        RECT 29.035 118.785 29.205 119.595 ;
        RECT 29.375 118.945 29.705 119.425 ;
        RECT 29.875 119.125 30.045 119.595 ;
        RECT 30.215 118.945 30.545 119.425 ;
        RECT 30.715 119.125 30.885 119.595 ;
        RECT 29.375 118.775 31.140 118.945 ;
        RECT 31.365 118.870 31.655 119.595 ;
        RECT 28.515 118.395 30.545 118.605 ;
        RECT 28.515 118.385 28.860 118.395 ;
        RECT 26.165 118.025 26.840 118.185 ;
        RECT 27.300 118.105 27.470 118.195 ;
        RECT 26.165 118.015 27.130 118.025 ;
        RECT 25.805 117.845 25.975 117.985 ;
        RECT 22.550 117.045 22.800 117.505 ;
        RECT 22.970 117.215 23.220 117.545 ;
        RECT 23.435 117.215 24.115 117.545 ;
        RECT 24.285 117.645 25.360 117.815 ;
        RECT 25.805 117.675 26.365 117.845 ;
        RECT 26.670 117.725 27.130 118.015 ;
        RECT 27.300 117.935 28.520 118.105 ;
        RECT 24.285 117.305 24.455 117.645 ;
        RECT 24.690 117.045 25.020 117.475 ;
        RECT 25.190 117.305 25.360 117.645 ;
        RECT 25.655 117.045 26.025 117.505 ;
        RECT 26.195 117.215 26.365 117.675 ;
        RECT 27.300 117.555 27.470 117.935 ;
        RECT 28.690 117.765 28.860 118.385 ;
        RECT 30.730 118.225 31.140 118.775 ;
        RECT 31.825 118.825 35.335 119.595 ;
        RECT 35.970 119.045 36.225 119.335 ;
        RECT 36.395 119.215 36.725 119.595 ;
        RECT 35.970 118.875 36.720 119.045 ;
        RECT 31.825 118.305 33.475 118.825 ;
        RECT 26.600 117.215 27.470 117.555 ;
        RECT 28.060 117.595 28.860 117.765 ;
        RECT 27.640 117.045 27.890 117.505 ;
        RECT 28.060 117.305 28.230 117.595 ;
        RECT 28.410 117.045 28.740 117.425 ;
        RECT 29.035 117.045 29.205 118.105 ;
        RECT 29.415 118.055 31.140 118.225 ;
        RECT 29.415 117.215 29.705 118.055 ;
        RECT 29.875 117.045 30.045 117.885 ;
        RECT 30.255 117.215 30.505 118.055 ;
        RECT 30.715 117.045 30.885 117.885 ;
        RECT 31.365 117.045 31.655 118.210 ;
        RECT 33.645 118.135 35.335 118.655 ;
        RECT 31.825 117.045 35.335 118.135 ;
        RECT 35.970 118.055 36.320 118.705 ;
        RECT 36.490 117.885 36.720 118.875 ;
        RECT 35.970 117.715 36.720 117.885 ;
        RECT 35.970 117.215 36.225 117.715 ;
        RECT 36.395 117.045 36.725 117.545 ;
        RECT 36.895 117.215 37.065 119.335 ;
        RECT 37.425 119.235 37.755 119.595 ;
        RECT 37.925 119.205 38.420 119.375 ;
        RECT 38.625 119.205 39.480 119.375 ;
        RECT 37.295 118.015 37.755 119.065 ;
        RECT 37.235 117.230 37.560 118.015 ;
        RECT 37.925 117.845 38.095 119.205 ;
        RECT 38.265 118.295 38.615 118.915 ;
        RECT 38.785 118.695 39.140 118.915 ;
        RECT 38.785 118.105 38.955 118.695 ;
        RECT 39.310 118.495 39.480 119.205 ;
        RECT 40.355 119.135 40.685 119.595 ;
        RECT 40.895 119.235 41.245 119.405 ;
        RECT 39.685 118.665 40.475 118.915 ;
        RECT 40.895 118.845 41.155 119.235 ;
        RECT 41.465 119.145 42.415 119.425 ;
        RECT 42.585 119.155 42.775 119.595 ;
        RECT 42.945 119.215 44.015 119.385 ;
        RECT 40.645 118.495 40.815 118.675 ;
        RECT 37.925 117.675 38.320 117.845 ;
        RECT 38.490 117.715 38.955 118.105 ;
        RECT 39.125 118.325 40.815 118.495 ;
        RECT 38.150 117.545 38.320 117.675 ;
        RECT 39.125 117.545 39.295 118.325 ;
        RECT 40.985 118.155 41.155 118.845 ;
        RECT 39.655 117.985 41.155 118.155 ;
        RECT 41.345 118.185 41.555 118.975 ;
        RECT 41.725 118.355 42.075 118.975 ;
        RECT 42.245 118.365 42.415 119.145 ;
        RECT 42.945 118.985 43.115 119.215 ;
        RECT 42.585 118.815 43.115 118.985 ;
        RECT 42.585 118.535 42.805 118.815 ;
        RECT 43.285 118.645 43.525 119.045 ;
        RECT 42.245 118.195 42.650 118.365 ;
        RECT 42.985 118.275 43.525 118.645 ;
        RECT 43.695 118.860 44.015 119.215 ;
        RECT 43.695 118.605 44.020 118.860 ;
        RECT 44.215 118.785 44.385 119.595 ;
        RECT 44.555 118.945 44.885 119.425 ;
        RECT 45.055 119.125 45.225 119.595 ;
        RECT 45.395 118.945 45.725 119.425 ;
        RECT 45.895 119.125 46.065 119.595 ;
        RECT 46.550 119.045 46.805 119.335 ;
        RECT 46.975 119.215 47.305 119.595 ;
        RECT 44.555 118.775 46.320 118.945 ;
        RECT 46.550 118.875 47.300 119.045 ;
        RECT 43.695 118.395 45.725 118.605 ;
        RECT 43.695 118.385 44.040 118.395 ;
        RECT 41.345 118.025 42.020 118.185 ;
        RECT 42.480 118.105 42.650 118.195 ;
        RECT 41.345 118.015 42.310 118.025 ;
        RECT 40.985 117.845 41.155 117.985 ;
        RECT 37.730 117.045 37.980 117.505 ;
        RECT 38.150 117.215 38.400 117.545 ;
        RECT 38.615 117.215 39.295 117.545 ;
        RECT 39.465 117.645 40.540 117.815 ;
        RECT 40.985 117.675 41.545 117.845 ;
        RECT 41.850 117.725 42.310 118.015 ;
        RECT 42.480 117.935 43.700 118.105 ;
        RECT 39.465 117.305 39.635 117.645 ;
        RECT 39.870 117.045 40.200 117.475 ;
        RECT 40.370 117.305 40.540 117.645 ;
        RECT 40.835 117.045 41.205 117.505 ;
        RECT 41.375 117.215 41.545 117.675 ;
        RECT 42.480 117.555 42.650 117.935 ;
        RECT 43.870 117.765 44.040 118.385 ;
        RECT 45.910 118.225 46.320 118.775 ;
        RECT 41.780 117.215 42.650 117.555 ;
        RECT 43.240 117.595 44.040 117.765 ;
        RECT 42.820 117.045 43.070 117.505 ;
        RECT 43.240 117.305 43.410 117.595 ;
        RECT 43.590 117.045 43.920 117.425 ;
        RECT 44.215 117.045 44.385 118.105 ;
        RECT 44.595 118.055 46.320 118.225 ;
        RECT 46.550 118.055 46.900 118.705 ;
        RECT 44.595 117.215 44.885 118.055 ;
        RECT 45.055 117.045 45.225 117.885 ;
        RECT 45.435 117.215 45.685 118.055 ;
        RECT 47.070 117.885 47.300 118.875 ;
        RECT 45.895 117.045 46.065 117.885 ;
        RECT 46.550 117.715 47.300 117.885 ;
        RECT 46.550 117.215 46.805 117.715 ;
        RECT 46.975 117.045 47.305 117.545 ;
        RECT 47.475 117.215 47.645 119.335 ;
        RECT 48.005 119.235 48.335 119.595 ;
        RECT 48.505 119.205 49.000 119.375 ;
        RECT 49.205 119.205 50.060 119.375 ;
        RECT 47.875 118.015 48.335 119.065 ;
        RECT 47.815 117.230 48.140 118.015 ;
        RECT 48.505 117.845 48.675 119.205 ;
        RECT 48.845 118.295 49.195 118.915 ;
        RECT 49.365 118.695 49.720 118.915 ;
        RECT 49.365 118.105 49.535 118.695 ;
        RECT 49.890 118.495 50.060 119.205 ;
        RECT 50.935 119.135 51.265 119.595 ;
        RECT 51.475 119.235 51.825 119.405 ;
        RECT 50.265 118.665 51.055 118.915 ;
        RECT 51.475 118.845 51.735 119.235 ;
        RECT 52.045 119.145 52.995 119.425 ;
        RECT 53.165 119.155 53.355 119.595 ;
        RECT 53.525 119.215 54.595 119.385 ;
        RECT 51.225 118.495 51.395 118.675 ;
        RECT 48.505 117.675 48.900 117.845 ;
        RECT 49.070 117.715 49.535 118.105 ;
        RECT 49.705 118.325 51.395 118.495 ;
        RECT 48.730 117.545 48.900 117.675 ;
        RECT 49.705 117.545 49.875 118.325 ;
        RECT 51.565 118.155 51.735 118.845 ;
        RECT 50.235 117.985 51.735 118.155 ;
        RECT 51.925 118.185 52.135 118.975 ;
        RECT 52.305 118.355 52.655 118.975 ;
        RECT 52.825 118.365 52.995 119.145 ;
        RECT 53.525 118.985 53.695 119.215 ;
        RECT 53.165 118.815 53.695 118.985 ;
        RECT 53.165 118.535 53.385 118.815 ;
        RECT 53.865 118.645 54.105 119.045 ;
        RECT 52.825 118.195 53.230 118.365 ;
        RECT 53.565 118.275 54.105 118.645 ;
        RECT 54.275 118.860 54.595 119.215 ;
        RECT 54.275 118.605 54.600 118.860 ;
        RECT 54.795 118.785 54.965 119.595 ;
        RECT 55.135 118.945 55.465 119.425 ;
        RECT 55.635 119.125 55.805 119.595 ;
        RECT 55.975 118.945 56.305 119.425 ;
        RECT 56.475 119.125 56.645 119.595 ;
        RECT 55.135 118.775 56.900 118.945 ;
        RECT 57.125 118.870 57.415 119.595 ;
        RECT 54.275 118.395 56.305 118.605 ;
        RECT 54.275 118.385 54.620 118.395 ;
        RECT 51.925 118.025 52.600 118.185 ;
        RECT 53.060 118.105 53.230 118.195 ;
        RECT 51.925 118.015 52.890 118.025 ;
        RECT 51.565 117.845 51.735 117.985 ;
        RECT 48.310 117.045 48.560 117.505 ;
        RECT 48.730 117.215 48.980 117.545 ;
        RECT 49.195 117.215 49.875 117.545 ;
        RECT 50.045 117.645 51.120 117.815 ;
        RECT 51.565 117.675 52.125 117.845 ;
        RECT 52.430 117.725 52.890 118.015 ;
        RECT 53.060 117.935 54.280 118.105 ;
        RECT 50.045 117.305 50.215 117.645 ;
        RECT 50.450 117.045 50.780 117.475 ;
        RECT 50.950 117.305 51.120 117.645 ;
        RECT 51.415 117.045 51.785 117.505 ;
        RECT 51.955 117.215 52.125 117.675 ;
        RECT 53.060 117.555 53.230 117.935 ;
        RECT 54.450 117.765 54.620 118.385 ;
        RECT 56.490 118.225 56.900 118.775 ;
        RECT 57.585 118.825 59.255 119.595 ;
        RECT 59.430 119.045 59.685 119.335 ;
        RECT 59.855 119.215 60.185 119.595 ;
        RECT 59.430 118.875 60.180 119.045 ;
        RECT 57.585 118.305 58.335 118.825 ;
        RECT 52.360 117.215 53.230 117.555 ;
        RECT 53.820 117.595 54.620 117.765 ;
        RECT 53.400 117.045 53.650 117.505 ;
        RECT 53.820 117.305 53.990 117.595 ;
        RECT 54.170 117.045 54.500 117.425 ;
        RECT 54.795 117.045 54.965 118.105 ;
        RECT 55.175 118.055 56.900 118.225 ;
        RECT 55.175 117.215 55.465 118.055 ;
        RECT 55.635 117.045 55.805 117.885 ;
        RECT 56.015 117.215 56.265 118.055 ;
        RECT 56.475 117.045 56.645 117.885 ;
        RECT 57.125 117.045 57.415 118.210 ;
        RECT 58.505 118.135 59.255 118.655 ;
        RECT 57.585 117.045 59.255 118.135 ;
        RECT 59.430 118.055 59.780 118.705 ;
        RECT 59.950 117.885 60.180 118.875 ;
        RECT 59.430 117.715 60.180 117.885 ;
        RECT 59.430 117.215 59.685 117.715 ;
        RECT 59.855 117.045 60.185 117.545 ;
        RECT 60.355 117.215 60.525 119.335 ;
        RECT 60.885 119.235 61.215 119.595 ;
        RECT 61.385 119.205 61.880 119.375 ;
        RECT 62.085 119.205 62.940 119.375 ;
        RECT 60.755 118.015 61.215 119.065 ;
        RECT 60.695 117.230 61.020 118.015 ;
        RECT 61.385 117.845 61.555 119.205 ;
        RECT 61.725 118.295 62.075 118.915 ;
        RECT 62.245 118.695 62.600 118.915 ;
        RECT 62.245 118.105 62.415 118.695 ;
        RECT 62.770 118.495 62.940 119.205 ;
        RECT 63.815 119.135 64.145 119.595 ;
        RECT 64.355 119.235 64.705 119.405 ;
        RECT 63.145 118.665 63.935 118.915 ;
        RECT 64.355 118.845 64.615 119.235 ;
        RECT 64.925 119.145 65.875 119.425 ;
        RECT 66.045 119.155 66.235 119.595 ;
        RECT 66.405 119.215 67.475 119.385 ;
        RECT 64.105 118.495 64.275 118.675 ;
        RECT 61.385 117.675 61.780 117.845 ;
        RECT 61.950 117.715 62.415 118.105 ;
        RECT 62.585 118.325 64.275 118.495 ;
        RECT 61.610 117.545 61.780 117.675 ;
        RECT 62.585 117.545 62.755 118.325 ;
        RECT 64.445 118.155 64.615 118.845 ;
        RECT 63.115 117.985 64.615 118.155 ;
        RECT 64.805 118.185 65.015 118.975 ;
        RECT 65.185 118.355 65.535 118.975 ;
        RECT 65.705 118.365 65.875 119.145 ;
        RECT 66.405 118.985 66.575 119.215 ;
        RECT 66.045 118.815 66.575 118.985 ;
        RECT 66.045 118.535 66.265 118.815 ;
        RECT 66.745 118.645 66.985 119.045 ;
        RECT 65.705 118.195 66.110 118.365 ;
        RECT 66.445 118.275 66.985 118.645 ;
        RECT 67.155 118.860 67.475 119.215 ;
        RECT 67.155 118.605 67.480 118.860 ;
        RECT 67.675 118.785 67.845 119.595 ;
        RECT 68.015 118.945 68.345 119.425 ;
        RECT 68.515 119.125 68.685 119.595 ;
        RECT 68.855 118.945 69.185 119.425 ;
        RECT 69.355 119.125 69.525 119.595 ;
        RECT 70.010 119.045 70.265 119.335 ;
        RECT 70.435 119.215 70.765 119.595 ;
        RECT 68.015 118.775 69.780 118.945 ;
        RECT 70.010 118.875 70.760 119.045 ;
        RECT 67.155 118.395 69.185 118.605 ;
        RECT 67.155 118.385 67.500 118.395 ;
        RECT 64.805 118.025 65.480 118.185 ;
        RECT 65.940 118.105 66.110 118.195 ;
        RECT 64.805 118.015 65.770 118.025 ;
        RECT 64.445 117.845 64.615 117.985 ;
        RECT 61.190 117.045 61.440 117.505 ;
        RECT 61.610 117.215 61.860 117.545 ;
        RECT 62.075 117.215 62.755 117.545 ;
        RECT 62.925 117.645 64.000 117.815 ;
        RECT 64.445 117.675 65.005 117.845 ;
        RECT 65.310 117.725 65.770 118.015 ;
        RECT 65.940 117.935 67.160 118.105 ;
        RECT 62.925 117.305 63.095 117.645 ;
        RECT 63.330 117.045 63.660 117.475 ;
        RECT 63.830 117.305 64.000 117.645 ;
        RECT 64.295 117.045 64.665 117.505 ;
        RECT 64.835 117.215 65.005 117.675 ;
        RECT 65.940 117.555 66.110 117.935 ;
        RECT 67.330 117.765 67.500 118.385 ;
        RECT 69.370 118.225 69.780 118.775 ;
        RECT 65.240 117.215 66.110 117.555 ;
        RECT 66.700 117.595 67.500 117.765 ;
        RECT 66.280 117.045 66.530 117.505 ;
        RECT 66.700 117.305 66.870 117.595 ;
        RECT 67.050 117.045 67.380 117.425 ;
        RECT 67.675 117.045 67.845 118.105 ;
        RECT 68.055 118.055 69.780 118.225 ;
        RECT 70.010 118.055 70.360 118.705 ;
        RECT 68.055 117.215 68.345 118.055 ;
        RECT 68.515 117.045 68.685 117.885 ;
        RECT 68.895 117.215 69.145 118.055 ;
        RECT 70.530 117.885 70.760 118.875 ;
        RECT 69.355 117.045 69.525 117.885 ;
        RECT 70.010 117.715 70.760 117.885 ;
        RECT 70.010 117.215 70.265 117.715 ;
        RECT 70.435 117.045 70.765 117.545 ;
        RECT 70.935 117.215 71.105 119.335 ;
        RECT 71.465 119.235 71.795 119.595 ;
        RECT 71.965 119.205 72.460 119.375 ;
        RECT 72.665 119.205 73.520 119.375 ;
        RECT 71.335 118.015 71.795 119.065 ;
        RECT 71.275 117.230 71.600 118.015 ;
        RECT 71.965 117.845 72.135 119.205 ;
        RECT 72.305 118.295 72.655 118.915 ;
        RECT 72.825 118.695 73.180 118.915 ;
        RECT 72.825 118.105 72.995 118.695 ;
        RECT 73.350 118.495 73.520 119.205 ;
        RECT 74.395 119.135 74.725 119.595 ;
        RECT 74.935 119.235 75.285 119.405 ;
        RECT 73.725 118.665 74.515 118.915 ;
        RECT 74.935 118.845 75.195 119.235 ;
        RECT 75.505 119.145 76.455 119.425 ;
        RECT 76.625 119.155 76.815 119.595 ;
        RECT 76.985 119.215 78.055 119.385 ;
        RECT 74.685 118.495 74.855 118.675 ;
        RECT 71.965 117.675 72.360 117.845 ;
        RECT 72.530 117.715 72.995 118.105 ;
        RECT 73.165 118.325 74.855 118.495 ;
        RECT 72.190 117.545 72.360 117.675 ;
        RECT 73.165 117.545 73.335 118.325 ;
        RECT 75.025 118.155 75.195 118.845 ;
        RECT 73.695 117.985 75.195 118.155 ;
        RECT 75.385 118.185 75.595 118.975 ;
        RECT 75.765 118.355 76.115 118.975 ;
        RECT 76.285 118.365 76.455 119.145 ;
        RECT 76.985 118.985 77.155 119.215 ;
        RECT 76.625 118.815 77.155 118.985 ;
        RECT 76.625 118.535 76.845 118.815 ;
        RECT 77.325 118.645 77.565 119.045 ;
        RECT 76.285 118.195 76.690 118.365 ;
        RECT 77.025 118.275 77.565 118.645 ;
        RECT 77.735 118.860 78.055 119.215 ;
        RECT 77.735 118.605 78.060 118.860 ;
        RECT 78.255 118.785 78.425 119.595 ;
        RECT 78.595 118.945 78.925 119.425 ;
        RECT 79.095 119.125 79.265 119.595 ;
        RECT 79.435 118.945 79.765 119.425 ;
        RECT 79.935 119.125 80.105 119.595 ;
        RECT 78.595 118.775 80.360 118.945 ;
        RECT 80.625 118.775 80.855 119.595 ;
        RECT 81.025 118.795 81.355 119.425 ;
        RECT 77.735 118.395 79.765 118.605 ;
        RECT 77.735 118.385 78.080 118.395 ;
        RECT 75.385 118.025 76.060 118.185 ;
        RECT 76.520 118.105 76.690 118.195 ;
        RECT 75.385 118.015 76.350 118.025 ;
        RECT 75.025 117.845 75.195 117.985 ;
        RECT 71.770 117.045 72.020 117.505 ;
        RECT 72.190 117.215 72.440 117.545 ;
        RECT 72.655 117.215 73.335 117.545 ;
        RECT 73.505 117.645 74.580 117.815 ;
        RECT 75.025 117.675 75.585 117.845 ;
        RECT 75.890 117.725 76.350 118.015 ;
        RECT 76.520 117.935 77.740 118.105 ;
        RECT 73.505 117.305 73.675 117.645 ;
        RECT 73.910 117.045 74.240 117.475 ;
        RECT 74.410 117.305 74.580 117.645 ;
        RECT 74.875 117.045 75.245 117.505 ;
        RECT 75.415 117.215 75.585 117.675 ;
        RECT 76.520 117.555 76.690 117.935 ;
        RECT 77.910 117.765 78.080 118.385 ;
        RECT 79.950 118.225 80.360 118.775 ;
        RECT 80.605 118.355 80.935 118.605 ;
        RECT 75.820 117.215 76.690 117.555 ;
        RECT 77.280 117.595 78.080 117.765 ;
        RECT 76.860 117.045 77.110 117.505 ;
        RECT 77.280 117.305 77.450 117.595 ;
        RECT 77.630 117.045 77.960 117.425 ;
        RECT 78.255 117.045 78.425 118.105 ;
        RECT 78.635 118.055 80.360 118.225 ;
        RECT 81.105 118.195 81.355 118.795 ;
        RECT 81.525 118.775 81.735 119.595 ;
        RECT 82.885 118.870 83.175 119.595 ;
        RECT 83.350 119.045 83.605 119.335 ;
        RECT 83.775 119.215 84.105 119.595 ;
        RECT 83.350 118.875 84.100 119.045 ;
        RECT 78.635 117.215 78.925 118.055 ;
        RECT 79.095 117.045 79.265 117.885 ;
        RECT 79.475 117.215 79.725 118.055 ;
        RECT 79.935 117.045 80.105 117.885 ;
        RECT 80.625 117.045 80.855 118.185 ;
        RECT 81.025 117.215 81.355 118.195 ;
        RECT 81.525 117.045 81.735 118.185 ;
        RECT 82.885 117.045 83.175 118.210 ;
        RECT 83.350 118.055 83.700 118.705 ;
        RECT 83.870 117.885 84.100 118.875 ;
        RECT 83.350 117.715 84.100 117.885 ;
        RECT 83.350 117.215 83.605 117.715 ;
        RECT 83.775 117.045 84.105 117.545 ;
        RECT 84.275 117.215 84.445 119.335 ;
        RECT 84.805 119.235 85.135 119.595 ;
        RECT 85.305 119.205 85.800 119.375 ;
        RECT 86.005 119.205 86.860 119.375 ;
        RECT 84.675 118.015 85.135 119.065 ;
        RECT 84.615 117.230 84.940 118.015 ;
        RECT 85.305 117.845 85.475 119.205 ;
        RECT 85.645 118.295 85.995 118.915 ;
        RECT 86.165 118.695 86.520 118.915 ;
        RECT 86.165 118.105 86.335 118.695 ;
        RECT 86.690 118.495 86.860 119.205 ;
        RECT 87.735 119.135 88.065 119.595 ;
        RECT 88.275 119.235 88.625 119.405 ;
        RECT 87.065 118.665 87.855 118.915 ;
        RECT 88.275 118.845 88.535 119.235 ;
        RECT 88.845 119.145 89.795 119.425 ;
        RECT 89.965 119.155 90.155 119.595 ;
        RECT 90.325 119.215 91.395 119.385 ;
        RECT 88.025 118.495 88.195 118.675 ;
        RECT 85.305 117.675 85.700 117.845 ;
        RECT 85.870 117.715 86.335 118.105 ;
        RECT 86.505 118.325 88.195 118.495 ;
        RECT 85.530 117.545 85.700 117.675 ;
        RECT 86.505 117.545 86.675 118.325 ;
        RECT 88.365 118.155 88.535 118.845 ;
        RECT 87.035 117.985 88.535 118.155 ;
        RECT 88.725 118.185 88.935 118.975 ;
        RECT 89.105 118.355 89.455 118.975 ;
        RECT 89.625 118.365 89.795 119.145 ;
        RECT 90.325 118.985 90.495 119.215 ;
        RECT 89.965 118.815 90.495 118.985 ;
        RECT 89.965 118.535 90.185 118.815 ;
        RECT 90.665 118.645 90.905 119.045 ;
        RECT 89.625 118.195 90.030 118.365 ;
        RECT 90.365 118.275 90.905 118.645 ;
        RECT 91.075 118.860 91.395 119.215 ;
        RECT 91.075 118.605 91.400 118.860 ;
        RECT 91.595 118.785 91.765 119.595 ;
        RECT 91.935 118.945 92.265 119.425 ;
        RECT 92.435 119.125 92.605 119.595 ;
        RECT 92.775 118.945 93.105 119.425 ;
        RECT 93.275 119.125 93.445 119.595 ;
        RECT 94.235 119.125 94.405 119.595 ;
        RECT 94.575 118.945 94.905 119.425 ;
        RECT 95.075 119.125 95.245 119.595 ;
        RECT 95.415 118.945 95.745 119.425 ;
        RECT 91.935 118.775 93.700 118.945 ;
        RECT 91.075 118.395 93.105 118.605 ;
        RECT 91.075 118.385 91.420 118.395 ;
        RECT 88.725 118.025 89.400 118.185 ;
        RECT 89.860 118.105 90.030 118.195 ;
        RECT 88.725 118.015 89.690 118.025 ;
        RECT 88.365 117.845 88.535 117.985 ;
        RECT 85.110 117.045 85.360 117.505 ;
        RECT 85.530 117.215 85.780 117.545 ;
        RECT 85.995 117.215 86.675 117.545 ;
        RECT 86.845 117.645 87.920 117.815 ;
        RECT 88.365 117.675 88.925 117.845 ;
        RECT 89.230 117.725 89.690 118.015 ;
        RECT 89.860 117.935 91.080 118.105 ;
        RECT 86.845 117.305 87.015 117.645 ;
        RECT 87.250 117.045 87.580 117.475 ;
        RECT 87.750 117.305 87.920 117.645 ;
        RECT 88.215 117.045 88.585 117.505 ;
        RECT 88.755 117.215 88.925 117.675 ;
        RECT 89.860 117.555 90.030 117.935 ;
        RECT 91.250 117.765 91.420 118.385 ;
        RECT 93.290 118.225 93.700 118.775 ;
        RECT 89.160 117.215 90.030 117.555 ;
        RECT 90.620 117.595 91.420 117.765 ;
        RECT 90.200 117.045 90.450 117.505 ;
        RECT 90.620 117.305 90.790 117.595 ;
        RECT 90.970 117.045 91.300 117.425 ;
        RECT 91.595 117.045 91.765 118.105 ;
        RECT 91.975 118.055 93.700 118.225 ;
        RECT 93.980 118.775 95.745 118.945 ;
        RECT 95.915 118.785 96.085 119.595 ;
        RECT 96.285 119.215 97.355 119.385 ;
        RECT 96.285 118.860 96.605 119.215 ;
        RECT 93.980 118.225 94.390 118.775 ;
        RECT 96.280 118.605 96.605 118.860 ;
        RECT 94.575 118.395 96.605 118.605 ;
        RECT 96.260 118.385 96.605 118.395 ;
        RECT 96.775 118.645 97.015 119.045 ;
        RECT 97.185 118.985 97.355 119.215 ;
        RECT 97.525 119.155 97.715 119.595 ;
        RECT 97.885 119.145 98.835 119.425 ;
        RECT 99.055 119.235 99.405 119.405 ;
        RECT 97.185 118.815 97.715 118.985 ;
        RECT 93.980 118.055 95.705 118.225 ;
        RECT 91.975 117.215 92.265 118.055 ;
        RECT 92.435 117.045 92.605 117.885 ;
        RECT 92.815 117.215 93.065 118.055 ;
        RECT 93.275 117.045 93.445 117.885 ;
        RECT 94.235 117.045 94.405 117.885 ;
        RECT 94.615 117.215 94.865 118.055 ;
        RECT 95.075 117.045 95.245 117.885 ;
        RECT 95.415 117.215 95.705 118.055 ;
        RECT 95.915 117.045 96.085 118.105 ;
        RECT 96.260 117.765 96.430 118.385 ;
        RECT 96.775 118.275 97.315 118.645 ;
        RECT 97.495 118.535 97.715 118.815 ;
        RECT 97.885 118.365 98.055 119.145 ;
        RECT 97.650 118.195 98.055 118.365 ;
        RECT 98.225 118.355 98.575 118.975 ;
        RECT 97.650 118.105 97.820 118.195 ;
        RECT 98.745 118.185 98.955 118.975 ;
        RECT 96.600 117.935 97.820 118.105 ;
        RECT 98.280 118.025 98.955 118.185 ;
        RECT 96.260 117.595 97.060 117.765 ;
        RECT 96.380 117.045 96.710 117.425 ;
        RECT 96.890 117.305 97.060 117.595 ;
        RECT 97.650 117.555 97.820 117.935 ;
        RECT 97.990 118.015 98.955 118.025 ;
        RECT 99.145 118.845 99.405 119.235 ;
        RECT 99.615 119.135 99.945 119.595 ;
        RECT 100.820 119.205 101.675 119.375 ;
        RECT 101.880 119.205 102.375 119.375 ;
        RECT 102.545 119.235 102.875 119.595 ;
        RECT 99.145 118.155 99.315 118.845 ;
        RECT 99.485 118.495 99.655 118.675 ;
        RECT 99.825 118.665 100.615 118.915 ;
        RECT 100.820 118.495 100.990 119.205 ;
        RECT 101.160 118.695 101.515 118.915 ;
        RECT 99.485 118.325 101.175 118.495 ;
        RECT 97.990 117.725 98.450 118.015 ;
        RECT 99.145 117.985 100.645 118.155 ;
        RECT 99.145 117.845 99.315 117.985 ;
        RECT 98.755 117.675 99.315 117.845 ;
        RECT 97.230 117.045 97.480 117.505 ;
        RECT 97.650 117.215 98.520 117.555 ;
        RECT 98.755 117.215 98.925 117.675 ;
        RECT 99.760 117.645 100.835 117.815 ;
        RECT 99.095 117.045 99.465 117.505 ;
        RECT 99.760 117.305 99.930 117.645 ;
        RECT 100.100 117.045 100.430 117.475 ;
        RECT 100.665 117.305 100.835 117.645 ;
        RECT 101.005 117.545 101.175 118.325 ;
        RECT 101.345 118.105 101.515 118.695 ;
        RECT 101.685 118.295 102.035 118.915 ;
        RECT 101.345 117.715 101.810 118.105 ;
        RECT 102.205 117.845 102.375 119.205 ;
        RECT 102.545 118.015 103.005 119.065 ;
        RECT 101.980 117.675 102.375 117.845 ;
        RECT 101.980 117.545 102.150 117.675 ;
        RECT 101.005 117.215 101.685 117.545 ;
        RECT 101.900 117.215 102.150 117.545 ;
        RECT 102.320 117.045 102.570 117.505 ;
        RECT 102.740 117.230 103.065 118.015 ;
        RECT 103.235 117.215 103.405 119.335 ;
        RECT 103.575 119.215 103.905 119.595 ;
        RECT 104.075 119.045 104.330 119.335 ;
        RECT 103.580 118.875 104.330 119.045 ;
        RECT 103.580 117.885 103.810 118.875 ;
        RECT 104.565 118.775 104.775 119.595 ;
        RECT 104.945 118.795 105.275 119.425 ;
        RECT 103.980 118.055 104.330 118.705 ;
        RECT 104.945 118.195 105.195 118.795 ;
        RECT 105.445 118.775 105.675 119.595 ;
        RECT 105.885 118.825 108.475 119.595 ;
        RECT 108.645 118.870 108.935 119.595 ;
        RECT 109.105 119.050 114.450 119.595 ;
        RECT 105.365 118.355 105.695 118.605 ;
        RECT 105.885 118.305 107.095 118.825 ;
        RECT 103.580 117.715 104.330 117.885 ;
        RECT 103.575 117.045 103.905 117.545 ;
        RECT 104.075 117.215 104.330 117.715 ;
        RECT 104.565 117.045 104.775 118.185 ;
        RECT 104.945 117.215 105.275 118.195 ;
        RECT 105.445 117.045 105.675 118.185 ;
        RECT 107.265 118.135 108.475 118.655 ;
        RECT 110.690 118.220 111.030 119.050 ;
        RECT 114.625 118.825 117.215 119.595 ;
        RECT 117.385 118.845 118.595 119.595 ;
        RECT 105.885 117.045 108.475 118.135 ;
        RECT 108.645 117.045 108.935 118.210 ;
        RECT 112.510 117.480 112.860 118.730 ;
        RECT 114.625 118.305 115.835 118.825 ;
        RECT 116.005 118.135 117.215 118.655 ;
        RECT 109.105 117.045 114.450 117.480 ;
        RECT 114.625 117.045 117.215 118.135 ;
        RECT 117.385 118.135 117.905 118.675 ;
        RECT 118.075 118.305 118.595 118.845 ;
        RECT 117.385 117.045 118.595 118.135 ;
        RECT 5.520 116.875 118.680 117.045 ;
        RECT 5.605 115.785 6.815 116.875 ;
        RECT 7.295 116.035 7.465 116.875 ;
        RECT 7.675 115.865 7.925 116.705 ;
        RECT 8.135 116.035 8.305 116.875 ;
        RECT 8.475 115.865 8.765 116.705 ;
        RECT 5.605 115.075 6.125 115.615 ;
        RECT 6.295 115.245 6.815 115.785 ;
        RECT 7.040 115.695 8.765 115.865 ;
        RECT 8.975 115.815 9.145 116.875 ;
        RECT 9.440 116.495 9.770 116.875 ;
        RECT 9.950 116.325 10.120 116.615 ;
        RECT 10.290 116.415 10.540 116.875 ;
        RECT 9.320 116.155 10.120 116.325 ;
        RECT 10.710 116.365 11.580 116.705 ;
        RECT 7.040 115.145 7.450 115.695 ;
        RECT 9.320 115.535 9.490 116.155 ;
        RECT 10.710 115.985 10.880 116.365 ;
        RECT 11.815 116.245 11.985 116.705 ;
        RECT 12.155 116.415 12.525 116.875 ;
        RECT 12.820 116.275 12.990 116.615 ;
        RECT 13.160 116.445 13.490 116.875 ;
        RECT 13.725 116.275 13.895 116.615 ;
        RECT 9.660 115.815 10.880 115.985 ;
        RECT 11.050 115.905 11.510 116.195 ;
        RECT 11.815 116.075 12.375 116.245 ;
        RECT 12.820 116.105 13.895 116.275 ;
        RECT 14.065 116.375 14.745 116.705 ;
        RECT 14.960 116.375 15.210 116.705 ;
        RECT 15.380 116.415 15.630 116.875 ;
        RECT 12.205 115.935 12.375 116.075 ;
        RECT 11.050 115.895 12.015 115.905 ;
        RECT 10.710 115.725 10.880 115.815 ;
        RECT 11.340 115.735 12.015 115.895 ;
        RECT 9.320 115.525 9.665 115.535 ;
        RECT 7.635 115.315 9.665 115.525 ;
        RECT 5.605 114.325 6.815 115.075 ;
        RECT 7.040 114.975 8.805 115.145 ;
        RECT 7.295 114.325 7.465 114.795 ;
        RECT 7.635 114.495 7.965 114.975 ;
        RECT 8.135 114.325 8.305 114.795 ;
        RECT 8.475 114.495 8.805 114.975 ;
        RECT 8.975 114.325 9.145 115.135 ;
        RECT 9.340 115.060 9.665 115.315 ;
        RECT 9.345 114.705 9.665 115.060 ;
        RECT 9.835 115.275 10.375 115.645 ;
        RECT 10.710 115.555 11.115 115.725 ;
        RECT 9.835 114.875 10.075 115.275 ;
        RECT 10.555 115.105 10.775 115.385 ;
        RECT 10.245 114.935 10.775 115.105 ;
        RECT 10.245 114.705 10.415 114.935 ;
        RECT 10.945 114.775 11.115 115.555 ;
        RECT 11.285 114.945 11.635 115.565 ;
        RECT 11.805 114.945 12.015 115.735 ;
        RECT 12.205 115.765 13.705 115.935 ;
        RECT 12.205 115.075 12.375 115.765 ;
        RECT 14.065 115.595 14.235 116.375 ;
        RECT 15.040 116.245 15.210 116.375 ;
        RECT 12.545 115.425 14.235 115.595 ;
        RECT 14.405 115.815 14.870 116.205 ;
        RECT 15.040 116.075 15.435 116.245 ;
        RECT 12.545 115.245 12.715 115.425 ;
        RECT 9.345 114.535 10.415 114.705 ;
        RECT 10.585 114.325 10.775 114.765 ;
        RECT 10.945 114.495 11.895 114.775 ;
        RECT 12.205 114.685 12.465 115.075 ;
        RECT 12.885 115.005 13.675 115.255 ;
        RECT 12.115 114.515 12.465 114.685 ;
        RECT 12.675 114.325 13.005 114.785 ;
        RECT 13.880 114.715 14.050 115.425 ;
        RECT 14.405 115.225 14.575 115.815 ;
        RECT 14.220 115.005 14.575 115.225 ;
        RECT 14.745 115.005 15.095 115.625 ;
        RECT 15.265 114.715 15.435 116.075 ;
        RECT 15.800 115.905 16.125 116.690 ;
        RECT 15.605 114.855 16.065 115.905 ;
        RECT 13.880 114.545 14.735 114.715 ;
        RECT 14.940 114.545 15.435 114.715 ;
        RECT 15.605 114.325 15.935 114.685 ;
        RECT 16.295 114.585 16.465 116.705 ;
        RECT 16.635 116.375 16.965 116.875 ;
        RECT 17.135 116.205 17.390 116.705 ;
        RECT 16.640 116.035 17.390 116.205 ;
        RECT 16.640 115.045 16.870 116.035 ;
        RECT 17.040 115.215 17.390 115.865 ;
        RECT 18.485 115.710 18.775 116.875 ;
        RECT 18.950 116.205 19.205 116.705 ;
        RECT 19.375 116.375 19.705 116.875 ;
        RECT 18.950 116.035 19.700 116.205 ;
        RECT 18.950 115.215 19.300 115.865 ;
        RECT 16.640 114.875 17.390 115.045 ;
        RECT 16.635 114.325 16.965 114.705 ;
        RECT 17.135 114.585 17.390 114.875 ;
        RECT 18.485 114.325 18.775 115.050 ;
        RECT 19.470 115.045 19.700 116.035 ;
        RECT 18.950 114.875 19.700 115.045 ;
        RECT 18.950 114.585 19.205 114.875 ;
        RECT 19.375 114.325 19.705 114.705 ;
        RECT 19.875 114.585 20.045 116.705 ;
        RECT 20.215 115.905 20.540 116.690 ;
        RECT 20.710 116.415 20.960 116.875 ;
        RECT 21.130 116.375 21.380 116.705 ;
        RECT 21.595 116.375 22.275 116.705 ;
        RECT 21.130 116.245 21.300 116.375 ;
        RECT 20.905 116.075 21.300 116.245 ;
        RECT 20.275 114.855 20.735 115.905 ;
        RECT 20.905 114.715 21.075 116.075 ;
        RECT 21.470 115.815 21.935 116.205 ;
        RECT 21.245 115.005 21.595 115.625 ;
        RECT 21.765 115.225 21.935 115.815 ;
        RECT 22.105 115.595 22.275 116.375 ;
        RECT 22.445 116.275 22.615 116.615 ;
        RECT 22.850 116.445 23.180 116.875 ;
        RECT 23.350 116.275 23.520 116.615 ;
        RECT 23.815 116.415 24.185 116.875 ;
        RECT 22.445 116.105 23.520 116.275 ;
        RECT 24.355 116.245 24.525 116.705 ;
        RECT 24.760 116.365 25.630 116.705 ;
        RECT 25.800 116.415 26.050 116.875 ;
        RECT 23.965 116.075 24.525 116.245 ;
        RECT 23.965 115.935 24.135 116.075 ;
        RECT 22.635 115.765 24.135 115.935 ;
        RECT 24.830 115.905 25.290 116.195 ;
        RECT 22.105 115.425 23.795 115.595 ;
        RECT 21.765 115.005 22.120 115.225 ;
        RECT 22.290 114.715 22.460 115.425 ;
        RECT 22.665 115.005 23.455 115.255 ;
        RECT 23.625 115.245 23.795 115.425 ;
        RECT 23.965 115.075 24.135 115.765 ;
        RECT 20.405 114.325 20.735 114.685 ;
        RECT 20.905 114.545 21.400 114.715 ;
        RECT 21.605 114.545 22.460 114.715 ;
        RECT 23.335 114.325 23.665 114.785 ;
        RECT 23.875 114.685 24.135 115.075 ;
        RECT 24.325 115.895 25.290 115.905 ;
        RECT 25.460 115.985 25.630 116.365 ;
        RECT 26.220 116.325 26.390 116.615 ;
        RECT 26.570 116.495 26.900 116.875 ;
        RECT 26.220 116.155 27.020 116.325 ;
        RECT 24.325 115.735 25.000 115.895 ;
        RECT 25.460 115.815 26.680 115.985 ;
        RECT 24.325 114.945 24.535 115.735 ;
        RECT 25.460 115.725 25.630 115.815 ;
        RECT 24.705 114.945 25.055 115.565 ;
        RECT 25.225 115.555 25.630 115.725 ;
        RECT 25.225 114.775 25.395 115.555 ;
        RECT 25.565 115.105 25.785 115.385 ;
        RECT 25.965 115.275 26.505 115.645 ;
        RECT 26.850 115.535 27.020 116.155 ;
        RECT 27.195 115.815 27.365 116.875 ;
        RECT 27.575 115.865 27.865 116.705 ;
        RECT 28.035 116.035 28.205 116.875 ;
        RECT 28.415 115.865 28.665 116.705 ;
        RECT 28.875 116.035 29.045 116.875 ;
        RECT 27.575 115.695 29.300 115.865 ;
        RECT 29.585 115.735 29.795 116.875 ;
        RECT 25.565 114.935 26.095 115.105 ;
        RECT 23.875 114.515 24.225 114.685 ;
        RECT 24.445 114.495 25.395 114.775 ;
        RECT 25.565 114.325 25.755 114.765 ;
        RECT 25.925 114.705 26.095 114.935 ;
        RECT 26.265 114.875 26.505 115.275 ;
        RECT 26.675 115.525 27.020 115.535 ;
        RECT 26.675 115.315 28.705 115.525 ;
        RECT 26.675 115.060 27.000 115.315 ;
        RECT 28.890 115.145 29.300 115.695 ;
        RECT 29.965 115.725 30.295 116.705 ;
        RECT 30.465 115.735 30.695 116.875 ;
        RECT 30.905 115.785 32.115 116.875 ;
        RECT 26.675 114.705 26.995 115.060 ;
        RECT 25.925 114.535 26.995 114.705 ;
        RECT 27.195 114.325 27.365 115.135 ;
        RECT 27.535 114.975 29.300 115.145 ;
        RECT 27.535 114.495 27.865 114.975 ;
        RECT 28.035 114.325 28.205 114.795 ;
        RECT 28.375 114.495 28.705 114.975 ;
        RECT 28.875 114.325 29.045 114.795 ;
        RECT 29.585 114.325 29.795 115.145 ;
        RECT 29.965 115.125 30.215 115.725 ;
        RECT 30.385 115.315 30.715 115.565 ;
        RECT 29.965 114.495 30.295 115.125 ;
        RECT 30.465 114.325 30.695 115.145 ;
        RECT 30.905 115.075 31.425 115.615 ;
        RECT 31.595 115.245 32.115 115.785 ;
        RECT 32.325 115.735 32.555 116.875 ;
        RECT 32.725 115.725 33.055 116.705 ;
        RECT 33.225 115.735 33.435 116.875 ;
        RECT 33.670 116.205 33.925 116.705 ;
        RECT 34.095 116.375 34.425 116.875 ;
        RECT 33.670 116.035 34.420 116.205 ;
        RECT 32.305 115.315 32.635 115.565 ;
        RECT 30.905 114.325 32.115 115.075 ;
        RECT 32.325 114.325 32.555 115.145 ;
        RECT 32.805 115.125 33.055 115.725 ;
        RECT 33.670 115.215 34.020 115.865 ;
        RECT 32.725 114.495 33.055 115.125 ;
        RECT 33.225 114.325 33.435 115.145 ;
        RECT 34.190 115.045 34.420 116.035 ;
        RECT 33.670 114.875 34.420 115.045 ;
        RECT 33.670 114.585 33.925 114.875 ;
        RECT 34.095 114.325 34.425 114.705 ;
        RECT 34.595 114.585 34.765 116.705 ;
        RECT 34.935 115.905 35.260 116.690 ;
        RECT 35.430 116.415 35.680 116.875 ;
        RECT 35.850 116.375 36.100 116.705 ;
        RECT 36.315 116.375 36.995 116.705 ;
        RECT 35.850 116.245 36.020 116.375 ;
        RECT 35.625 116.075 36.020 116.245 ;
        RECT 34.995 114.855 35.455 115.905 ;
        RECT 35.625 114.715 35.795 116.075 ;
        RECT 36.190 115.815 36.655 116.205 ;
        RECT 35.965 115.005 36.315 115.625 ;
        RECT 36.485 115.225 36.655 115.815 ;
        RECT 36.825 115.595 36.995 116.375 ;
        RECT 37.165 116.275 37.335 116.615 ;
        RECT 37.570 116.445 37.900 116.875 ;
        RECT 38.070 116.275 38.240 116.615 ;
        RECT 38.535 116.415 38.905 116.875 ;
        RECT 37.165 116.105 38.240 116.275 ;
        RECT 39.075 116.245 39.245 116.705 ;
        RECT 39.480 116.365 40.350 116.705 ;
        RECT 40.520 116.415 40.770 116.875 ;
        RECT 38.685 116.075 39.245 116.245 ;
        RECT 38.685 115.935 38.855 116.075 ;
        RECT 37.355 115.765 38.855 115.935 ;
        RECT 39.550 115.905 40.010 116.195 ;
        RECT 36.825 115.425 38.515 115.595 ;
        RECT 36.485 115.005 36.840 115.225 ;
        RECT 37.010 114.715 37.180 115.425 ;
        RECT 37.385 115.005 38.175 115.255 ;
        RECT 38.345 115.245 38.515 115.425 ;
        RECT 38.685 115.075 38.855 115.765 ;
        RECT 35.125 114.325 35.455 114.685 ;
        RECT 35.625 114.545 36.120 114.715 ;
        RECT 36.325 114.545 37.180 114.715 ;
        RECT 38.055 114.325 38.385 114.785 ;
        RECT 38.595 114.685 38.855 115.075 ;
        RECT 39.045 115.895 40.010 115.905 ;
        RECT 40.180 115.985 40.350 116.365 ;
        RECT 40.940 116.325 41.110 116.615 ;
        RECT 41.290 116.495 41.620 116.875 ;
        RECT 40.940 116.155 41.740 116.325 ;
        RECT 39.045 115.735 39.720 115.895 ;
        RECT 40.180 115.815 41.400 115.985 ;
        RECT 39.045 114.945 39.255 115.735 ;
        RECT 40.180 115.725 40.350 115.815 ;
        RECT 39.425 114.945 39.775 115.565 ;
        RECT 39.945 115.555 40.350 115.725 ;
        RECT 39.945 114.775 40.115 115.555 ;
        RECT 40.285 115.105 40.505 115.385 ;
        RECT 40.685 115.275 41.225 115.645 ;
        RECT 41.570 115.535 41.740 116.155 ;
        RECT 41.915 115.815 42.085 116.875 ;
        RECT 42.295 115.865 42.585 116.705 ;
        RECT 42.755 116.035 42.925 116.875 ;
        RECT 43.135 115.865 43.385 116.705 ;
        RECT 43.595 116.035 43.765 116.875 ;
        RECT 42.295 115.695 44.020 115.865 ;
        RECT 44.245 115.710 44.535 116.875 ;
        RECT 44.705 115.800 44.975 116.705 ;
        RECT 45.145 116.115 45.475 116.875 ;
        RECT 45.655 115.945 45.825 116.705 ;
        RECT 46.550 116.205 46.805 116.705 ;
        RECT 46.975 116.375 47.305 116.875 ;
        RECT 46.550 116.035 47.300 116.205 ;
        RECT 40.285 114.935 40.815 115.105 ;
        RECT 38.595 114.515 38.945 114.685 ;
        RECT 39.165 114.495 40.115 114.775 ;
        RECT 40.285 114.325 40.475 114.765 ;
        RECT 40.645 114.705 40.815 114.935 ;
        RECT 40.985 114.875 41.225 115.275 ;
        RECT 41.395 115.525 41.740 115.535 ;
        RECT 41.395 115.315 43.425 115.525 ;
        RECT 41.395 115.060 41.720 115.315 ;
        RECT 43.610 115.145 44.020 115.695 ;
        RECT 41.395 114.705 41.715 115.060 ;
        RECT 40.645 114.535 41.715 114.705 ;
        RECT 41.915 114.325 42.085 115.135 ;
        RECT 42.255 114.975 44.020 115.145 ;
        RECT 42.255 114.495 42.585 114.975 ;
        RECT 42.755 114.325 42.925 114.795 ;
        RECT 43.095 114.495 43.425 114.975 ;
        RECT 43.595 114.325 43.765 114.795 ;
        RECT 44.245 114.325 44.535 115.050 ;
        RECT 44.705 115.000 44.875 115.800 ;
        RECT 45.160 115.775 45.825 115.945 ;
        RECT 45.160 115.630 45.330 115.775 ;
        RECT 45.045 115.300 45.330 115.630 ;
        RECT 45.160 115.045 45.330 115.300 ;
        RECT 45.565 115.225 45.895 115.595 ;
        RECT 46.550 115.215 46.900 115.865 ;
        RECT 47.070 115.045 47.300 116.035 ;
        RECT 44.705 114.495 44.965 115.000 ;
        RECT 45.160 114.875 45.825 115.045 ;
        RECT 45.145 114.325 45.475 114.705 ;
        RECT 45.655 114.495 45.825 114.875 ;
        RECT 46.550 114.875 47.300 115.045 ;
        RECT 46.550 114.585 46.805 114.875 ;
        RECT 46.975 114.325 47.305 114.705 ;
        RECT 47.475 114.585 47.645 116.705 ;
        RECT 47.815 115.905 48.140 116.690 ;
        RECT 48.310 116.415 48.560 116.875 ;
        RECT 48.730 116.375 48.980 116.705 ;
        RECT 49.195 116.375 49.875 116.705 ;
        RECT 48.730 116.245 48.900 116.375 ;
        RECT 48.505 116.075 48.900 116.245 ;
        RECT 47.875 114.855 48.335 115.905 ;
        RECT 48.505 114.715 48.675 116.075 ;
        RECT 49.070 115.815 49.535 116.205 ;
        RECT 48.845 115.005 49.195 115.625 ;
        RECT 49.365 115.225 49.535 115.815 ;
        RECT 49.705 115.595 49.875 116.375 ;
        RECT 50.045 116.275 50.215 116.615 ;
        RECT 50.450 116.445 50.780 116.875 ;
        RECT 50.950 116.275 51.120 116.615 ;
        RECT 51.415 116.415 51.785 116.875 ;
        RECT 50.045 116.105 51.120 116.275 ;
        RECT 51.955 116.245 52.125 116.705 ;
        RECT 52.360 116.365 53.230 116.705 ;
        RECT 53.400 116.415 53.650 116.875 ;
        RECT 51.565 116.075 52.125 116.245 ;
        RECT 51.565 115.935 51.735 116.075 ;
        RECT 50.235 115.765 51.735 115.935 ;
        RECT 52.430 115.905 52.890 116.195 ;
        RECT 49.705 115.425 51.395 115.595 ;
        RECT 49.365 115.005 49.720 115.225 ;
        RECT 49.890 114.715 50.060 115.425 ;
        RECT 50.265 115.005 51.055 115.255 ;
        RECT 51.225 115.245 51.395 115.425 ;
        RECT 51.565 115.075 51.735 115.765 ;
        RECT 48.005 114.325 48.335 114.685 ;
        RECT 48.505 114.545 49.000 114.715 ;
        RECT 49.205 114.545 50.060 114.715 ;
        RECT 50.935 114.325 51.265 114.785 ;
        RECT 51.475 114.685 51.735 115.075 ;
        RECT 51.925 115.895 52.890 115.905 ;
        RECT 53.060 115.985 53.230 116.365 ;
        RECT 53.820 116.325 53.990 116.615 ;
        RECT 54.170 116.495 54.500 116.875 ;
        RECT 53.820 116.155 54.620 116.325 ;
        RECT 51.925 115.735 52.600 115.895 ;
        RECT 53.060 115.815 54.280 115.985 ;
        RECT 51.925 114.945 52.135 115.735 ;
        RECT 53.060 115.725 53.230 115.815 ;
        RECT 52.305 114.945 52.655 115.565 ;
        RECT 52.825 115.555 53.230 115.725 ;
        RECT 52.825 114.775 52.995 115.555 ;
        RECT 53.165 115.105 53.385 115.385 ;
        RECT 53.565 115.275 54.105 115.645 ;
        RECT 54.450 115.535 54.620 116.155 ;
        RECT 54.795 115.815 54.965 116.875 ;
        RECT 55.175 115.865 55.465 116.705 ;
        RECT 55.635 116.035 55.805 116.875 ;
        RECT 56.015 115.865 56.265 116.705 ;
        RECT 56.475 116.035 56.645 116.875 ;
        RECT 55.175 115.695 56.900 115.865 ;
        RECT 53.165 114.935 53.695 115.105 ;
        RECT 51.475 114.515 51.825 114.685 ;
        RECT 52.045 114.495 52.995 114.775 ;
        RECT 53.165 114.325 53.355 114.765 ;
        RECT 53.525 114.705 53.695 114.935 ;
        RECT 53.865 114.875 54.105 115.275 ;
        RECT 54.275 115.525 54.620 115.535 ;
        RECT 54.275 115.315 56.305 115.525 ;
        RECT 54.275 115.060 54.600 115.315 ;
        RECT 56.490 115.145 56.900 115.695 ;
        RECT 54.275 114.705 54.595 115.060 ;
        RECT 53.525 114.535 54.595 114.705 ;
        RECT 54.795 114.325 54.965 115.135 ;
        RECT 55.135 114.975 56.900 115.145 ;
        RECT 57.125 115.800 57.395 116.705 ;
        RECT 57.565 116.115 57.895 116.875 ;
        RECT 58.075 115.945 58.245 116.705 ;
        RECT 59.430 116.205 59.685 116.705 ;
        RECT 59.855 116.375 60.185 116.875 ;
        RECT 59.430 116.035 60.180 116.205 ;
        RECT 57.125 115.000 57.295 115.800 ;
        RECT 57.580 115.775 58.245 115.945 ;
        RECT 57.580 115.630 57.750 115.775 ;
        RECT 57.465 115.300 57.750 115.630 ;
        RECT 57.580 115.045 57.750 115.300 ;
        RECT 57.985 115.225 58.315 115.595 ;
        RECT 59.430 115.215 59.780 115.865 ;
        RECT 59.950 115.045 60.180 116.035 ;
        RECT 55.135 114.495 55.465 114.975 ;
        RECT 55.635 114.325 55.805 114.795 ;
        RECT 55.975 114.495 56.305 114.975 ;
        RECT 56.475 114.325 56.645 114.795 ;
        RECT 57.125 114.495 57.385 115.000 ;
        RECT 57.580 114.875 58.245 115.045 ;
        RECT 57.565 114.325 57.895 114.705 ;
        RECT 58.075 114.495 58.245 114.875 ;
        RECT 59.430 114.875 60.180 115.045 ;
        RECT 59.430 114.585 59.685 114.875 ;
        RECT 59.855 114.325 60.185 114.705 ;
        RECT 60.355 114.585 60.525 116.705 ;
        RECT 60.695 115.905 61.020 116.690 ;
        RECT 61.190 116.415 61.440 116.875 ;
        RECT 61.610 116.375 61.860 116.705 ;
        RECT 62.075 116.375 62.755 116.705 ;
        RECT 61.610 116.245 61.780 116.375 ;
        RECT 61.385 116.075 61.780 116.245 ;
        RECT 60.755 114.855 61.215 115.905 ;
        RECT 61.385 114.715 61.555 116.075 ;
        RECT 61.950 115.815 62.415 116.205 ;
        RECT 61.725 115.005 62.075 115.625 ;
        RECT 62.245 115.225 62.415 115.815 ;
        RECT 62.585 115.595 62.755 116.375 ;
        RECT 62.925 116.275 63.095 116.615 ;
        RECT 63.330 116.445 63.660 116.875 ;
        RECT 63.830 116.275 64.000 116.615 ;
        RECT 64.295 116.415 64.665 116.875 ;
        RECT 62.925 116.105 64.000 116.275 ;
        RECT 64.835 116.245 65.005 116.705 ;
        RECT 65.240 116.365 66.110 116.705 ;
        RECT 66.280 116.415 66.530 116.875 ;
        RECT 64.445 116.075 65.005 116.245 ;
        RECT 64.445 115.935 64.615 116.075 ;
        RECT 63.115 115.765 64.615 115.935 ;
        RECT 65.310 115.905 65.770 116.195 ;
        RECT 62.585 115.425 64.275 115.595 ;
        RECT 62.245 115.005 62.600 115.225 ;
        RECT 62.770 114.715 62.940 115.425 ;
        RECT 63.145 115.005 63.935 115.255 ;
        RECT 64.105 115.245 64.275 115.425 ;
        RECT 64.445 115.075 64.615 115.765 ;
        RECT 60.885 114.325 61.215 114.685 ;
        RECT 61.385 114.545 61.880 114.715 ;
        RECT 62.085 114.545 62.940 114.715 ;
        RECT 63.815 114.325 64.145 114.785 ;
        RECT 64.355 114.685 64.615 115.075 ;
        RECT 64.805 115.895 65.770 115.905 ;
        RECT 65.940 115.985 66.110 116.365 ;
        RECT 66.700 116.325 66.870 116.615 ;
        RECT 67.050 116.495 67.380 116.875 ;
        RECT 66.700 116.155 67.500 116.325 ;
        RECT 64.805 115.735 65.480 115.895 ;
        RECT 65.940 115.815 67.160 115.985 ;
        RECT 64.805 114.945 65.015 115.735 ;
        RECT 65.940 115.725 66.110 115.815 ;
        RECT 65.185 114.945 65.535 115.565 ;
        RECT 65.705 115.555 66.110 115.725 ;
        RECT 65.705 114.775 65.875 115.555 ;
        RECT 66.045 115.105 66.265 115.385 ;
        RECT 66.445 115.275 66.985 115.645 ;
        RECT 67.330 115.535 67.500 116.155 ;
        RECT 67.675 115.815 67.845 116.875 ;
        RECT 68.055 115.865 68.345 116.705 ;
        RECT 68.515 116.035 68.685 116.875 ;
        RECT 68.895 115.865 69.145 116.705 ;
        RECT 69.355 116.035 69.525 116.875 ;
        RECT 68.055 115.695 69.780 115.865 ;
        RECT 70.005 115.710 70.295 116.875 ;
        RECT 70.465 115.800 70.735 116.705 ;
        RECT 70.905 116.115 71.235 116.875 ;
        RECT 71.415 115.945 71.585 116.705 ;
        RECT 66.045 114.935 66.575 115.105 ;
        RECT 64.355 114.515 64.705 114.685 ;
        RECT 64.925 114.495 65.875 114.775 ;
        RECT 66.045 114.325 66.235 114.765 ;
        RECT 66.405 114.705 66.575 114.935 ;
        RECT 66.745 114.875 66.985 115.275 ;
        RECT 67.155 115.525 67.500 115.535 ;
        RECT 67.155 115.315 69.185 115.525 ;
        RECT 67.155 115.060 67.480 115.315 ;
        RECT 69.370 115.145 69.780 115.695 ;
        RECT 67.155 114.705 67.475 115.060 ;
        RECT 66.405 114.535 67.475 114.705 ;
        RECT 67.675 114.325 67.845 115.135 ;
        RECT 68.015 114.975 69.780 115.145 ;
        RECT 68.015 114.495 68.345 114.975 ;
        RECT 68.515 114.325 68.685 114.795 ;
        RECT 68.855 114.495 69.185 114.975 ;
        RECT 69.355 114.325 69.525 114.795 ;
        RECT 70.005 114.325 70.295 115.050 ;
        RECT 70.465 115.000 70.635 115.800 ;
        RECT 70.920 115.775 71.585 115.945 ;
        RECT 70.920 115.630 71.090 115.775 ;
        RECT 71.905 115.735 72.115 116.875 ;
        RECT 70.805 115.300 71.090 115.630 ;
        RECT 72.285 115.725 72.615 116.705 ;
        RECT 72.785 115.735 73.015 116.875 ;
        RECT 73.225 115.785 74.435 116.875 ;
        RECT 70.920 115.045 71.090 115.300 ;
        RECT 71.325 115.225 71.655 115.595 ;
        RECT 70.465 114.495 70.725 115.000 ;
        RECT 70.920 114.875 71.585 115.045 ;
        RECT 70.905 114.325 71.235 114.705 ;
        RECT 71.415 114.495 71.585 114.875 ;
        RECT 71.905 114.325 72.115 115.145 ;
        RECT 72.285 115.125 72.535 115.725 ;
        RECT 72.705 115.315 73.035 115.565 ;
        RECT 72.285 114.495 72.615 115.125 ;
        RECT 72.785 114.325 73.015 115.145 ;
        RECT 73.225 115.075 73.745 115.615 ;
        RECT 73.915 115.245 74.435 115.785 ;
        RECT 74.645 115.735 74.875 116.875 ;
        RECT 75.045 115.725 75.375 116.705 ;
        RECT 75.545 115.735 75.755 116.875 ;
        RECT 75.990 116.205 76.245 116.705 ;
        RECT 76.415 116.375 76.745 116.875 ;
        RECT 75.990 116.035 76.740 116.205 ;
        RECT 74.625 115.315 74.955 115.565 ;
        RECT 73.225 114.325 74.435 115.075 ;
        RECT 74.645 114.325 74.875 115.145 ;
        RECT 75.125 115.125 75.375 115.725 ;
        RECT 75.990 115.215 76.340 115.865 ;
        RECT 75.045 114.495 75.375 115.125 ;
        RECT 75.545 114.325 75.755 115.145 ;
        RECT 76.510 115.045 76.740 116.035 ;
        RECT 75.990 114.875 76.740 115.045 ;
        RECT 75.990 114.585 76.245 114.875 ;
        RECT 76.415 114.325 76.745 114.705 ;
        RECT 76.915 114.585 77.085 116.705 ;
        RECT 77.255 115.905 77.580 116.690 ;
        RECT 77.750 116.415 78.000 116.875 ;
        RECT 78.170 116.375 78.420 116.705 ;
        RECT 78.635 116.375 79.315 116.705 ;
        RECT 78.170 116.245 78.340 116.375 ;
        RECT 77.945 116.075 78.340 116.245 ;
        RECT 77.315 114.855 77.775 115.905 ;
        RECT 77.945 114.715 78.115 116.075 ;
        RECT 78.510 115.815 78.975 116.205 ;
        RECT 78.285 115.005 78.635 115.625 ;
        RECT 78.805 115.225 78.975 115.815 ;
        RECT 79.145 115.595 79.315 116.375 ;
        RECT 79.485 116.275 79.655 116.615 ;
        RECT 79.890 116.445 80.220 116.875 ;
        RECT 80.390 116.275 80.560 116.615 ;
        RECT 80.855 116.415 81.225 116.875 ;
        RECT 79.485 116.105 80.560 116.275 ;
        RECT 81.395 116.245 81.565 116.705 ;
        RECT 81.800 116.365 82.670 116.705 ;
        RECT 82.840 116.415 83.090 116.875 ;
        RECT 81.005 116.075 81.565 116.245 ;
        RECT 81.005 115.935 81.175 116.075 ;
        RECT 79.675 115.765 81.175 115.935 ;
        RECT 81.870 115.905 82.330 116.195 ;
        RECT 79.145 115.425 80.835 115.595 ;
        RECT 78.805 115.005 79.160 115.225 ;
        RECT 79.330 114.715 79.500 115.425 ;
        RECT 79.705 115.005 80.495 115.255 ;
        RECT 80.665 115.245 80.835 115.425 ;
        RECT 81.005 115.075 81.175 115.765 ;
        RECT 77.445 114.325 77.775 114.685 ;
        RECT 77.945 114.545 78.440 114.715 ;
        RECT 78.645 114.545 79.500 114.715 ;
        RECT 80.375 114.325 80.705 114.785 ;
        RECT 80.915 114.685 81.175 115.075 ;
        RECT 81.365 115.895 82.330 115.905 ;
        RECT 82.500 115.985 82.670 116.365 ;
        RECT 83.260 116.325 83.430 116.615 ;
        RECT 83.610 116.495 83.940 116.875 ;
        RECT 83.260 116.155 84.060 116.325 ;
        RECT 81.365 115.735 82.040 115.895 ;
        RECT 82.500 115.815 83.720 115.985 ;
        RECT 81.365 114.945 81.575 115.735 ;
        RECT 82.500 115.725 82.670 115.815 ;
        RECT 81.745 114.945 82.095 115.565 ;
        RECT 82.265 115.555 82.670 115.725 ;
        RECT 82.265 114.775 82.435 115.555 ;
        RECT 82.605 115.105 82.825 115.385 ;
        RECT 83.005 115.275 83.545 115.645 ;
        RECT 83.890 115.535 84.060 116.155 ;
        RECT 84.235 115.815 84.405 116.875 ;
        RECT 84.615 115.865 84.905 116.705 ;
        RECT 85.075 116.035 85.245 116.875 ;
        RECT 85.455 115.865 85.705 116.705 ;
        RECT 85.915 116.035 86.085 116.875 ;
        RECT 84.615 115.695 86.340 115.865 ;
        RECT 82.605 114.935 83.135 115.105 ;
        RECT 80.915 114.515 81.265 114.685 ;
        RECT 81.485 114.495 82.435 114.775 ;
        RECT 82.605 114.325 82.795 114.765 ;
        RECT 82.965 114.705 83.135 114.935 ;
        RECT 83.305 114.875 83.545 115.275 ;
        RECT 83.715 115.525 84.060 115.535 ;
        RECT 83.715 115.315 85.745 115.525 ;
        RECT 83.715 115.060 84.040 115.315 ;
        RECT 85.930 115.145 86.340 115.695 ;
        RECT 83.715 114.705 84.035 115.060 ;
        RECT 82.965 114.535 84.035 114.705 ;
        RECT 84.235 114.325 84.405 115.135 ;
        RECT 84.575 114.975 86.340 115.145 ;
        RECT 86.565 115.800 86.835 116.705 ;
        RECT 87.005 116.115 87.335 116.875 ;
        RECT 87.515 115.945 87.685 116.705 ;
        RECT 86.565 115.000 86.735 115.800 ;
        RECT 87.020 115.775 87.685 115.945 ;
        RECT 87.020 115.630 87.190 115.775 ;
        RECT 87.985 115.735 88.215 116.875 ;
        RECT 88.385 115.725 88.715 116.705 ;
        RECT 88.885 115.735 89.095 116.875 ;
        RECT 89.875 115.945 90.045 116.705 ;
        RECT 90.225 116.115 90.555 116.875 ;
        RECT 89.875 115.775 90.540 115.945 ;
        RECT 90.725 115.800 90.995 116.705 ;
        RECT 86.905 115.300 87.190 115.630 ;
        RECT 87.020 115.045 87.190 115.300 ;
        RECT 87.425 115.225 87.755 115.595 ;
        RECT 87.965 115.315 88.295 115.565 ;
        RECT 84.575 114.495 84.905 114.975 ;
        RECT 85.075 114.325 85.245 114.795 ;
        RECT 85.415 114.495 85.745 114.975 ;
        RECT 85.915 114.325 86.085 114.795 ;
        RECT 86.565 114.495 86.825 115.000 ;
        RECT 87.020 114.875 87.685 115.045 ;
        RECT 87.005 114.325 87.335 114.705 ;
        RECT 87.515 114.495 87.685 114.875 ;
        RECT 87.985 114.325 88.215 115.145 ;
        RECT 88.465 115.125 88.715 115.725 ;
        RECT 90.370 115.630 90.540 115.775 ;
        RECT 89.805 115.225 90.135 115.595 ;
        RECT 90.370 115.300 90.655 115.630 ;
        RECT 88.385 114.495 88.715 115.125 ;
        RECT 88.885 114.325 89.095 115.145 ;
        RECT 90.370 115.045 90.540 115.300 ;
        RECT 89.875 114.875 90.540 115.045 ;
        RECT 90.825 115.000 90.995 115.800 ;
        RECT 91.165 115.785 92.375 116.875 ;
        RECT 89.875 114.495 90.045 114.875 ;
        RECT 90.225 114.325 90.555 114.705 ;
        RECT 90.735 114.495 90.995 115.000 ;
        RECT 91.165 115.075 91.685 115.615 ;
        RECT 91.855 115.245 92.375 115.785 ;
        RECT 92.585 115.735 92.815 116.875 ;
        RECT 92.985 115.725 93.315 116.705 ;
        RECT 93.485 115.735 93.695 116.875 ;
        RECT 94.475 115.945 94.645 116.705 ;
        RECT 94.825 116.115 95.155 116.875 ;
        RECT 94.475 115.775 95.140 115.945 ;
        RECT 95.325 115.800 95.595 116.705 ;
        RECT 92.565 115.315 92.895 115.565 ;
        RECT 91.165 114.325 92.375 115.075 ;
        RECT 92.585 114.325 92.815 115.145 ;
        RECT 93.065 115.125 93.315 115.725 ;
        RECT 94.970 115.630 95.140 115.775 ;
        RECT 94.405 115.225 94.735 115.595 ;
        RECT 94.970 115.300 95.255 115.630 ;
        RECT 92.985 114.495 93.315 115.125 ;
        RECT 93.485 114.325 93.695 115.145 ;
        RECT 94.970 115.045 95.140 115.300 ;
        RECT 94.475 114.875 95.140 115.045 ;
        RECT 95.425 115.000 95.595 115.800 ;
        RECT 95.765 115.710 96.055 116.875 ;
        RECT 96.230 116.205 96.485 116.705 ;
        RECT 96.655 116.375 96.985 116.875 ;
        RECT 96.230 116.035 96.980 116.205 ;
        RECT 96.230 115.215 96.580 115.865 ;
        RECT 94.475 114.495 94.645 114.875 ;
        RECT 94.825 114.325 95.155 114.705 ;
        RECT 95.335 114.495 95.595 115.000 ;
        RECT 95.765 114.325 96.055 115.050 ;
        RECT 96.750 115.045 96.980 116.035 ;
        RECT 96.230 114.875 96.980 115.045 ;
        RECT 96.230 114.585 96.485 114.875 ;
        RECT 96.655 114.325 96.985 114.705 ;
        RECT 97.155 114.585 97.325 116.705 ;
        RECT 97.495 115.905 97.820 116.690 ;
        RECT 97.990 116.415 98.240 116.875 ;
        RECT 98.410 116.375 98.660 116.705 ;
        RECT 98.875 116.375 99.555 116.705 ;
        RECT 98.410 116.245 98.580 116.375 ;
        RECT 98.185 116.075 98.580 116.245 ;
        RECT 97.555 114.855 98.015 115.905 ;
        RECT 98.185 114.715 98.355 116.075 ;
        RECT 98.750 115.815 99.215 116.205 ;
        RECT 98.525 115.005 98.875 115.625 ;
        RECT 99.045 115.225 99.215 115.815 ;
        RECT 99.385 115.595 99.555 116.375 ;
        RECT 99.725 116.275 99.895 116.615 ;
        RECT 100.130 116.445 100.460 116.875 ;
        RECT 100.630 116.275 100.800 116.615 ;
        RECT 101.095 116.415 101.465 116.875 ;
        RECT 99.725 116.105 100.800 116.275 ;
        RECT 101.635 116.245 101.805 116.705 ;
        RECT 102.040 116.365 102.910 116.705 ;
        RECT 103.080 116.415 103.330 116.875 ;
        RECT 101.245 116.075 101.805 116.245 ;
        RECT 101.245 115.935 101.415 116.075 ;
        RECT 99.915 115.765 101.415 115.935 ;
        RECT 102.110 115.905 102.570 116.195 ;
        RECT 99.385 115.425 101.075 115.595 ;
        RECT 99.045 115.005 99.400 115.225 ;
        RECT 99.570 114.715 99.740 115.425 ;
        RECT 99.945 115.005 100.735 115.255 ;
        RECT 100.905 115.245 101.075 115.425 ;
        RECT 101.245 115.075 101.415 115.765 ;
        RECT 97.685 114.325 98.015 114.685 ;
        RECT 98.185 114.545 98.680 114.715 ;
        RECT 98.885 114.545 99.740 114.715 ;
        RECT 100.615 114.325 100.945 114.785 ;
        RECT 101.155 114.685 101.415 115.075 ;
        RECT 101.605 115.895 102.570 115.905 ;
        RECT 102.740 115.985 102.910 116.365 ;
        RECT 103.500 116.325 103.670 116.615 ;
        RECT 103.850 116.495 104.180 116.875 ;
        RECT 103.500 116.155 104.300 116.325 ;
        RECT 101.605 115.735 102.280 115.895 ;
        RECT 102.740 115.815 103.960 115.985 ;
        RECT 101.605 114.945 101.815 115.735 ;
        RECT 102.740 115.725 102.910 115.815 ;
        RECT 101.985 114.945 102.335 115.565 ;
        RECT 102.505 115.555 102.910 115.725 ;
        RECT 102.505 114.775 102.675 115.555 ;
        RECT 102.845 115.105 103.065 115.385 ;
        RECT 103.245 115.275 103.785 115.645 ;
        RECT 104.130 115.535 104.300 116.155 ;
        RECT 104.475 115.815 104.645 116.875 ;
        RECT 104.855 115.865 105.145 116.705 ;
        RECT 105.315 116.035 105.485 116.875 ;
        RECT 105.695 115.865 105.945 116.705 ;
        RECT 106.155 116.035 106.325 116.875 ;
        RECT 106.810 116.205 107.065 116.705 ;
        RECT 107.235 116.375 107.565 116.875 ;
        RECT 106.810 116.035 107.560 116.205 ;
        RECT 104.855 115.695 106.580 115.865 ;
        RECT 102.845 114.935 103.375 115.105 ;
        RECT 101.155 114.515 101.505 114.685 ;
        RECT 101.725 114.495 102.675 114.775 ;
        RECT 102.845 114.325 103.035 114.765 ;
        RECT 103.205 114.705 103.375 114.935 ;
        RECT 103.545 114.875 103.785 115.275 ;
        RECT 103.955 115.525 104.300 115.535 ;
        RECT 103.955 115.315 105.985 115.525 ;
        RECT 103.955 115.060 104.280 115.315 ;
        RECT 106.170 115.145 106.580 115.695 ;
        RECT 106.810 115.215 107.160 115.865 ;
        RECT 103.955 114.705 104.275 115.060 ;
        RECT 103.205 114.535 104.275 114.705 ;
        RECT 104.475 114.325 104.645 115.135 ;
        RECT 104.815 114.975 106.580 115.145 ;
        RECT 107.330 115.045 107.560 116.035 ;
        RECT 104.815 114.495 105.145 114.975 ;
        RECT 105.315 114.325 105.485 114.795 ;
        RECT 105.655 114.495 105.985 114.975 ;
        RECT 106.810 114.875 107.560 115.045 ;
        RECT 106.155 114.325 106.325 114.795 ;
        RECT 106.810 114.585 107.065 114.875 ;
        RECT 107.235 114.325 107.565 114.705 ;
        RECT 107.735 114.585 107.905 116.705 ;
        RECT 108.075 115.905 108.400 116.690 ;
        RECT 108.570 116.415 108.820 116.875 ;
        RECT 108.990 116.375 109.240 116.705 ;
        RECT 109.455 116.375 110.135 116.705 ;
        RECT 108.990 116.245 109.160 116.375 ;
        RECT 108.765 116.075 109.160 116.245 ;
        RECT 108.135 114.855 108.595 115.905 ;
        RECT 108.765 114.715 108.935 116.075 ;
        RECT 109.330 115.815 109.795 116.205 ;
        RECT 109.105 115.005 109.455 115.625 ;
        RECT 109.625 115.225 109.795 115.815 ;
        RECT 109.965 115.595 110.135 116.375 ;
        RECT 110.305 116.275 110.475 116.615 ;
        RECT 110.710 116.445 111.040 116.875 ;
        RECT 111.210 116.275 111.380 116.615 ;
        RECT 111.675 116.415 112.045 116.875 ;
        RECT 110.305 116.105 111.380 116.275 ;
        RECT 112.215 116.245 112.385 116.705 ;
        RECT 112.620 116.365 113.490 116.705 ;
        RECT 113.660 116.415 113.910 116.875 ;
        RECT 111.825 116.075 112.385 116.245 ;
        RECT 111.825 115.935 111.995 116.075 ;
        RECT 110.495 115.765 111.995 115.935 ;
        RECT 112.690 115.905 113.150 116.195 ;
        RECT 109.965 115.425 111.655 115.595 ;
        RECT 109.625 115.005 109.980 115.225 ;
        RECT 110.150 114.715 110.320 115.425 ;
        RECT 110.525 115.005 111.315 115.255 ;
        RECT 111.485 115.245 111.655 115.425 ;
        RECT 111.825 115.075 111.995 115.765 ;
        RECT 108.265 114.325 108.595 114.685 ;
        RECT 108.765 114.545 109.260 114.715 ;
        RECT 109.465 114.545 110.320 114.715 ;
        RECT 111.195 114.325 111.525 114.785 ;
        RECT 111.735 114.685 111.995 115.075 ;
        RECT 112.185 115.895 113.150 115.905 ;
        RECT 113.320 115.985 113.490 116.365 ;
        RECT 114.080 116.325 114.250 116.615 ;
        RECT 114.430 116.495 114.760 116.875 ;
        RECT 114.080 116.155 114.880 116.325 ;
        RECT 112.185 115.735 112.860 115.895 ;
        RECT 113.320 115.815 114.540 115.985 ;
        RECT 112.185 114.945 112.395 115.735 ;
        RECT 113.320 115.725 113.490 115.815 ;
        RECT 112.565 114.945 112.915 115.565 ;
        RECT 113.085 115.555 113.490 115.725 ;
        RECT 113.085 114.775 113.255 115.555 ;
        RECT 113.425 115.105 113.645 115.385 ;
        RECT 113.825 115.275 114.365 115.645 ;
        RECT 114.710 115.535 114.880 116.155 ;
        RECT 115.055 115.815 115.225 116.875 ;
        RECT 115.435 115.865 115.725 116.705 ;
        RECT 115.895 116.035 116.065 116.875 ;
        RECT 116.275 115.865 116.525 116.705 ;
        RECT 116.735 116.035 116.905 116.875 ;
        RECT 115.435 115.695 117.160 115.865 ;
        RECT 113.425 114.935 113.955 115.105 ;
        RECT 111.735 114.515 112.085 114.685 ;
        RECT 112.305 114.495 113.255 114.775 ;
        RECT 113.425 114.325 113.615 114.765 ;
        RECT 113.785 114.705 113.955 114.935 ;
        RECT 114.125 114.875 114.365 115.275 ;
        RECT 114.535 115.525 114.880 115.535 ;
        RECT 114.535 115.315 116.565 115.525 ;
        RECT 114.535 115.060 114.860 115.315 ;
        RECT 116.750 115.145 117.160 115.695 ;
        RECT 117.385 115.785 118.595 116.875 ;
        RECT 117.385 115.245 117.905 115.785 ;
        RECT 114.535 114.705 114.855 115.060 ;
        RECT 113.785 114.535 114.855 114.705 ;
        RECT 115.055 114.325 115.225 115.135 ;
        RECT 115.395 114.975 117.160 115.145 ;
        RECT 118.075 115.075 118.595 115.615 ;
        RECT 115.395 114.495 115.725 114.975 ;
        RECT 115.895 114.325 116.065 114.795 ;
        RECT 116.235 114.495 116.565 114.975 ;
        RECT 116.735 114.325 116.905 114.795 ;
        RECT 117.385 114.325 118.595 115.075 ;
        RECT 5.520 114.155 118.680 114.325 ;
        RECT 5.605 113.405 6.815 114.155 ;
        RECT 7.295 113.685 7.465 114.155 ;
        RECT 7.635 113.505 7.965 113.985 ;
        RECT 8.135 113.685 8.305 114.155 ;
        RECT 8.475 113.505 8.805 113.985 ;
        RECT 5.605 112.865 6.125 113.405 ;
        RECT 7.040 113.335 8.805 113.505 ;
        RECT 8.975 113.345 9.145 114.155 ;
        RECT 9.345 113.775 10.415 113.945 ;
        RECT 9.345 113.420 9.665 113.775 ;
        RECT 6.295 112.695 6.815 113.235 ;
        RECT 5.605 111.605 6.815 112.695 ;
        RECT 7.040 112.785 7.450 113.335 ;
        RECT 9.340 113.165 9.665 113.420 ;
        RECT 7.635 112.955 9.665 113.165 ;
        RECT 9.320 112.945 9.665 112.955 ;
        RECT 9.835 113.205 10.075 113.605 ;
        RECT 10.245 113.545 10.415 113.775 ;
        RECT 10.585 113.715 10.775 114.155 ;
        RECT 10.945 113.705 11.895 113.985 ;
        RECT 12.115 113.795 12.465 113.965 ;
        RECT 10.245 113.375 10.775 113.545 ;
        RECT 7.040 112.615 8.765 112.785 ;
        RECT 7.295 111.605 7.465 112.445 ;
        RECT 7.675 111.775 7.925 112.615 ;
        RECT 8.135 111.605 8.305 112.445 ;
        RECT 8.475 111.775 8.765 112.615 ;
        RECT 8.975 111.605 9.145 112.665 ;
        RECT 9.320 112.325 9.490 112.945 ;
        RECT 9.835 112.835 10.375 113.205 ;
        RECT 10.555 113.095 10.775 113.375 ;
        RECT 10.945 112.925 11.115 113.705 ;
        RECT 10.710 112.755 11.115 112.925 ;
        RECT 11.285 112.915 11.635 113.535 ;
        RECT 10.710 112.665 10.880 112.755 ;
        RECT 11.805 112.745 12.015 113.535 ;
        RECT 9.660 112.495 10.880 112.665 ;
        RECT 11.340 112.585 12.015 112.745 ;
        RECT 9.320 112.155 10.120 112.325 ;
        RECT 9.440 111.605 9.770 111.985 ;
        RECT 9.950 111.865 10.120 112.155 ;
        RECT 10.710 112.115 10.880 112.495 ;
        RECT 11.050 112.575 12.015 112.585 ;
        RECT 12.205 113.405 12.465 113.795 ;
        RECT 12.675 113.695 13.005 114.155 ;
        RECT 13.880 113.765 14.735 113.935 ;
        RECT 14.940 113.765 15.435 113.935 ;
        RECT 15.605 113.795 15.935 114.155 ;
        RECT 12.205 112.715 12.375 113.405 ;
        RECT 12.545 113.055 12.715 113.235 ;
        RECT 12.885 113.225 13.675 113.475 ;
        RECT 13.880 113.055 14.050 113.765 ;
        RECT 14.220 113.255 14.575 113.475 ;
        RECT 12.545 112.885 14.235 113.055 ;
        RECT 11.050 112.285 11.510 112.575 ;
        RECT 12.205 112.545 13.705 112.715 ;
        RECT 12.205 112.405 12.375 112.545 ;
        RECT 11.815 112.235 12.375 112.405 ;
        RECT 10.290 111.605 10.540 112.065 ;
        RECT 10.710 111.775 11.580 112.115 ;
        RECT 11.815 111.775 11.985 112.235 ;
        RECT 12.820 112.205 13.895 112.375 ;
        RECT 12.155 111.605 12.525 112.065 ;
        RECT 12.820 111.865 12.990 112.205 ;
        RECT 13.160 111.605 13.490 112.035 ;
        RECT 13.725 111.865 13.895 112.205 ;
        RECT 14.065 112.105 14.235 112.885 ;
        RECT 14.405 112.665 14.575 113.255 ;
        RECT 14.745 112.855 15.095 113.475 ;
        RECT 14.405 112.275 14.870 112.665 ;
        RECT 15.265 112.405 15.435 113.765 ;
        RECT 15.605 112.575 16.065 113.625 ;
        RECT 15.040 112.235 15.435 112.405 ;
        RECT 15.040 112.105 15.210 112.235 ;
        RECT 14.065 111.775 14.745 112.105 ;
        RECT 14.960 111.775 15.210 112.105 ;
        RECT 15.380 111.605 15.630 112.065 ;
        RECT 15.800 111.790 16.125 112.575 ;
        RECT 16.295 111.775 16.465 113.895 ;
        RECT 16.635 113.775 16.965 114.155 ;
        RECT 17.135 113.605 17.390 113.895 ;
        RECT 16.640 113.435 17.390 113.605 ;
        RECT 16.640 112.445 16.870 113.435 ;
        RECT 17.625 113.335 17.835 114.155 ;
        RECT 18.005 113.355 18.335 113.985 ;
        RECT 17.040 112.615 17.390 113.265 ;
        RECT 18.005 112.755 18.255 113.355 ;
        RECT 18.505 113.335 18.735 114.155 ;
        RECT 18.945 113.405 20.155 114.155 ;
        RECT 20.325 113.480 20.585 113.985 ;
        RECT 20.765 113.775 21.095 114.155 ;
        RECT 21.275 113.605 21.445 113.985 ;
        RECT 18.425 112.915 18.755 113.165 ;
        RECT 18.945 112.865 19.465 113.405 ;
        RECT 16.640 112.275 17.390 112.445 ;
        RECT 16.635 111.605 16.965 112.105 ;
        RECT 17.135 111.775 17.390 112.275 ;
        RECT 17.625 111.605 17.835 112.745 ;
        RECT 18.005 111.775 18.335 112.755 ;
        RECT 18.505 111.605 18.735 112.745 ;
        RECT 19.635 112.695 20.155 113.235 ;
        RECT 18.945 111.605 20.155 112.695 ;
        RECT 20.325 112.680 20.495 113.480 ;
        RECT 20.780 113.435 21.445 113.605 ;
        RECT 21.705 113.480 21.965 113.985 ;
        RECT 22.145 113.775 22.475 114.155 ;
        RECT 22.655 113.605 22.825 113.985 ;
        RECT 20.780 113.180 20.950 113.435 ;
        RECT 20.665 112.850 20.950 113.180 ;
        RECT 21.185 112.885 21.515 113.255 ;
        RECT 20.780 112.705 20.950 112.850 ;
        RECT 20.325 111.775 20.595 112.680 ;
        RECT 20.780 112.535 21.445 112.705 ;
        RECT 20.765 111.605 21.095 112.365 ;
        RECT 21.275 111.775 21.445 112.535 ;
        RECT 21.705 112.680 21.875 113.480 ;
        RECT 22.160 113.435 22.825 113.605 ;
        RECT 22.160 113.180 22.330 113.435 ;
        RECT 23.125 113.335 23.355 114.155 ;
        RECT 23.525 113.355 23.855 113.985 ;
        RECT 22.045 112.850 22.330 113.180 ;
        RECT 22.565 112.885 22.895 113.255 ;
        RECT 23.105 112.915 23.435 113.165 ;
        RECT 22.160 112.705 22.330 112.850 ;
        RECT 23.605 112.755 23.855 113.355 ;
        RECT 24.025 113.335 24.235 114.155 ;
        RECT 24.465 113.405 25.675 114.155 ;
        RECT 25.845 113.480 26.105 113.985 ;
        RECT 26.285 113.775 26.615 114.155 ;
        RECT 26.795 113.605 26.965 113.985 ;
        RECT 24.465 112.865 24.985 113.405 ;
        RECT 21.705 111.775 21.975 112.680 ;
        RECT 22.160 112.535 22.825 112.705 ;
        RECT 22.145 111.605 22.475 112.365 ;
        RECT 22.655 111.775 22.825 112.535 ;
        RECT 23.125 111.605 23.355 112.745 ;
        RECT 23.525 111.775 23.855 112.755 ;
        RECT 24.025 111.605 24.235 112.745 ;
        RECT 25.155 112.695 25.675 113.235 ;
        RECT 24.465 111.605 25.675 112.695 ;
        RECT 25.845 112.680 26.015 113.480 ;
        RECT 26.300 113.435 26.965 113.605 ;
        RECT 26.300 113.180 26.470 113.435 ;
        RECT 27.225 113.385 30.735 114.155 ;
        RECT 31.365 113.430 31.655 114.155 ;
        RECT 31.915 113.605 32.085 113.985 ;
        RECT 32.265 113.775 32.595 114.155 ;
        RECT 31.915 113.435 32.580 113.605 ;
        RECT 32.775 113.480 33.035 113.985 ;
        RECT 26.185 112.850 26.470 113.180 ;
        RECT 26.705 112.885 27.035 113.255 ;
        RECT 27.225 112.865 28.875 113.385 ;
        RECT 26.300 112.705 26.470 112.850 ;
        RECT 25.845 111.775 26.115 112.680 ;
        RECT 26.300 112.535 26.965 112.705 ;
        RECT 29.045 112.695 30.735 113.215 ;
        RECT 31.845 112.885 32.175 113.255 ;
        RECT 32.410 113.180 32.580 113.435 ;
        RECT 32.410 112.850 32.695 113.180 ;
        RECT 26.285 111.605 26.615 112.365 ;
        RECT 26.795 111.775 26.965 112.535 ;
        RECT 27.225 111.605 30.735 112.695 ;
        RECT 31.365 111.605 31.655 112.770 ;
        RECT 32.410 112.705 32.580 112.850 ;
        RECT 31.915 112.535 32.580 112.705 ;
        RECT 32.865 112.680 33.035 113.480 ;
        RECT 33.205 113.385 36.715 114.155 ;
        RECT 36.885 113.405 38.095 114.155 ;
        RECT 38.265 113.480 38.525 113.985 ;
        RECT 38.705 113.775 39.035 114.155 ;
        RECT 39.215 113.605 39.385 113.985 ;
        RECT 33.205 112.865 34.855 113.385 ;
        RECT 35.025 112.695 36.715 113.215 ;
        RECT 36.885 112.865 37.405 113.405 ;
        RECT 37.575 112.695 38.095 113.235 ;
        RECT 31.915 111.775 32.085 112.535 ;
        RECT 32.265 111.605 32.595 112.365 ;
        RECT 32.765 111.775 33.035 112.680 ;
        RECT 33.205 111.605 36.715 112.695 ;
        RECT 36.885 111.605 38.095 112.695 ;
        RECT 38.265 112.680 38.435 113.480 ;
        RECT 38.720 113.435 39.385 113.605 ;
        RECT 38.720 113.180 38.890 113.435 ;
        RECT 39.705 113.335 39.915 114.155 ;
        RECT 40.085 113.355 40.415 113.985 ;
        RECT 38.605 112.850 38.890 113.180 ;
        RECT 39.125 112.885 39.455 113.255 ;
        RECT 38.720 112.705 38.890 112.850 ;
        RECT 40.085 112.755 40.335 113.355 ;
        RECT 40.585 113.335 40.815 114.155 ;
        RECT 41.025 113.385 44.535 114.155 ;
        RECT 40.505 112.915 40.835 113.165 ;
        RECT 41.025 112.865 42.675 113.385 ;
        RECT 44.765 113.335 44.975 114.155 ;
        RECT 45.145 113.355 45.475 113.985 ;
        RECT 38.265 111.775 38.535 112.680 ;
        RECT 38.720 112.535 39.385 112.705 ;
        RECT 38.705 111.605 39.035 112.365 ;
        RECT 39.215 111.775 39.385 112.535 ;
        RECT 39.705 111.605 39.915 112.745 ;
        RECT 40.085 111.775 40.415 112.755 ;
        RECT 40.585 111.605 40.815 112.745 ;
        RECT 42.845 112.695 44.535 113.215 ;
        RECT 45.145 112.755 45.395 113.355 ;
        RECT 45.645 113.335 45.875 114.155 ;
        RECT 46.085 113.385 48.675 114.155 ;
        RECT 49.305 113.480 49.565 113.985 ;
        RECT 49.745 113.775 50.075 114.155 ;
        RECT 50.255 113.605 50.425 113.985 ;
        RECT 45.565 112.915 45.895 113.165 ;
        RECT 46.085 112.865 47.295 113.385 ;
        RECT 41.025 111.605 44.535 112.695 ;
        RECT 44.765 111.605 44.975 112.745 ;
        RECT 45.145 111.775 45.475 112.755 ;
        RECT 45.645 111.605 45.875 112.745 ;
        RECT 47.465 112.695 48.675 113.215 ;
        RECT 46.085 111.605 48.675 112.695 ;
        RECT 49.305 112.680 49.475 113.480 ;
        RECT 49.760 113.435 50.425 113.605 ;
        RECT 49.760 113.180 49.930 113.435 ;
        RECT 50.835 113.355 51.165 114.155 ;
        RECT 51.335 113.505 51.505 113.985 ;
        RECT 51.675 113.675 52.005 114.155 ;
        RECT 52.175 113.505 52.345 113.985 ;
        RECT 52.595 113.675 52.835 114.155 ;
        RECT 53.015 113.505 53.185 113.985 ;
        RECT 51.335 113.335 52.345 113.505 ;
        RECT 52.550 113.335 53.185 113.505 ;
        RECT 54.405 113.335 54.635 114.155 ;
        RECT 54.805 113.355 55.135 113.985 ;
        RECT 49.645 112.850 49.930 113.180 ;
        RECT 50.165 112.885 50.495 113.255 ;
        RECT 49.760 112.705 49.930 112.850 ;
        RECT 51.335 112.795 51.830 113.335 ;
        RECT 52.550 113.165 52.720 113.335 ;
        RECT 52.220 112.995 52.720 113.165 ;
        RECT 49.305 111.775 49.575 112.680 ;
        RECT 49.760 112.535 50.425 112.705 ;
        RECT 49.745 111.605 50.075 112.365 ;
        RECT 50.255 111.775 50.425 112.535 ;
        RECT 50.835 111.605 51.165 112.755 ;
        RECT 51.335 112.625 52.345 112.795 ;
        RECT 51.335 111.775 51.505 112.625 ;
        RECT 51.675 111.605 52.005 112.405 ;
        RECT 52.175 111.775 52.345 112.625 ;
        RECT 52.550 112.755 52.720 112.995 ;
        RECT 52.890 112.925 53.270 113.165 ;
        RECT 54.385 112.915 54.715 113.165 ;
        RECT 54.885 112.755 55.135 113.355 ;
        RECT 55.305 113.335 55.515 114.155 ;
        RECT 55.785 113.335 56.015 114.155 ;
        RECT 56.185 113.355 56.515 113.985 ;
        RECT 55.765 112.915 56.095 113.165 ;
        RECT 56.265 112.755 56.515 113.355 ;
        RECT 56.685 113.335 56.895 114.155 ;
        RECT 57.125 113.430 57.415 114.155 ;
        RECT 57.585 113.610 62.930 114.155 ;
        RECT 59.170 112.780 59.510 113.610 ;
        RECT 63.565 113.480 63.825 113.985 ;
        RECT 64.005 113.775 64.335 114.155 ;
        RECT 64.515 113.605 64.685 113.985 ;
        RECT 52.550 112.585 53.265 112.755 ;
        RECT 52.525 111.605 52.765 112.405 ;
        RECT 52.935 111.775 53.265 112.585 ;
        RECT 54.405 111.605 54.635 112.745 ;
        RECT 54.805 111.775 55.135 112.755 ;
        RECT 55.305 111.605 55.515 112.745 ;
        RECT 55.785 111.605 56.015 112.745 ;
        RECT 56.185 111.775 56.515 112.755 ;
        RECT 56.685 111.605 56.895 112.745 ;
        RECT 57.125 111.605 57.415 112.770 ;
        RECT 60.990 112.040 61.340 113.290 ;
        RECT 63.565 112.680 63.735 113.480 ;
        RECT 64.020 113.435 64.685 113.605 ;
        RECT 64.020 113.180 64.190 113.435 ;
        RECT 64.945 113.385 66.615 114.155 ;
        RECT 63.905 112.850 64.190 113.180 ;
        RECT 64.425 112.885 64.755 113.255 ;
        RECT 64.945 112.865 65.695 113.385 ;
        RECT 67.305 113.335 67.515 114.155 ;
        RECT 67.685 113.355 68.015 113.985 ;
        RECT 64.020 112.705 64.190 112.850 ;
        RECT 57.585 111.605 62.930 112.040 ;
        RECT 63.565 111.775 63.835 112.680 ;
        RECT 64.020 112.535 64.685 112.705 ;
        RECT 65.865 112.695 66.615 113.215 ;
        RECT 67.685 112.755 67.935 113.355 ;
        RECT 68.185 113.335 68.415 114.155 ;
        RECT 68.625 113.385 70.295 114.155 ;
        RECT 68.105 112.915 68.435 113.165 ;
        RECT 68.625 112.865 69.375 113.385 ;
        RECT 71.075 113.355 71.405 114.155 ;
        RECT 71.575 113.505 71.745 113.985 ;
        RECT 71.915 113.675 72.245 114.155 ;
        RECT 72.415 113.505 72.585 113.985 ;
        RECT 72.835 113.675 73.075 114.155 ;
        RECT 73.255 113.505 73.425 113.985 ;
        RECT 71.575 113.335 72.585 113.505 ;
        RECT 72.790 113.335 73.425 113.505 ;
        RECT 73.685 113.405 74.895 114.155 ;
        RECT 75.065 113.480 75.325 113.985 ;
        RECT 75.505 113.775 75.835 114.155 ;
        RECT 76.015 113.605 76.185 113.985 ;
        RECT 64.005 111.605 64.335 112.365 ;
        RECT 64.515 111.775 64.685 112.535 ;
        RECT 64.945 111.605 66.615 112.695 ;
        RECT 67.305 111.605 67.515 112.745 ;
        RECT 67.685 111.775 68.015 112.755 ;
        RECT 68.185 111.605 68.415 112.745 ;
        RECT 69.545 112.695 70.295 113.215 ;
        RECT 71.575 113.135 72.070 113.335 ;
        RECT 72.790 113.165 72.960 113.335 ;
        RECT 71.575 112.965 72.075 113.135 ;
        RECT 72.460 112.995 72.960 113.165 ;
        RECT 71.575 112.795 72.070 112.965 ;
        RECT 68.625 111.605 70.295 112.695 ;
        RECT 71.075 111.605 71.405 112.755 ;
        RECT 71.575 112.625 72.585 112.795 ;
        RECT 71.575 111.775 71.745 112.625 ;
        RECT 71.915 111.605 72.245 112.405 ;
        RECT 72.415 111.775 72.585 112.625 ;
        RECT 72.790 112.755 72.960 112.995 ;
        RECT 73.130 112.925 73.510 113.165 ;
        RECT 73.685 112.865 74.205 113.405 ;
        RECT 72.790 112.585 73.505 112.755 ;
        RECT 74.375 112.695 74.895 113.235 ;
        RECT 72.765 111.605 73.005 112.405 ;
        RECT 73.175 111.775 73.505 112.585 ;
        RECT 73.685 111.605 74.895 112.695 ;
        RECT 75.065 112.680 75.235 113.480 ;
        RECT 75.520 113.435 76.185 113.605 ;
        RECT 75.520 113.180 75.690 113.435 ;
        RECT 76.445 113.385 79.955 114.155 ;
        RECT 81.045 113.480 81.305 113.985 ;
        RECT 81.485 113.775 81.815 114.155 ;
        RECT 81.995 113.605 82.165 113.985 ;
        RECT 75.405 112.850 75.690 113.180 ;
        RECT 75.925 112.885 76.255 113.255 ;
        RECT 76.445 112.865 78.095 113.385 ;
        RECT 75.520 112.705 75.690 112.850 ;
        RECT 75.065 111.775 75.335 112.680 ;
        RECT 75.520 112.535 76.185 112.705 ;
        RECT 78.265 112.695 79.955 113.215 ;
        RECT 75.505 111.605 75.835 112.365 ;
        RECT 76.015 111.775 76.185 112.535 ;
        RECT 76.445 111.605 79.955 112.695 ;
        RECT 81.045 112.680 81.215 113.480 ;
        RECT 81.500 113.435 82.165 113.605 ;
        RECT 81.500 113.180 81.670 113.435 ;
        RECT 82.885 113.430 83.175 114.155 ;
        RECT 83.345 113.610 88.690 114.155 ;
        RECT 88.865 113.610 94.210 114.155 ;
        RECT 81.385 112.850 81.670 113.180 ;
        RECT 81.905 112.885 82.235 113.255 ;
        RECT 81.500 112.705 81.670 112.850 ;
        RECT 84.930 112.780 85.270 113.610 ;
        RECT 81.045 111.775 81.315 112.680 ;
        RECT 81.500 112.535 82.165 112.705 ;
        RECT 81.485 111.605 81.815 112.365 ;
        RECT 81.995 111.775 82.165 112.535 ;
        RECT 82.885 111.605 83.175 112.770 ;
        RECT 86.750 112.040 87.100 113.290 ;
        RECT 90.450 112.780 90.790 113.610 ;
        RECT 94.385 113.385 96.975 114.155 ;
        RECT 97.695 113.605 97.865 113.985 ;
        RECT 98.045 113.775 98.375 114.155 ;
        RECT 97.695 113.435 98.360 113.605 ;
        RECT 98.555 113.480 98.815 113.985 ;
        RECT 92.270 112.040 92.620 113.290 ;
        RECT 94.385 112.865 95.595 113.385 ;
        RECT 95.765 112.695 96.975 113.215 ;
        RECT 97.625 112.885 97.955 113.255 ;
        RECT 98.190 113.180 98.360 113.435 ;
        RECT 98.190 112.850 98.475 113.180 ;
        RECT 98.190 112.705 98.360 112.850 ;
        RECT 83.345 111.605 88.690 112.040 ;
        RECT 88.865 111.605 94.210 112.040 ;
        RECT 94.385 111.605 96.975 112.695 ;
        RECT 97.695 112.535 98.360 112.705 ;
        RECT 98.645 112.680 98.815 113.480 ;
        RECT 99.995 113.605 100.165 113.985 ;
        RECT 100.345 113.775 100.675 114.155 ;
        RECT 99.995 113.435 100.660 113.605 ;
        RECT 100.855 113.480 101.115 113.985 ;
        RECT 99.925 112.885 100.255 113.255 ;
        RECT 100.490 113.180 100.660 113.435 ;
        RECT 100.490 112.850 100.775 113.180 ;
        RECT 100.490 112.705 100.660 112.850 ;
        RECT 97.695 111.775 97.865 112.535 ;
        RECT 98.045 111.605 98.375 112.365 ;
        RECT 98.545 111.775 98.815 112.680 ;
        RECT 99.995 112.535 100.660 112.705 ;
        RECT 100.945 112.680 101.115 113.480 ;
        RECT 101.325 113.335 101.555 114.155 ;
        RECT 101.725 113.355 102.055 113.985 ;
        RECT 101.305 112.915 101.635 113.165 ;
        RECT 101.805 112.755 102.055 113.355 ;
        RECT 102.225 113.335 102.435 114.155 ;
        RECT 102.665 113.385 104.335 114.155 ;
        RECT 104.595 113.605 104.765 113.985 ;
        RECT 104.945 113.775 105.275 114.155 ;
        RECT 104.595 113.435 105.260 113.605 ;
        RECT 105.455 113.480 105.715 113.985 ;
        RECT 102.665 112.865 103.415 113.385 ;
        RECT 99.995 111.775 100.165 112.535 ;
        RECT 100.345 111.605 100.675 112.365 ;
        RECT 100.845 111.775 101.115 112.680 ;
        RECT 101.325 111.605 101.555 112.745 ;
        RECT 101.725 111.775 102.055 112.755 ;
        RECT 102.225 111.605 102.435 112.745 ;
        RECT 103.585 112.695 104.335 113.215 ;
        RECT 104.525 112.885 104.855 113.255 ;
        RECT 105.090 113.180 105.260 113.435 ;
        RECT 105.090 112.850 105.375 113.180 ;
        RECT 105.090 112.705 105.260 112.850 ;
        RECT 102.665 111.605 104.335 112.695 ;
        RECT 104.595 112.535 105.260 112.705 ;
        RECT 105.545 112.680 105.715 113.480 ;
        RECT 105.885 113.385 108.475 114.155 ;
        RECT 108.645 113.430 108.935 114.155 ;
        RECT 105.885 112.865 107.095 113.385 ;
        RECT 109.145 113.335 109.375 114.155 ;
        RECT 109.545 113.355 109.875 113.985 ;
        RECT 107.265 112.695 108.475 113.215 ;
        RECT 109.125 112.915 109.455 113.165 ;
        RECT 104.595 111.775 104.765 112.535 ;
        RECT 104.945 111.605 105.275 112.365 ;
        RECT 105.445 111.775 105.715 112.680 ;
        RECT 105.885 111.605 108.475 112.695 ;
        RECT 108.645 111.605 108.935 112.770 ;
        RECT 109.625 112.755 109.875 113.355 ;
        RECT 110.045 113.335 110.255 114.155 ;
        RECT 111.445 113.335 111.675 114.155 ;
        RECT 111.845 113.355 112.175 113.985 ;
        RECT 111.425 112.915 111.755 113.165 ;
        RECT 111.925 112.755 112.175 113.355 ;
        RECT 112.345 113.335 112.555 114.155 ;
        RECT 112.785 113.385 116.295 114.155 ;
        RECT 117.385 113.405 118.595 114.155 ;
        RECT 112.785 112.865 114.435 113.385 ;
        RECT 109.145 111.605 109.375 112.745 ;
        RECT 109.545 111.775 109.875 112.755 ;
        RECT 110.045 111.605 110.255 112.745 ;
        RECT 111.445 111.605 111.675 112.745 ;
        RECT 111.845 111.775 112.175 112.755 ;
        RECT 112.345 111.605 112.555 112.745 ;
        RECT 114.605 112.695 116.295 113.215 ;
        RECT 112.785 111.605 116.295 112.695 ;
        RECT 117.385 112.695 117.905 113.235 ;
        RECT 118.075 112.865 118.595 113.405 ;
        RECT 117.385 111.605 118.595 112.695 ;
        RECT 5.520 111.435 118.680 111.605 ;
        RECT 5.605 110.345 6.815 111.435 ;
        RECT 6.985 110.345 9.575 111.435 ;
        RECT 5.605 109.635 6.125 110.175 ;
        RECT 6.295 109.805 6.815 110.345 ;
        RECT 6.985 109.655 8.195 110.175 ;
        RECT 8.365 109.825 9.575 110.345 ;
        RECT 9.835 110.505 10.005 111.265 ;
        RECT 10.185 110.675 10.515 111.435 ;
        RECT 9.835 110.335 10.500 110.505 ;
        RECT 10.685 110.360 10.955 111.265 ;
        RECT 10.330 110.190 10.500 110.335 ;
        RECT 9.765 109.785 10.095 110.155 ;
        RECT 10.330 109.860 10.615 110.190 ;
        RECT 5.605 108.885 6.815 109.635 ;
        RECT 6.985 108.885 9.575 109.655 ;
        RECT 10.330 109.605 10.500 109.860 ;
        RECT 9.835 109.435 10.500 109.605 ;
        RECT 10.785 109.560 10.955 110.360 ;
        RECT 11.215 110.505 11.385 111.265 ;
        RECT 11.565 110.675 11.895 111.435 ;
        RECT 11.215 110.335 11.880 110.505 ;
        RECT 12.065 110.360 12.335 111.265 ;
        RECT 11.710 110.190 11.880 110.335 ;
        RECT 11.145 109.785 11.475 110.155 ;
        RECT 11.710 109.860 11.995 110.190 ;
        RECT 11.710 109.605 11.880 109.860 ;
        RECT 9.835 109.055 10.005 109.435 ;
        RECT 10.185 108.885 10.515 109.265 ;
        RECT 10.695 109.055 10.955 109.560 ;
        RECT 11.215 109.435 11.880 109.605 ;
        RECT 12.165 109.560 12.335 110.360 ;
        RECT 12.565 110.295 12.775 111.435 ;
        RECT 12.945 110.285 13.275 111.265 ;
        RECT 13.445 110.295 13.675 111.435 ;
        RECT 13.885 110.345 17.395 111.435 ;
        RECT 11.215 109.055 11.385 109.435 ;
        RECT 11.565 108.885 11.895 109.265 ;
        RECT 12.075 109.055 12.335 109.560 ;
        RECT 12.565 108.885 12.775 109.705 ;
        RECT 12.945 109.685 13.195 110.285 ;
        RECT 13.365 109.875 13.695 110.125 ;
        RECT 12.945 109.055 13.275 109.685 ;
        RECT 13.445 108.885 13.675 109.705 ;
        RECT 13.885 109.655 15.535 110.175 ;
        RECT 15.705 109.825 17.395 110.345 ;
        RECT 18.485 110.270 18.775 111.435 ;
        RECT 18.945 111.000 24.290 111.435 ;
        RECT 24.465 111.000 29.810 111.435 ;
        RECT 13.885 108.885 17.395 109.655 ;
        RECT 18.485 108.885 18.775 109.610 ;
        RECT 20.530 109.430 20.870 110.260 ;
        RECT 22.350 109.750 22.700 111.000 ;
        RECT 26.050 109.430 26.390 110.260 ;
        RECT 27.870 109.750 28.220 111.000 ;
        RECT 29.985 110.465 30.245 111.435 ;
        RECT 18.945 108.885 24.290 109.430 ;
        RECT 24.465 108.885 29.810 109.430 ;
        RECT 29.985 109.175 30.225 110.125 ;
        RECT 30.415 110.090 30.745 111.265 ;
        RECT 30.915 110.465 31.195 111.435 ;
        RECT 31.455 110.690 31.725 111.435 ;
        RECT 32.355 111.430 38.630 111.435 ;
        RECT 31.895 110.520 32.185 111.260 ;
        RECT 32.355 110.705 32.610 111.430 ;
        RECT 32.795 110.535 33.055 111.260 ;
        RECT 33.225 110.705 33.470 111.430 ;
        RECT 33.655 110.535 33.915 111.260 ;
        RECT 34.085 110.705 34.330 111.430 ;
        RECT 34.515 110.535 34.775 111.260 ;
        RECT 34.945 110.705 35.190 111.430 ;
        RECT 35.360 110.535 35.620 111.260 ;
        RECT 35.790 110.705 36.050 111.430 ;
        RECT 36.220 110.535 36.480 111.260 ;
        RECT 36.650 110.705 36.910 111.430 ;
        RECT 37.080 110.535 37.340 111.260 ;
        RECT 37.510 110.705 37.770 111.430 ;
        RECT 37.940 110.535 38.200 111.260 ;
        RECT 38.370 110.635 38.630 111.430 ;
        RECT 32.795 110.520 38.200 110.535 ;
        RECT 31.455 110.295 38.200 110.520 ;
        RECT 30.415 109.560 31.195 110.090 ;
        RECT 31.455 109.735 32.620 110.295 ;
        RECT 38.800 110.125 39.050 111.260 ;
        RECT 39.230 110.625 39.490 111.435 ;
        RECT 39.665 110.125 39.910 111.265 ;
        RECT 40.090 110.625 40.385 111.435 ;
        RECT 40.565 110.345 44.075 111.435 ;
        RECT 32.790 109.875 39.910 110.125 ;
        RECT 31.425 109.705 32.620 109.735 ;
        RECT 31.425 109.565 38.200 109.705 ;
        RECT 30.415 109.055 30.740 109.560 ;
        RECT 31.455 109.535 38.200 109.565 ;
        RECT 30.910 108.885 31.195 109.390 ;
        RECT 31.455 108.885 31.755 109.365 ;
        RECT 31.925 109.080 32.185 109.535 ;
        RECT 32.355 108.885 32.615 109.365 ;
        RECT 32.795 109.080 33.055 109.535 ;
        RECT 33.225 108.885 33.475 109.365 ;
        RECT 33.655 109.080 33.915 109.535 ;
        RECT 34.085 108.885 34.335 109.365 ;
        RECT 34.515 109.080 34.775 109.535 ;
        RECT 34.945 108.885 35.190 109.365 ;
        RECT 35.360 109.080 35.635 109.535 ;
        RECT 35.805 108.885 36.050 109.365 ;
        RECT 36.220 109.080 36.480 109.535 ;
        RECT 36.650 108.885 36.910 109.365 ;
        RECT 37.080 109.080 37.340 109.535 ;
        RECT 37.510 108.885 37.770 109.365 ;
        RECT 37.940 109.080 38.200 109.535 ;
        RECT 38.370 108.885 38.630 109.445 ;
        RECT 38.800 109.065 39.050 109.875 ;
        RECT 39.230 108.885 39.490 109.410 ;
        RECT 39.660 109.065 39.910 109.875 ;
        RECT 40.080 109.565 40.395 110.125 ;
        RECT 40.565 109.655 42.215 110.175 ;
        RECT 42.385 109.825 44.075 110.345 ;
        RECT 44.245 110.270 44.535 111.435 ;
        RECT 44.705 111.000 50.050 111.435 ;
        RECT 40.090 108.885 40.395 109.395 ;
        RECT 40.565 108.885 44.075 109.655 ;
        RECT 44.245 108.885 44.535 109.610 ;
        RECT 46.290 109.430 46.630 110.260 ;
        RECT 48.110 109.750 48.460 111.000 ;
        RECT 50.225 110.345 51.435 111.435 ;
        RECT 50.225 109.635 50.745 110.175 ;
        RECT 50.915 109.805 51.435 110.345 ;
        RECT 51.645 110.295 51.875 111.435 ;
        RECT 52.045 110.285 52.375 111.265 ;
        RECT 52.545 110.295 52.755 111.435 ;
        RECT 52.985 111.000 58.330 111.435 ;
        RECT 58.505 111.000 63.850 111.435 ;
        RECT 64.025 111.000 69.370 111.435 ;
        RECT 51.625 109.875 51.955 110.125 ;
        RECT 44.705 108.885 50.050 109.430 ;
        RECT 50.225 108.885 51.435 109.635 ;
        RECT 51.645 108.885 51.875 109.705 ;
        RECT 52.125 109.685 52.375 110.285 ;
        RECT 52.045 109.055 52.375 109.685 ;
        RECT 52.545 108.885 52.755 109.705 ;
        RECT 54.570 109.430 54.910 110.260 ;
        RECT 56.390 109.750 56.740 111.000 ;
        RECT 60.090 109.430 60.430 110.260 ;
        RECT 61.910 109.750 62.260 111.000 ;
        RECT 65.610 109.430 65.950 110.260 ;
        RECT 67.430 109.750 67.780 111.000 ;
        RECT 70.005 110.270 70.295 111.435 ;
        RECT 70.465 111.000 75.810 111.435 ;
        RECT 75.985 111.000 81.330 111.435 ;
        RECT 52.985 108.885 58.330 109.430 ;
        RECT 58.505 108.885 63.850 109.430 ;
        RECT 64.025 108.885 69.370 109.430 ;
        RECT 70.005 108.885 70.295 109.610 ;
        RECT 72.050 109.430 72.390 110.260 ;
        RECT 73.870 109.750 74.220 111.000 ;
        RECT 77.570 109.430 77.910 110.260 ;
        RECT 79.390 109.750 79.740 111.000 ;
        RECT 81.505 110.345 85.015 111.435 ;
        RECT 86.115 110.625 86.410 111.435 ;
        RECT 81.505 109.655 83.155 110.175 ;
        RECT 83.325 109.825 85.015 110.345 ;
        RECT 86.590 110.125 86.835 111.265 ;
        RECT 87.010 110.625 87.270 111.435 ;
        RECT 87.870 111.430 94.145 111.435 ;
        RECT 87.450 110.125 87.700 111.260 ;
        RECT 87.870 110.635 88.130 111.430 ;
        RECT 88.300 110.535 88.560 111.260 ;
        RECT 88.730 110.705 88.990 111.430 ;
        RECT 89.160 110.535 89.420 111.260 ;
        RECT 89.590 110.705 89.850 111.430 ;
        RECT 90.020 110.535 90.280 111.260 ;
        RECT 90.450 110.705 90.710 111.430 ;
        RECT 90.880 110.535 91.140 111.260 ;
        RECT 91.310 110.705 91.555 111.430 ;
        RECT 91.725 110.535 91.985 111.260 ;
        RECT 92.170 110.705 92.415 111.430 ;
        RECT 92.585 110.535 92.845 111.260 ;
        RECT 93.030 110.705 93.275 111.430 ;
        RECT 93.445 110.535 93.705 111.260 ;
        RECT 93.890 110.705 94.145 111.430 ;
        RECT 88.300 110.520 93.705 110.535 ;
        RECT 94.315 110.520 94.605 111.260 ;
        RECT 94.775 110.690 95.045 111.435 ;
        RECT 88.300 110.295 95.045 110.520 ;
        RECT 70.465 108.885 75.810 109.430 ;
        RECT 75.985 108.885 81.330 109.430 ;
        RECT 81.505 108.885 85.015 109.655 ;
        RECT 86.105 109.565 86.420 110.125 ;
        RECT 86.590 109.875 93.710 110.125 ;
        RECT 86.105 108.885 86.410 109.395 ;
        RECT 86.590 109.065 86.840 109.875 ;
        RECT 87.010 108.885 87.270 109.410 ;
        RECT 87.450 109.065 87.700 109.875 ;
        RECT 93.880 109.705 95.045 110.295 ;
        RECT 95.765 110.270 96.055 111.435 ;
        RECT 96.225 110.345 97.895 111.435 ;
        RECT 88.300 109.535 95.045 109.705 ;
        RECT 96.225 109.655 96.975 110.175 ;
        RECT 97.145 109.825 97.895 110.345 ;
        RECT 98.105 110.295 98.335 111.435 ;
        RECT 98.505 110.285 98.835 111.265 ;
        RECT 99.005 110.295 99.215 111.435 ;
        RECT 99.445 111.000 104.790 111.435 ;
        RECT 98.085 109.875 98.415 110.125 ;
        RECT 87.870 108.885 88.130 109.445 ;
        RECT 88.300 109.080 88.560 109.535 ;
        RECT 88.730 108.885 88.990 109.365 ;
        RECT 89.160 109.080 89.420 109.535 ;
        RECT 89.590 108.885 89.850 109.365 ;
        RECT 90.020 109.080 90.280 109.535 ;
        RECT 90.450 108.885 90.695 109.365 ;
        RECT 90.865 109.080 91.140 109.535 ;
        RECT 91.310 108.885 91.555 109.365 ;
        RECT 91.725 109.080 91.985 109.535 ;
        RECT 92.165 108.885 92.415 109.365 ;
        RECT 92.585 109.080 92.845 109.535 ;
        RECT 93.025 108.885 93.275 109.365 ;
        RECT 93.445 109.080 93.705 109.535 ;
        RECT 93.885 108.885 94.145 109.365 ;
        RECT 94.315 109.080 94.575 109.535 ;
        RECT 94.745 108.885 95.045 109.365 ;
        RECT 95.765 108.885 96.055 109.610 ;
        RECT 96.225 108.885 97.895 109.655 ;
        RECT 98.105 108.885 98.335 109.705 ;
        RECT 98.585 109.685 98.835 110.285 ;
        RECT 98.505 109.055 98.835 109.685 ;
        RECT 99.005 108.885 99.215 109.705 ;
        RECT 101.030 109.430 101.370 110.260 ;
        RECT 102.850 109.750 103.200 111.000 ;
        RECT 104.965 110.345 106.635 111.435 ;
        RECT 106.810 110.765 107.065 111.265 ;
        RECT 107.235 110.935 107.565 111.435 ;
        RECT 106.810 110.595 107.560 110.765 ;
        RECT 104.965 109.655 105.715 110.175 ;
        RECT 105.885 109.825 106.635 110.345 ;
        RECT 106.810 109.775 107.160 110.425 ;
        RECT 99.445 108.885 104.790 109.430 ;
        RECT 104.965 108.885 106.635 109.655 ;
        RECT 107.330 109.605 107.560 110.595 ;
        RECT 106.810 109.435 107.560 109.605 ;
        RECT 106.810 109.145 107.065 109.435 ;
        RECT 107.235 108.885 107.565 109.265 ;
        RECT 107.735 109.145 107.905 111.265 ;
        RECT 108.075 110.465 108.400 111.250 ;
        RECT 108.570 110.975 108.820 111.435 ;
        RECT 108.990 110.935 109.240 111.265 ;
        RECT 109.455 110.935 110.135 111.265 ;
        RECT 108.990 110.805 109.160 110.935 ;
        RECT 108.765 110.635 109.160 110.805 ;
        RECT 108.135 109.415 108.595 110.465 ;
        RECT 108.765 109.275 108.935 110.635 ;
        RECT 109.330 110.375 109.795 110.765 ;
        RECT 109.105 109.565 109.455 110.185 ;
        RECT 109.625 109.785 109.795 110.375 ;
        RECT 109.965 110.155 110.135 110.935 ;
        RECT 110.305 110.835 110.475 111.175 ;
        RECT 110.710 111.005 111.040 111.435 ;
        RECT 111.210 110.835 111.380 111.175 ;
        RECT 111.675 110.975 112.045 111.435 ;
        RECT 110.305 110.665 111.380 110.835 ;
        RECT 112.215 110.805 112.385 111.265 ;
        RECT 112.620 110.925 113.490 111.265 ;
        RECT 113.660 110.975 113.910 111.435 ;
        RECT 111.825 110.635 112.385 110.805 ;
        RECT 111.825 110.495 111.995 110.635 ;
        RECT 110.495 110.325 111.995 110.495 ;
        RECT 112.690 110.465 113.150 110.755 ;
        RECT 109.965 109.985 111.655 110.155 ;
        RECT 109.625 109.565 109.980 109.785 ;
        RECT 110.150 109.275 110.320 109.985 ;
        RECT 110.525 109.565 111.315 109.815 ;
        RECT 111.485 109.805 111.655 109.985 ;
        RECT 111.825 109.635 111.995 110.325 ;
        RECT 108.265 108.885 108.595 109.245 ;
        RECT 108.765 109.105 109.260 109.275 ;
        RECT 109.465 109.105 110.320 109.275 ;
        RECT 111.195 108.885 111.525 109.345 ;
        RECT 111.735 109.245 111.995 109.635 ;
        RECT 112.185 110.455 113.150 110.465 ;
        RECT 113.320 110.545 113.490 110.925 ;
        RECT 114.080 110.885 114.250 111.175 ;
        RECT 114.430 111.055 114.760 111.435 ;
        RECT 114.080 110.715 114.880 110.885 ;
        RECT 112.185 110.295 112.860 110.455 ;
        RECT 113.320 110.375 114.540 110.545 ;
        RECT 112.185 109.505 112.395 110.295 ;
        RECT 113.320 110.285 113.490 110.375 ;
        RECT 112.565 109.505 112.915 110.125 ;
        RECT 113.085 110.115 113.490 110.285 ;
        RECT 113.085 109.335 113.255 110.115 ;
        RECT 113.425 109.665 113.645 109.945 ;
        RECT 113.825 109.835 114.365 110.205 ;
        RECT 114.710 110.095 114.880 110.715 ;
        RECT 115.055 110.375 115.225 111.435 ;
        RECT 115.435 110.425 115.725 111.265 ;
        RECT 115.895 110.595 116.065 111.435 ;
        RECT 116.275 110.425 116.525 111.265 ;
        RECT 116.735 110.595 116.905 111.435 ;
        RECT 115.435 110.255 117.160 110.425 ;
        RECT 113.425 109.495 113.955 109.665 ;
        RECT 111.735 109.075 112.085 109.245 ;
        RECT 112.305 109.055 113.255 109.335 ;
        RECT 113.425 108.885 113.615 109.325 ;
        RECT 113.785 109.265 113.955 109.495 ;
        RECT 114.125 109.435 114.365 109.835 ;
        RECT 114.535 110.085 114.880 110.095 ;
        RECT 114.535 109.875 116.565 110.085 ;
        RECT 114.535 109.620 114.860 109.875 ;
        RECT 116.750 109.705 117.160 110.255 ;
        RECT 117.385 110.345 118.595 111.435 ;
        RECT 117.385 109.805 117.905 110.345 ;
        RECT 114.535 109.265 114.855 109.620 ;
        RECT 113.785 109.095 114.855 109.265 ;
        RECT 115.055 108.885 115.225 109.695 ;
        RECT 115.395 109.535 117.160 109.705 ;
        RECT 118.075 109.635 118.595 110.175 ;
        RECT 115.395 109.055 115.725 109.535 ;
        RECT 115.895 108.885 116.065 109.355 ;
        RECT 116.235 109.055 116.565 109.535 ;
        RECT 116.735 108.885 116.905 109.355 ;
        RECT 117.385 108.885 118.595 109.635 ;
        RECT 5.520 108.715 118.680 108.885 ;
        RECT 5.605 107.965 6.815 108.715 ;
        RECT 6.985 108.170 12.330 108.715 ;
        RECT 12.505 108.170 17.850 108.715 ;
        RECT 5.605 107.425 6.125 107.965 ;
        RECT 6.295 107.255 6.815 107.795 ;
        RECT 8.570 107.340 8.910 108.170 ;
        RECT 5.605 106.165 6.815 107.255 ;
        RECT 10.390 106.600 10.740 107.850 ;
        RECT 14.090 107.340 14.430 108.170 ;
        RECT 18.030 107.975 18.285 108.545 ;
        RECT 18.455 108.315 18.785 108.715 ;
        RECT 19.210 108.180 19.740 108.545 ;
        RECT 19.210 108.145 19.385 108.180 ;
        RECT 18.455 107.975 19.385 108.145 ;
        RECT 15.910 106.600 16.260 107.850 ;
        RECT 18.030 107.305 18.200 107.975 ;
        RECT 18.455 107.805 18.625 107.975 ;
        RECT 18.370 107.475 18.625 107.805 ;
        RECT 18.850 107.475 19.045 107.805 ;
        RECT 6.985 106.165 12.330 106.600 ;
        RECT 12.505 106.165 17.850 106.600 ;
        RECT 18.030 106.335 18.365 107.305 ;
        RECT 18.535 106.165 18.705 107.305 ;
        RECT 18.875 106.505 19.045 107.475 ;
        RECT 19.215 106.845 19.385 107.975 ;
        RECT 19.555 107.185 19.725 107.985 ;
        RECT 19.930 107.695 20.205 108.545 ;
        RECT 19.925 107.525 20.205 107.695 ;
        RECT 19.930 107.385 20.205 107.525 ;
        RECT 20.375 107.185 20.565 108.545 ;
        RECT 20.745 108.180 21.255 108.715 ;
        RECT 21.475 107.905 21.720 108.510 ;
        RECT 22.165 107.945 23.835 108.715 ;
        RECT 24.005 108.040 24.265 108.545 ;
        RECT 24.445 108.335 24.775 108.715 ;
        RECT 24.955 108.165 25.125 108.545 ;
        RECT 25.385 108.170 30.730 108.715 ;
        RECT 20.765 107.735 21.995 107.905 ;
        RECT 19.555 107.015 20.565 107.185 ;
        RECT 20.735 107.170 21.485 107.360 ;
        RECT 19.215 106.675 20.340 106.845 ;
        RECT 20.735 106.505 20.905 107.170 ;
        RECT 21.655 106.925 21.995 107.735 ;
        RECT 22.165 107.425 22.915 107.945 ;
        RECT 23.085 107.255 23.835 107.775 ;
        RECT 18.875 106.335 20.905 106.505 ;
        RECT 21.075 106.165 21.245 106.925 ;
        RECT 21.480 106.515 21.995 106.925 ;
        RECT 22.165 106.165 23.835 107.255 ;
        RECT 24.005 107.240 24.175 108.040 ;
        RECT 24.460 107.995 25.125 108.165 ;
        RECT 24.460 107.740 24.630 107.995 ;
        RECT 24.345 107.410 24.630 107.740 ;
        RECT 24.865 107.445 25.195 107.815 ;
        RECT 24.460 107.265 24.630 107.410 ;
        RECT 26.970 107.340 27.310 108.170 ;
        RECT 31.365 107.990 31.655 108.715 ;
        RECT 31.915 108.165 32.085 108.545 ;
        RECT 32.265 108.335 32.595 108.715 ;
        RECT 31.915 107.995 32.580 108.165 ;
        RECT 32.775 108.040 33.035 108.545 ;
        RECT 24.005 106.335 24.275 107.240 ;
        RECT 24.460 107.095 25.125 107.265 ;
        RECT 24.445 106.165 24.775 106.925 ;
        RECT 24.955 106.335 25.125 107.095 ;
        RECT 28.790 106.600 29.140 107.850 ;
        RECT 31.845 107.445 32.175 107.815 ;
        RECT 32.410 107.740 32.580 107.995 ;
        RECT 32.410 107.410 32.695 107.740 ;
        RECT 25.385 106.165 30.730 106.600 ;
        RECT 31.365 106.165 31.655 107.330 ;
        RECT 32.410 107.265 32.580 107.410 ;
        RECT 31.915 107.095 32.580 107.265 ;
        RECT 32.865 107.240 33.035 108.040 ;
        RECT 33.205 107.945 35.795 108.715 ;
        RECT 36.800 108.005 37.055 108.535 ;
        RECT 37.235 108.255 37.520 108.715 ;
        RECT 33.205 107.425 34.415 107.945 ;
        RECT 34.585 107.255 35.795 107.775 ;
        RECT 31.915 106.335 32.085 107.095 ;
        RECT 32.265 106.165 32.595 106.925 ;
        RECT 32.765 106.335 33.035 107.240 ;
        RECT 33.205 106.165 35.795 107.255 ;
        RECT 36.800 107.145 36.980 108.005 ;
        RECT 37.700 107.805 37.950 108.455 ;
        RECT 37.150 107.475 37.950 107.805 ;
        RECT 36.800 106.675 37.055 107.145 ;
        RECT 36.715 106.505 37.055 106.675 ;
        RECT 36.800 106.475 37.055 106.505 ;
        RECT 37.235 106.165 37.520 106.965 ;
        RECT 37.700 106.885 37.950 107.475 ;
        RECT 38.150 108.120 38.470 108.450 ;
        RECT 38.650 108.235 39.310 108.715 ;
        RECT 39.510 108.325 40.360 108.495 ;
        RECT 38.150 107.225 38.340 108.120 ;
        RECT 38.660 107.795 39.320 108.065 ;
        RECT 38.990 107.735 39.320 107.795 ;
        RECT 38.510 107.565 38.840 107.625 ;
        RECT 39.510 107.565 39.680 108.325 ;
        RECT 40.920 108.255 41.240 108.715 ;
        RECT 41.440 108.075 41.690 108.505 ;
        RECT 41.980 108.275 42.390 108.715 ;
        RECT 42.560 108.335 43.575 108.535 ;
        RECT 39.850 107.905 41.100 108.075 ;
        RECT 39.850 107.785 40.180 107.905 ;
        RECT 38.510 107.395 40.410 107.565 ;
        RECT 38.150 107.055 40.070 107.225 ;
        RECT 38.150 107.035 38.470 107.055 ;
        RECT 37.700 106.375 38.030 106.885 ;
        RECT 38.300 106.425 38.470 107.035 ;
        RECT 40.240 106.885 40.410 107.395 ;
        RECT 40.580 107.325 40.760 107.735 ;
        RECT 40.930 107.145 41.100 107.905 ;
        RECT 38.640 106.165 38.970 106.855 ;
        RECT 39.200 106.715 40.410 106.885 ;
        RECT 40.580 106.835 41.100 107.145 ;
        RECT 41.270 107.735 41.690 108.075 ;
        RECT 41.980 107.735 42.390 108.065 ;
        RECT 41.270 106.965 41.460 107.735 ;
        RECT 42.560 107.605 42.730 108.335 ;
        RECT 43.875 108.165 44.045 108.495 ;
        RECT 44.215 108.335 44.545 108.715 ;
        RECT 42.900 107.785 43.250 108.155 ;
        RECT 42.560 107.565 42.980 107.605 ;
        RECT 41.630 107.395 42.980 107.565 ;
        RECT 41.630 107.235 41.880 107.395 ;
        RECT 42.390 106.965 42.640 107.225 ;
        RECT 41.270 106.715 42.640 106.965 ;
        RECT 39.200 106.425 39.440 106.715 ;
        RECT 40.240 106.635 40.410 106.715 ;
        RECT 39.640 106.165 40.060 106.545 ;
        RECT 40.240 106.385 40.870 106.635 ;
        RECT 41.340 106.165 41.670 106.545 ;
        RECT 41.840 106.425 42.010 106.715 ;
        RECT 42.810 106.550 42.980 107.395 ;
        RECT 43.430 107.225 43.650 108.095 ;
        RECT 43.875 107.975 44.570 108.165 ;
        RECT 43.150 106.845 43.650 107.225 ;
        RECT 43.820 107.175 44.230 107.795 ;
        RECT 44.400 107.005 44.570 107.975 ;
        RECT 43.875 106.835 44.570 107.005 ;
        RECT 42.190 106.165 42.570 106.545 ;
        RECT 42.810 106.380 43.640 106.550 ;
        RECT 43.875 106.335 44.045 106.835 ;
        RECT 44.215 106.165 44.545 106.665 ;
        RECT 44.760 106.335 44.985 108.455 ;
        RECT 45.155 108.335 45.485 108.715 ;
        RECT 45.655 108.165 45.825 108.455 ;
        RECT 45.160 107.995 45.825 108.165 ;
        RECT 46.635 108.165 46.805 108.455 ;
        RECT 46.975 108.335 47.305 108.715 ;
        RECT 46.635 107.995 47.300 108.165 ;
        RECT 45.160 107.005 45.390 107.995 ;
        RECT 45.560 107.175 45.910 107.825 ;
        RECT 46.550 107.175 46.900 107.825 ;
        RECT 47.070 107.005 47.300 107.995 ;
        RECT 45.160 106.835 45.825 107.005 ;
        RECT 45.155 106.165 45.485 106.665 ;
        RECT 45.655 106.335 45.825 106.835 ;
        RECT 46.635 106.835 47.300 107.005 ;
        RECT 46.635 106.335 46.805 106.835 ;
        RECT 46.975 106.165 47.305 106.665 ;
        RECT 47.475 106.335 47.700 108.455 ;
        RECT 47.915 108.335 48.245 108.715 ;
        RECT 48.415 108.165 48.585 108.495 ;
        RECT 48.885 108.335 49.900 108.535 ;
        RECT 47.890 107.975 48.585 108.165 ;
        RECT 47.890 107.005 48.060 107.975 ;
        RECT 48.230 107.175 48.640 107.795 ;
        RECT 48.810 107.225 49.030 108.095 ;
        RECT 49.210 107.785 49.560 108.155 ;
        RECT 49.730 107.605 49.900 108.335 ;
        RECT 50.070 108.275 50.480 108.715 ;
        RECT 50.770 108.075 51.020 108.505 ;
        RECT 51.220 108.255 51.540 108.715 ;
        RECT 52.100 108.325 52.950 108.495 ;
        RECT 50.070 107.735 50.480 108.065 ;
        RECT 50.770 107.735 51.190 108.075 ;
        RECT 49.480 107.565 49.900 107.605 ;
        RECT 49.480 107.395 50.830 107.565 ;
        RECT 47.890 106.835 48.585 107.005 ;
        RECT 48.810 106.845 49.310 107.225 ;
        RECT 47.915 106.165 48.245 106.665 ;
        RECT 48.415 106.335 48.585 106.835 ;
        RECT 49.480 106.550 49.650 107.395 ;
        RECT 50.580 107.235 50.830 107.395 ;
        RECT 49.820 106.965 50.070 107.225 ;
        RECT 51.000 106.965 51.190 107.735 ;
        RECT 49.820 106.715 51.190 106.965 ;
        RECT 51.360 107.905 52.610 108.075 ;
        RECT 51.360 107.145 51.530 107.905 ;
        RECT 52.280 107.785 52.610 107.905 ;
        RECT 51.700 107.325 51.880 107.735 ;
        RECT 52.780 107.565 52.950 108.325 ;
        RECT 53.150 108.235 53.810 108.715 ;
        RECT 53.990 108.120 54.310 108.450 ;
        RECT 53.140 107.795 53.800 108.065 ;
        RECT 53.140 107.735 53.470 107.795 ;
        RECT 53.620 107.565 53.950 107.625 ;
        RECT 52.050 107.395 53.950 107.565 ;
        RECT 51.360 106.835 51.880 107.145 ;
        RECT 52.050 106.885 52.220 107.395 ;
        RECT 54.120 107.225 54.310 108.120 ;
        RECT 52.390 107.055 54.310 107.225 ;
        RECT 53.990 107.035 54.310 107.055 ;
        RECT 54.510 107.805 54.760 108.455 ;
        RECT 54.940 108.255 55.225 108.715 ;
        RECT 55.405 108.005 55.660 108.535 ;
        RECT 54.510 107.475 55.310 107.805 ;
        RECT 52.050 106.715 53.260 106.885 ;
        RECT 48.820 106.380 49.650 106.550 ;
        RECT 49.890 106.165 50.270 106.545 ;
        RECT 50.450 106.425 50.620 106.715 ;
        RECT 52.050 106.635 52.220 106.715 ;
        RECT 50.790 106.165 51.120 106.545 ;
        RECT 51.590 106.385 52.220 106.635 ;
        RECT 52.400 106.165 52.820 106.545 ;
        RECT 53.020 106.425 53.260 106.715 ;
        RECT 53.490 106.165 53.820 106.855 ;
        RECT 53.990 106.425 54.160 107.035 ;
        RECT 54.510 106.885 54.760 107.475 ;
        RECT 55.480 107.145 55.660 108.005 ;
        RECT 57.125 107.990 57.415 108.715 ;
        RECT 57.585 108.170 62.930 108.715 ;
        RECT 59.170 107.340 59.510 108.170 ;
        RECT 64.025 108.040 64.285 108.545 ;
        RECT 64.465 108.335 64.795 108.715 ;
        RECT 64.975 108.165 65.145 108.545 ;
        RECT 54.430 106.375 54.760 106.885 ;
        RECT 54.940 106.165 55.225 106.965 ;
        RECT 55.405 106.675 55.660 107.145 ;
        RECT 55.405 106.505 55.745 106.675 ;
        RECT 55.405 106.475 55.660 106.505 ;
        RECT 57.125 106.165 57.415 107.330 ;
        RECT 60.990 106.600 61.340 107.850 ;
        RECT 64.025 107.240 64.195 108.040 ;
        RECT 64.480 107.995 65.145 108.165 ;
        RECT 64.480 107.740 64.650 107.995 ;
        RECT 65.925 107.895 66.135 108.715 ;
        RECT 66.305 107.915 66.635 108.545 ;
        RECT 64.365 107.410 64.650 107.740 ;
        RECT 64.885 107.445 65.215 107.815 ;
        RECT 64.480 107.265 64.650 107.410 ;
        RECT 66.305 107.315 66.555 107.915 ;
        RECT 66.805 107.895 67.035 108.715 ;
        RECT 67.245 108.170 72.590 108.715 ;
        RECT 72.765 108.170 78.110 108.715 ;
        RECT 66.725 107.475 67.055 107.725 ;
        RECT 68.830 107.340 69.170 108.170 ;
        RECT 57.585 106.165 62.930 106.600 ;
        RECT 64.025 106.335 64.295 107.240 ;
        RECT 64.480 107.095 65.145 107.265 ;
        RECT 64.465 106.165 64.795 106.925 ;
        RECT 64.975 106.335 65.145 107.095 ;
        RECT 65.925 106.165 66.135 107.305 ;
        RECT 66.305 106.335 66.635 107.315 ;
        RECT 66.805 106.165 67.035 107.305 ;
        RECT 70.650 106.600 71.000 107.850 ;
        RECT 74.350 107.340 74.690 108.170 ;
        RECT 78.285 107.965 79.495 108.715 ;
        RECT 79.665 108.040 79.925 108.545 ;
        RECT 80.105 108.335 80.435 108.715 ;
        RECT 80.615 108.165 80.785 108.545 ;
        RECT 76.170 106.600 76.520 107.850 ;
        RECT 78.285 107.425 78.805 107.965 ;
        RECT 78.975 107.255 79.495 107.795 ;
        RECT 67.245 106.165 72.590 106.600 ;
        RECT 72.765 106.165 78.110 106.600 ;
        RECT 78.285 106.165 79.495 107.255 ;
        RECT 79.665 107.240 79.835 108.040 ;
        RECT 80.120 107.995 80.785 108.165 ;
        RECT 80.120 107.740 80.290 107.995 ;
        RECT 81.045 107.945 82.715 108.715 ;
        RECT 82.885 107.990 83.175 108.715 ;
        RECT 80.005 107.410 80.290 107.740 ;
        RECT 80.525 107.445 80.855 107.815 ;
        RECT 81.045 107.425 81.795 107.945 ;
        RECT 84.080 107.905 84.325 108.510 ;
        RECT 84.545 108.180 85.055 108.715 ;
        RECT 80.120 107.265 80.290 107.410 ;
        RECT 79.665 106.335 79.935 107.240 ;
        RECT 80.120 107.095 80.785 107.265 ;
        RECT 81.965 107.255 82.715 107.775 ;
        RECT 83.805 107.735 85.035 107.905 ;
        RECT 80.105 106.165 80.435 106.925 ;
        RECT 80.615 106.335 80.785 107.095 ;
        RECT 81.045 106.165 82.715 107.255 ;
        RECT 82.885 106.165 83.175 107.330 ;
        RECT 83.805 106.925 84.145 107.735 ;
        RECT 84.315 107.170 85.065 107.360 ;
        RECT 83.805 106.515 84.320 106.925 ;
        RECT 84.555 106.165 84.725 106.925 ;
        RECT 84.895 106.505 85.065 107.170 ;
        RECT 85.235 107.185 85.425 108.545 ;
        RECT 85.595 108.035 85.870 108.545 ;
        RECT 86.060 108.180 86.590 108.545 ;
        RECT 87.015 108.315 87.345 108.715 ;
        RECT 86.415 108.145 86.590 108.180 ;
        RECT 85.595 107.865 85.875 108.035 ;
        RECT 85.595 107.385 85.870 107.865 ;
        RECT 86.075 107.185 86.245 107.985 ;
        RECT 85.235 107.015 86.245 107.185 ;
        RECT 86.415 107.975 87.345 108.145 ;
        RECT 87.515 107.975 87.770 108.545 ;
        RECT 86.415 106.845 86.585 107.975 ;
        RECT 87.175 107.805 87.345 107.975 ;
        RECT 85.460 106.675 86.585 106.845 ;
        RECT 86.755 107.475 86.950 107.805 ;
        RECT 87.175 107.475 87.430 107.805 ;
        RECT 86.755 106.505 86.925 107.475 ;
        RECT 87.600 107.305 87.770 107.975 ;
        RECT 87.985 107.895 88.215 108.715 ;
        RECT 88.385 107.915 88.715 108.545 ;
        RECT 87.965 107.475 88.295 107.725 ;
        RECT 88.465 107.315 88.715 107.915 ;
        RECT 88.885 107.895 89.095 108.715 ;
        RECT 89.325 107.945 92.835 108.715 ;
        RECT 93.095 108.165 93.265 108.545 ;
        RECT 93.445 108.335 93.775 108.715 ;
        RECT 93.095 107.995 93.760 108.165 ;
        RECT 93.955 108.040 94.215 108.545 ;
        RECT 89.325 107.425 90.975 107.945 ;
        RECT 84.895 106.335 86.925 106.505 ;
        RECT 87.095 106.165 87.265 107.305 ;
        RECT 87.435 106.335 87.770 107.305 ;
        RECT 87.985 106.165 88.215 107.305 ;
        RECT 88.385 106.335 88.715 107.315 ;
        RECT 88.885 106.165 89.095 107.305 ;
        RECT 91.145 107.255 92.835 107.775 ;
        RECT 93.025 107.445 93.355 107.815 ;
        RECT 93.590 107.740 93.760 107.995 ;
        RECT 93.590 107.410 93.875 107.740 ;
        RECT 93.590 107.265 93.760 107.410 ;
        RECT 89.325 106.165 92.835 107.255 ;
        RECT 93.095 107.095 93.760 107.265 ;
        RECT 94.045 107.240 94.215 108.040 ;
        RECT 93.095 106.335 93.265 107.095 ;
        RECT 93.445 106.165 93.775 106.925 ;
        RECT 93.945 106.335 94.215 107.240 ;
        RECT 95.305 108.040 95.565 108.545 ;
        RECT 95.745 108.335 96.075 108.715 ;
        RECT 96.255 108.165 96.425 108.545 ;
        RECT 95.305 107.240 95.475 108.040 ;
        RECT 95.760 107.995 96.425 108.165 ;
        RECT 95.760 107.740 95.930 107.995 ;
        RECT 97.185 107.895 97.415 108.715 ;
        RECT 97.585 107.915 97.915 108.545 ;
        RECT 95.645 107.410 95.930 107.740 ;
        RECT 96.165 107.445 96.495 107.815 ;
        RECT 97.165 107.475 97.495 107.725 ;
        RECT 95.760 107.265 95.930 107.410 ;
        RECT 97.665 107.315 97.915 107.915 ;
        RECT 98.085 107.895 98.295 108.715 ;
        RECT 99.360 108.005 99.615 108.535 ;
        RECT 99.795 108.255 100.080 108.715 ;
        RECT 95.305 106.335 95.575 107.240 ;
        RECT 95.760 107.095 96.425 107.265 ;
        RECT 95.745 106.165 96.075 106.925 ;
        RECT 96.255 106.335 96.425 107.095 ;
        RECT 97.185 106.165 97.415 107.305 ;
        RECT 97.585 106.335 97.915 107.315 ;
        RECT 98.085 106.165 98.295 107.305 ;
        RECT 99.360 107.145 99.540 108.005 ;
        RECT 100.260 107.805 100.510 108.455 ;
        RECT 99.710 107.475 100.510 107.805 ;
        RECT 99.360 106.675 99.615 107.145 ;
        RECT 99.275 106.505 99.615 106.675 ;
        RECT 99.360 106.475 99.615 106.505 ;
        RECT 99.795 106.165 100.080 106.965 ;
        RECT 100.260 106.885 100.510 107.475 ;
        RECT 100.710 108.120 101.030 108.450 ;
        RECT 101.210 108.235 101.870 108.715 ;
        RECT 102.070 108.325 102.920 108.495 ;
        RECT 100.710 107.225 100.900 108.120 ;
        RECT 101.220 107.795 101.880 108.065 ;
        RECT 101.550 107.735 101.880 107.795 ;
        RECT 101.070 107.565 101.400 107.625 ;
        RECT 102.070 107.565 102.240 108.325 ;
        RECT 103.480 108.255 103.800 108.715 ;
        RECT 104.000 108.075 104.250 108.505 ;
        RECT 104.540 108.275 104.950 108.715 ;
        RECT 105.120 108.335 106.135 108.535 ;
        RECT 102.410 107.905 103.660 108.075 ;
        RECT 102.410 107.785 102.740 107.905 ;
        RECT 101.070 107.395 102.970 107.565 ;
        RECT 100.710 107.055 102.630 107.225 ;
        RECT 100.710 107.035 101.030 107.055 ;
        RECT 100.260 106.375 100.590 106.885 ;
        RECT 100.860 106.425 101.030 107.035 ;
        RECT 102.800 106.885 102.970 107.395 ;
        RECT 103.140 107.325 103.320 107.735 ;
        RECT 103.490 107.145 103.660 107.905 ;
        RECT 101.200 106.165 101.530 106.855 ;
        RECT 101.760 106.715 102.970 106.885 ;
        RECT 103.140 106.835 103.660 107.145 ;
        RECT 103.830 107.735 104.250 108.075 ;
        RECT 104.540 107.735 104.950 108.065 ;
        RECT 103.830 106.965 104.020 107.735 ;
        RECT 105.120 107.605 105.290 108.335 ;
        RECT 106.435 108.165 106.605 108.495 ;
        RECT 106.775 108.335 107.105 108.715 ;
        RECT 105.460 107.785 105.810 108.155 ;
        RECT 105.120 107.565 105.540 107.605 ;
        RECT 104.190 107.395 105.540 107.565 ;
        RECT 104.190 107.235 104.440 107.395 ;
        RECT 104.950 106.965 105.200 107.225 ;
        RECT 103.830 106.715 105.200 106.965 ;
        RECT 101.760 106.425 102.000 106.715 ;
        RECT 102.800 106.635 102.970 106.715 ;
        RECT 102.200 106.165 102.620 106.545 ;
        RECT 102.800 106.385 103.430 106.635 ;
        RECT 103.900 106.165 104.230 106.545 ;
        RECT 104.400 106.425 104.570 106.715 ;
        RECT 105.370 106.550 105.540 107.395 ;
        RECT 105.990 107.225 106.210 108.095 ;
        RECT 106.435 107.975 107.130 108.165 ;
        RECT 105.710 106.845 106.210 107.225 ;
        RECT 106.380 107.175 106.790 107.795 ;
        RECT 106.960 107.005 107.130 107.975 ;
        RECT 106.435 106.835 107.130 107.005 ;
        RECT 104.750 106.165 105.130 106.545 ;
        RECT 105.370 106.380 106.200 106.550 ;
        RECT 106.435 106.335 106.605 106.835 ;
        RECT 106.775 106.165 107.105 106.665 ;
        RECT 107.320 106.335 107.545 108.455 ;
        RECT 107.715 108.335 108.045 108.715 ;
        RECT 108.215 108.165 108.385 108.455 ;
        RECT 107.720 107.995 108.385 108.165 ;
        RECT 107.720 107.005 107.950 107.995 ;
        RECT 108.645 107.990 108.935 108.715 ;
        RECT 109.605 107.895 109.835 108.715 ;
        RECT 110.005 107.915 110.335 108.545 ;
        RECT 108.120 107.175 108.470 107.825 ;
        RECT 109.585 107.475 109.915 107.725 ;
        RECT 107.720 106.835 108.385 107.005 ;
        RECT 107.715 106.165 108.045 106.665 ;
        RECT 108.215 106.335 108.385 106.835 ;
        RECT 108.645 106.165 108.935 107.330 ;
        RECT 110.085 107.315 110.335 107.915 ;
        RECT 110.505 107.895 110.715 108.715 ;
        RECT 110.945 108.040 111.205 108.545 ;
        RECT 111.385 108.335 111.715 108.715 ;
        RECT 111.895 108.165 112.065 108.545 ;
        RECT 109.605 106.165 109.835 107.305 ;
        RECT 110.005 106.335 110.335 107.315 ;
        RECT 110.505 106.165 110.715 107.305 ;
        RECT 110.945 107.240 111.115 108.040 ;
        RECT 111.400 107.995 112.065 108.165 ;
        RECT 111.400 107.740 111.570 107.995 ;
        RECT 112.325 107.945 115.835 108.715 ;
        RECT 116.005 107.965 117.215 108.715 ;
        RECT 117.385 107.965 118.595 108.715 ;
        RECT 111.285 107.410 111.570 107.740 ;
        RECT 111.805 107.445 112.135 107.815 ;
        RECT 112.325 107.425 113.975 107.945 ;
        RECT 111.400 107.265 111.570 107.410 ;
        RECT 110.945 106.335 111.215 107.240 ;
        RECT 111.400 107.095 112.065 107.265 ;
        RECT 114.145 107.255 115.835 107.775 ;
        RECT 116.005 107.425 116.525 107.965 ;
        RECT 116.695 107.255 117.215 107.795 ;
        RECT 111.385 106.165 111.715 106.925 ;
        RECT 111.895 106.335 112.065 107.095 ;
        RECT 112.325 106.165 115.835 107.255 ;
        RECT 116.005 106.165 117.215 107.255 ;
        RECT 117.385 107.255 117.905 107.795 ;
        RECT 118.075 107.425 118.595 107.965 ;
        RECT 117.385 106.165 118.595 107.255 ;
        RECT 5.520 105.995 118.680 106.165 ;
        RECT 5.605 104.905 6.815 105.995 ;
        RECT 6.985 105.560 12.330 105.995 ;
        RECT 5.605 104.195 6.125 104.735 ;
        RECT 6.295 104.365 6.815 104.905 ;
        RECT 5.605 103.445 6.815 104.195 ;
        RECT 8.570 103.990 8.910 104.820 ;
        RECT 10.390 104.310 10.740 105.560 ;
        RECT 12.505 104.905 16.015 105.995 ;
        RECT 12.505 104.215 14.155 104.735 ;
        RECT 14.325 104.385 16.015 104.905 ;
        RECT 16.645 104.920 16.915 105.825 ;
        RECT 17.085 105.235 17.415 105.995 ;
        RECT 17.595 105.065 17.765 105.825 ;
        RECT 6.985 103.445 12.330 103.990 ;
        RECT 12.505 103.445 16.015 104.215 ;
        RECT 16.645 104.120 16.815 104.920 ;
        RECT 17.100 104.895 17.765 105.065 ;
        RECT 17.100 104.750 17.270 104.895 ;
        RECT 18.485 104.830 18.775 105.995 ;
        RECT 18.985 104.855 19.215 105.995 ;
        RECT 19.385 104.845 19.715 105.825 ;
        RECT 19.885 104.855 20.095 105.995 ;
        RECT 21.335 105.325 21.505 105.825 ;
        RECT 21.675 105.495 22.005 105.995 ;
        RECT 21.335 105.155 22.000 105.325 ;
        RECT 16.985 104.420 17.270 104.750 ;
        RECT 17.100 104.165 17.270 104.420 ;
        RECT 17.505 104.345 17.835 104.715 ;
        RECT 18.965 104.435 19.295 104.685 ;
        RECT 16.645 103.615 16.905 104.120 ;
        RECT 17.100 103.995 17.765 104.165 ;
        RECT 17.085 103.445 17.415 103.825 ;
        RECT 17.595 103.615 17.765 103.995 ;
        RECT 18.485 103.445 18.775 104.170 ;
        RECT 18.985 103.445 19.215 104.265 ;
        RECT 19.465 104.245 19.715 104.845 ;
        RECT 21.250 104.335 21.600 104.985 ;
        RECT 19.385 103.615 19.715 104.245 ;
        RECT 19.885 103.445 20.095 104.265 ;
        RECT 21.770 104.165 22.000 105.155 ;
        RECT 21.335 103.995 22.000 104.165 ;
        RECT 21.335 103.705 21.505 103.995 ;
        RECT 21.675 103.445 22.005 103.825 ;
        RECT 22.175 103.705 22.400 105.825 ;
        RECT 22.615 105.495 22.945 105.995 ;
        RECT 23.115 105.325 23.285 105.825 ;
        RECT 23.520 105.610 24.350 105.780 ;
        RECT 24.590 105.615 24.970 105.995 ;
        RECT 22.590 105.155 23.285 105.325 ;
        RECT 22.590 104.185 22.760 105.155 ;
        RECT 22.930 104.365 23.340 104.985 ;
        RECT 23.510 104.935 24.010 105.315 ;
        RECT 22.590 103.995 23.285 104.185 ;
        RECT 23.510 104.065 23.730 104.935 ;
        RECT 24.180 104.765 24.350 105.610 ;
        RECT 25.150 105.445 25.320 105.735 ;
        RECT 25.490 105.615 25.820 105.995 ;
        RECT 26.290 105.525 26.920 105.775 ;
        RECT 27.100 105.615 27.520 105.995 ;
        RECT 26.750 105.445 26.920 105.525 ;
        RECT 27.720 105.445 27.960 105.735 ;
        RECT 24.520 105.195 25.890 105.445 ;
        RECT 24.520 104.935 24.770 105.195 ;
        RECT 25.280 104.765 25.530 104.925 ;
        RECT 24.180 104.595 25.530 104.765 ;
        RECT 24.180 104.555 24.600 104.595 ;
        RECT 23.910 104.005 24.260 104.375 ;
        RECT 22.615 103.445 22.945 103.825 ;
        RECT 23.115 103.665 23.285 103.995 ;
        RECT 24.430 103.825 24.600 104.555 ;
        RECT 25.700 104.425 25.890 105.195 ;
        RECT 24.770 104.095 25.180 104.425 ;
        RECT 25.470 104.085 25.890 104.425 ;
        RECT 26.060 105.015 26.580 105.325 ;
        RECT 26.750 105.275 27.960 105.445 ;
        RECT 28.190 105.305 28.520 105.995 ;
        RECT 26.060 104.255 26.230 105.015 ;
        RECT 26.400 104.425 26.580 104.835 ;
        RECT 26.750 104.765 26.920 105.275 ;
        RECT 28.690 105.125 28.860 105.735 ;
        RECT 29.130 105.275 29.460 105.785 ;
        RECT 28.690 105.105 29.010 105.125 ;
        RECT 27.090 104.935 29.010 105.105 ;
        RECT 26.750 104.595 28.650 104.765 ;
        RECT 26.980 104.255 27.310 104.375 ;
        RECT 26.060 104.085 27.310 104.255 ;
        RECT 23.585 103.625 24.600 103.825 ;
        RECT 24.770 103.445 25.180 103.885 ;
        RECT 25.470 103.655 25.720 104.085 ;
        RECT 25.920 103.445 26.240 103.905 ;
        RECT 27.480 103.835 27.650 104.595 ;
        RECT 28.320 104.535 28.650 104.595 ;
        RECT 27.840 104.365 28.170 104.425 ;
        RECT 27.840 104.095 28.500 104.365 ;
        RECT 28.820 104.040 29.010 104.935 ;
        RECT 26.800 103.665 27.650 103.835 ;
        RECT 27.850 103.445 28.510 103.925 ;
        RECT 28.690 103.710 29.010 104.040 ;
        RECT 29.210 104.685 29.460 105.275 ;
        RECT 29.640 105.195 29.925 105.995 ;
        RECT 30.105 105.015 30.360 105.685 ;
        RECT 30.995 105.325 31.165 105.825 ;
        RECT 31.335 105.495 31.665 105.995 ;
        RECT 30.995 105.155 31.660 105.325 ;
        RECT 29.210 104.355 30.010 104.685 ;
        RECT 29.210 103.705 29.460 104.355 ;
        RECT 30.180 104.155 30.360 105.015 ;
        RECT 30.910 104.335 31.260 104.985 ;
        RECT 31.430 104.165 31.660 105.155 ;
        RECT 30.105 103.955 30.360 104.155 ;
        RECT 30.995 103.995 31.660 104.165 ;
        RECT 29.640 103.445 29.925 103.905 ;
        RECT 30.105 103.785 30.445 103.955 ;
        RECT 30.105 103.625 30.360 103.785 ;
        RECT 30.995 103.705 31.165 103.995 ;
        RECT 31.335 103.445 31.665 103.825 ;
        RECT 31.835 103.705 32.060 105.825 ;
        RECT 32.275 105.495 32.605 105.995 ;
        RECT 32.775 105.325 32.945 105.825 ;
        RECT 33.180 105.610 34.010 105.780 ;
        RECT 34.250 105.615 34.630 105.995 ;
        RECT 32.250 105.155 32.945 105.325 ;
        RECT 32.250 104.185 32.420 105.155 ;
        RECT 32.590 104.365 33.000 104.985 ;
        RECT 33.170 104.935 33.670 105.315 ;
        RECT 32.250 103.995 32.945 104.185 ;
        RECT 33.170 104.065 33.390 104.935 ;
        RECT 33.840 104.765 34.010 105.610 ;
        RECT 34.810 105.445 34.980 105.735 ;
        RECT 35.150 105.615 35.480 105.995 ;
        RECT 35.950 105.525 36.580 105.775 ;
        RECT 36.760 105.615 37.180 105.995 ;
        RECT 36.410 105.445 36.580 105.525 ;
        RECT 37.380 105.445 37.620 105.735 ;
        RECT 34.180 105.195 35.550 105.445 ;
        RECT 34.180 104.935 34.430 105.195 ;
        RECT 34.940 104.765 35.190 104.925 ;
        RECT 33.840 104.595 35.190 104.765 ;
        RECT 33.840 104.555 34.260 104.595 ;
        RECT 33.570 104.005 33.920 104.375 ;
        RECT 32.275 103.445 32.605 103.825 ;
        RECT 32.775 103.665 32.945 103.995 ;
        RECT 34.090 103.825 34.260 104.555 ;
        RECT 35.360 104.425 35.550 105.195 ;
        RECT 34.430 104.095 34.840 104.425 ;
        RECT 35.130 104.085 35.550 104.425 ;
        RECT 35.720 105.015 36.240 105.325 ;
        RECT 36.410 105.275 37.620 105.445 ;
        RECT 37.850 105.305 38.180 105.995 ;
        RECT 35.720 104.255 35.890 105.015 ;
        RECT 36.060 104.425 36.240 104.835 ;
        RECT 36.410 104.765 36.580 105.275 ;
        RECT 38.350 105.125 38.520 105.735 ;
        RECT 38.790 105.275 39.120 105.785 ;
        RECT 38.350 105.105 38.670 105.125 ;
        RECT 36.750 104.935 38.670 105.105 ;
        RECT 36.410 104.595 38.310 104.765 ;
        RECT 36.640 104.255 36.970 104.375 ;
        RECT 35.720 104.085 36.970 104.255 ;
        RECT 33.245 103.625 34.260 103.825 ;
        RECT 34.430 103.445 34.840 103.885 ;
        RECT 35.130 103.655 35.380 104.085 ;
        RECT 35.580 103.445 35.900 103.905 ;
        RECT 37.140 103.835 37.310 104.595 ;
        RECT 37.980 104.535 38.310 104.595 ;
        RECT 37.500 104.365 37.830 104.425 ;
        RECT 37.500 104.095 38.160 104.365 ;
        RECT 38.480 104.040 38.670 104.935 ;
        RECT 36.460 103.665 37.310 103.835 ;
        RECT 37.510 103.445 38.170 103.925 ;
        RECT 38.350 103.710 38.670 104.040 ;
        RECT 38.870 104.685 39.120 105.275 ;
        RECT 39.300 105.195 39.585 105.995 ;
        RECT 39.765 105.015 40.020 105.685 ;
        RECT 38.870 104.355 39.670 104.685 ;
        RECT 38.870 103.705 39.120 104.355 ;
        RECT 39.840 104.155 40.020 105.015 ;
        RECT 41.545 104.855 41.755 105.995 ;
        RECT 41.925 104.845 42.255 105.825 ;
        RECT 42.425 104.855 42.655 105.995 ;
        RECT 42.925 104.855 43.135 105.995 ;
        RECT 43.305 104.845 43.635 105.825 ;
        RECT 43.805 104.855 44.035 105.995 ;
        RECT 39.765 103.955 40.020 104.155 ;
        RECT 39.300 103.445 39.585 103.905 ;
        RECT 39.765 103.785 40.105 103.955 ;
        RECT 39.765 103.625 40.020 103.785 ;
        RECT 41.545 103.445 41.755 104.265 ;
        RECT 41.925 104.245 42.175 104.845 ;
        RECT 42.345 104.435 42.675 104.685 ;
        RECT 41.925 103.615 42.255 104.245 ;
        RECT 42.425 103.445 42.655 104.265 ;
        RECT 42.925 103.445 43.135 104.265 ;
        RECT 43.305 104.245 43.555 104.845 ;
        RECT 44.245 104.830 44.535 105.995 ;
        RECT 44.705 104.920 44.975 105.825 ;
        RECT 45.145 105.235 45.475 105.995 ;
        RECT 45.655 105.065 45.825 105.825 ;
        RECT 43.725 104.435 44.055 104.685 ;
        RECT 43.305 103.615 43.635 104.245 ;
        RECT 43.805 103.445 44.035 104.265 ;
        RECT 44.245 103.445 44.535 104.170 ;
        RECT 44.705 104.120 44.875 104.920 ;
        RECT 45.160 104.895 45.825 105.065 ;
        RECT 46.545 105.235 47.060 105.645 ;
        RECT 47.295 105.235 47.465 105.995 ;
        RECT 47.635 105.655 49.665 105.825 ;
        RECT 45.160 104.750 45.330 104.895 ;
        RECT 45.045 104.420 45.330 104.750 ;
        RECT 45.160 104.165 45.330 104.420 ;
        RECT 45.565 104.345 45.895 104.715 ;
        RECT 46.545 104.425 46.885 105.235 ;
        RECT 47.635 104.990 47.805 105.655 ;
        RECT 48.200 105.315 49.325 105.485 ;
        RECT 47.055 104.800 47.805 104.990 ;
        RECT 47.975 104.975 48.985 105.145 ;
        RECT 46.545 104.255 47.775 104.425 ;
        RECT 44.705 103.615 44.965 104.120 ;
        RECT 45.160 103.995 45.825 104.165 ;
        RECT 45.145 103.445 45.475 103.825 ;
        RECT 45.655 103.615 45.825 103.995 ;
        RECT 46.820 103.650 47.065 104.255 ;
        RECT 47.285 103.445 47.795 103.980 ;
        RECT 47.975 103.615 48.165 104.975 ;
        RECT 48.335 104.635 48.610 104.775 ;
        RECT 48.335 104.465 48.615 104.635 ;
        RECT 48.335 103.615 48.610 104.465 ;
        RECT 48.815 104.175 48.985 104.975 ;
        RECT 49.155 104.185 49.325 105.315 ;
        RECT 49.495 104.685 49.665 105.655 ;
        RECT 49.835 104.855 50.005 105.995 ;
        RECT 50.175 104.855 50.510 105.825 ;
        RECT 50.775 105.325 50.945 105.825 ;
        RECT 51.115 105.495 51.445 105.995 ;
        RECT 50.775 105.155 51.440 105.325 ;
        RECT 49.495 104.355 49.690 104.685 ;
        RECT 49.915 104.355 50.170 104.685 ;
        RECT 49.915 104.185 50.085 104.355 ;
        RECT 50.340 104.185 50.510 104.855 ;
        RECT 50.690 104.335 51.040 104.985 ;
        RECT 49.155 104.015 50.085 104.185 ;
        RECT 49.155 103.980 49.330 104.015 ;
        RECT 48.800 103.615 49.330 103.980 ;
        RECT 49.755 103.445 50.085 103.845 ;
        RECT 50.255 103.615 50.510 104.185 ;
        RECT 51.210 104.165 51.440 105.155 ;
        RECT 50.775 103.995 51.440 104.165 ;
        RECT 50.775 103.705 50.945 103.995 ;
        RECT 51.115 103.445 51.445 103.825 ;
        RECT 51.615 103.705 51.840 105.825 ;
        RECT 52.055 105.495 52.385 105.995 ;
        RECT 52.555 105.325 52.725 105.825 ;
        RECT 52.960 105.610 53.790 105.780 ;
        RECT 54.030 105.615 54.410 105.995 ;
        RECT 52.030 105.155 52.725 105.325 ;
        RECT 52.030 104.185 52.200 105.155 ;
        RECT 52.370 104.365 52.780 104.985 ;
        RECT 52.950 104.935 53.450 105.315 ;
        RECT 52.030 103.995 52.725 104.185 ;
        RECT 52.950 104.065 53.170 104.935 ;
        RECT 53.620 104.765 53.790 105.610 ;
        RECT 54.590 105.445 54.760 105.735 ;
        RECT 54.930 105.615 55.260 105.995 ;
        RECT 55.730 105.525 56.360 105.775 ;
        RECT 56.540 105.615 56.960 105.995 ;
        RECT 56.190 105.445 56.360 105.525 ;
        RECT 57.160 105.445 57.400 105.735 ;
        RECT 53.960 105.195 55.330 105.445 ;
        RECT 53.960 104.935 54.210 105.195 ;
        RECT 54.720 104.765 54.970 104.925 ;
        RECT 53.620 104.595 54.970 104.765 ;
        RECT 53.620 104.555 54.040 104.595 ;
        RECT 53.350 104.005 53.700 104.375 ;
        RECT 52.055 103.445 52.385 103.825 ;
        RECT 52.555 103.665 52.725 103.995 ;
        RECT 53.870 103.825 54.040 104.555 ;
        RECT 55.140 104.425 55.330 105.195 ;
        RECT 54.210 104.095 54.620 104.425 ;
        RECT 54.910 104.085 55.330 104.425 ;
        RECT 55.500 105.015 56.020 105.325 ;
        RECT 56.190 105.275 57.400 105.445 ;
        RECT 57.630 105.305 57.960 105.995 ;
        RECT 55.500 104.255 55.670 105.015 ;
        RECT 55.840 104.425 56.020 104.835 ;
        RECT 56.190 104.765 56.360 105.275 ;
        RECT 58.130 105.125 58.300 105.735 ;
        RECT 58.570 105.275 58.900 105.785 ;
        RECT 58.130 105.105 58.450 105.125 ;
        RECT 56.530 104.935 58.450 105.105 ;
        RECT 56.190 104.595 58.090 104.765 ;
        RECT 56.420 104.255 56.750 104.375 ;
        RECT 55.500 104.085 56.750 104.255 ;
        RECT 53.025 103.625 54.040 103.825 ;
        RECT 54.210 103.445 54.620 103.885 ;
        RECT 54.910 103.655 55.160 104.085 ;
        RECT 55.360 103.445 55.680 103.905 ;
        RECT 56.920 103.835 57.090 104.595 ;
        RECT 57.760 104.535 58.090 104.595 ;
        RECT 57.280 104.365 57.610 104.425 ;
        RECT 57.280 104.095 57.940 104.365 ;
        RECT 58.260 104.040 58.450 104.935 ;
        RECT 56.240 103.665 57.090 103.835 ;
        RECT 57.290 103.445 57.950 103.925 ;
        RECT 58.130 103.710 58.450 104.040 ;
        RECT 58.650 104.685 58.900 105.275 ;
        RECT 59.080 105.195 59.365 105.995 ;
        RECT 59.545 105.015 59.800 105.685 ;
        RECT 60.435 105.325 60.605 105.825 ;
        RECT 60.775 105.495 61.105 105.995 ;
        RECT 60.435 105.155 61.100 105.325 ;
        RECT 58.650 104.355 59.450 104.685 ;
        RECT 58.650 103.705 58.900 104.355 ;
        RECT 59.620 104.155 59.800 105.015 ;
        RECT 60.350 104.335 60.700 104.985 ;
        RECT 60.870 104.165 61.100 105.155 ;
        RECT 59.545 103.955 59.800 104.155 ;
        RECT 60.435 103.995 61.100 104.165 ;
        RECT 59.080 103.445 59.365 103.905 ;
        RECT 59.545 103.785 59.885 103.955 ;
        RECT 59.545 103.625 59.800 103.785 ;
        RECT 60.435 103.705 60.605 103.995 ;
        RECT 60.775 103.445 61.105 103.825 ;
        RECT 61.275 103.705 61.500 105.825 ;
        RECT 61.715 105.495 62.045 105.995 ;
        RECT 62.215 105.325 62.385 105.825 ;
        RECT 62.620 105.610 63.450 105.780 ;
        RECT 63.690 105.615 64.070 105.995 ;
        RECT 61.690 105.155 62.385 105.325 ;
        RECT 61.690 104.185 61.860 105.155 ;
        RECT 62.030 104.365 62.440 104.985 ;
        RECT 62.610 104.935 63.110 105.315 ;
        RECT 61.690 103.995 62.385 104.185 ;
        RECT 62.610 104.065 62.830 104.935 ;
        RECT 63.280 104.765 63.450 105.610 ;
        RECT 64.250 105.445 64.420 105.735 ;
        RECT 64.590 105.615 64.920 105.995 ;
        RECT 65.390 105.525 66.020 105.775 ;
        RECT 66.200 105.615 66.620 105.995 ;
        RECT 65.850 105.445 66.020 105.525 ;
        RECT 66.820 105.445 67.060 105.735 ;
        RECT 63.620 105.195 64.990 105.445 ;
        RECT 63.620 104.935 63.870 105.195 ;
        RECT 64.380 104.765 64.630 104.925 ;
        RECT 63.280 104.595 64.630 104.765 ;
        RECT 63.280 104.555 63.700 104.595 ;
        RECT 63.010 104.005 63.360 104.375 ;
        RECT 61.715 103.445 62.045 103.825 ;
        RECT 62.215 103.665 62.385 103.995 ;
        RECT 63.530 103.825 63.700 104.555 ;
        RECT 64.800 104.425 64.990 105.195 ;
        RECT 63.870 104.095 64.280 104.425 ;
        RECT 64.570 104.085 64.990 104.425 ;
        RECT 65.160 105.015 65.680 105.325 ;
        RECT 65.850 105.275 67.060 105.445 ;
        RECT 67.290 105.305 67.620 105.995 ;
        RECT 65.160 104.255 65.330 105.015 ;
        RECT 65.500 104.425 65.680 104.835 ;
        RECT 65.850 104.765 66.020 105.275 ;
        RECT 67.790 105.125 67.960 105.735 ;
        RECT 68.230 105.275 68.560 105.785 ;
        RECT 67.790 105.105 68.110 105.125 ;
        RECT 66.190 104.935 68.110 105.105 ;
        RECT 65.850 104.595 67.750 104.765 ;
        RECT 66.080 104.255 66.410 104.375 ;
        RECT 65.160 104.085 66.410 104.255 ;
        RECT 62.685 103.625 63.700 103.825 ;
        RECT 63.870 103.445 64.280 103.885 ;
        RECT 64.570 103.655 64.820 104.085 ;
        RECT 65.020 103.445 65.340 103.905 ;
        RECT 66.580 103.835 66.750 104.595 ;
        RECT 67.420 104.535 67.750 104.595 ;
        RECT 66.940 104.365 67.270 104.425 ;
        RECT 66.940 104.095 67.600 104.365 ;
        RECT 67.920 104.040 68.110 104.935 ;
        RECT 65.900 103.665 66.750 103.835 ;
        RECT 66.950 103.445 67.610 103.925 ;
        RECT 67.790 103.710 68.110 104.040 ;
        RECT 68.310 104.685 68.560 105.275 ;
        RECT 68.740 105.195 69.025 105.995 ;
        RECT 69.205 105.015 69.460 105.685 ;
        RECT 68.310 104.355 69.110 104.685 ;
        RECT 68.310 103.705 68.560 104.355 ;
        RECT 69.280 104.155 69.460 105.015 ;
        RECT 70.005 104.830 70.295 105.995 ;
        RECT 70.525 104.855 70.735 105.995 ;
        RECT 70.905 104.845 71.235 105.825 ;
        RECT 71.405 104.855 71.635 105.995 ;
        RECT 71.845 104.905 75.355 105.995 ;
        RECT 76.535 105.325 76.705 105.825 ;
        RECT 76.875 105.495 77.205 105.995 ;
        RECT 76.535 105.155 77.200 105.325 ;
        RECT 69.205 103.955 69.460 104.155 ;
        RECT 68.740 103.445 69.025 103.905 ;
        RECT 69.205 103.785 69.545 103.955 ;
        RECT 69.205 103.625 69.460 103.785 ;
        RECT 70.005 103.445 70.295 104.170 ;
        RECT 70.525 103.445 70.735 104.265 ;
        RECT 70.905 104.245 71.155 104.845 ;
        RECT 71.325 104.435 71.655 104.685 ;
        RECT 70.905 103.615 71.235 104.245 ;
        RECT 71.405 103.445 71.635 104.265 ;
        RECT 71.845 104.215 73.495 104.735 ;
        RECT 73.665 104.385 75.355 104.905 ;
        RECT 76.450 104.335 76.800 104.985 ;
        RECT 71.845 103.445 75.355 104.215 ;
        RECT 76.970 104.165 77.200 105.155 ;
        RECT 76.535 103.995 77.200 104.165 ;
        RECT 76.535 103.705 76.705 103.995 ;
        RECT 76.875 103.445 77.205 103.825 ;
        RECT 77.375 103.705 77.600 105.825 ;
        RECT 77.815 105.495 78.145 105.995 ;
        RECT 78.315 105.325 78.485 105.825 ;
        RECT 78.720 105.610 79.550 105.780 ;
        RECT 79.790 105.615 80.170 105.995 ;
        RECT 77.790 105.155 78.485 105.325 ;
        RECT 77.790 104.185 77.960 105.155 ;
        RECT 78.130 104.365 78.540 104.985 ;
        RECT 78.710 104.935 79.210 105.315 ;
        RECT 77.790 103.995 78.485 104.185 ;
        RECT 78.710 104.065 78.930 104.935 ;
        RECT 79.380 104.765 79.550 105.610 ;
        RECT 80.350 105.445 80.520 105.735 ;
        RECT 80.690 105.615 81.020 105.995 ;
        RECT 81.490 105.525 82.120 105.775 ;
        RECT 82.300 105.615 82.720 105.995 ;
        RECT 81.950 105.445 82.120 105.525 ;
        RECT 82.920 105.445 83.160 105.735 ;
        RECT 79.720 105.195 81.090 105.445 ;
        RECT 79.720 104.935 79.970 105.195 ;
        RECT 80.480 104.765 80.730 104.925 ;
        RECT 79.380 104.595 80.730 104.765 ;
        RECT 79.380 104.555 79.800 104.595 ;
        RECT 79.110 104.005 79.460 104.375 ;
        RECT 77.815 103.445 78.145 103.825 ;
        RECT 78.315 103.665 78.485 103.995 ;
        RECT 79.630 103.825 79.800 104.555 ;
        RECT 80.900 104.425 81.090 105.195 ;
        RECT 79.970 104.095 80.380 104.425 ;
        RECT 80.670 104.085 81.090 104.425 ;
        RECT 81.260 105.015 81.780 105.325 ;
        RECT 81.950 105.275 83.160 105.445 ;
        RECT 83.390 105.305 83.720 105.995 ;
        RECT 81.260 104.255 81.430 105.015 ;
        RECT 81.600 104.425 81.780 104.835 ;
        RECT 81.950 104.765 82.120 105.275 ;
        RECT 83.890 105.125 84.060 105.735 ;
        RECT 84.330 105.275 84.660 105.785 ;
        RECT 83.890 105.105 84.210 105.125 ;
        RECT 82.290 104.935 84.210 105.105 ;
        RECT 81.950 104.595 83.850 104.765 ;
        RECT 82.180 104.255 82.510 104.375 ;
        RECT 81.260 104.085 82.510 104.255 ;
        RECT 78.785 103.625 79.800 103.825 ;
        RECT 79.970 103.445 80.380 103.885 ;
        RECT 80.670 103.655 80.920 104.085 ;
        RECT 81.120 103.445 81.440 103.905 ;
        RECT 82.680 103.835 82.850 104.595 ;
        RECT 83.520 104.535 83.850 104.595 ;
        RECT 83.040 104.365 83.370 104.425 ;
        RECT 83.040 104.095 83.700 104.365 ;
        RECT 84.020 104.040 84.210 104.935 ;
        RECT 82.000 103.665 82.850 103.835 ;
        RECT 83.050 103.445 83.710 103.925 ;
        RECT 83.890 103.710 84.210 104.040 ;
        RECT 84.410 104.685 84.660 105.275 ;
        RECT 84.840 105.195 85.125 105.995 ;
        RECT 85.305 105.655 85.560 105.685 ;
        RECT 85.305 105.485 85.645 105.655 ;
        RECT 85.305 105.015 85.560 105.485 ;
        RECT 86.195 105.325 86.365 105.825 ;
        RECT 86.535 105.495 86.865 105.995 ;
        RECT 86.195 105.155 86.860 105.325 ;
        RECT 84.410 104.355 85.210 104.685 ;
        RECT 84.410 103.705 84.660 104.355 ;
        RECT 85.380 104.155 85.560 105.015 ;
        RECT 86.110 104.335 86.460 104.985 ;
        RECT 86.630 104.165 86.860 105.155 ;
        RECT 84.840 103.445 85.125 103.905 ;
        RECT 85.305 103.625 85.560 104.155 ;
        RECT 86.195 103.995 86.860 104.165 ;
        RECT 86.195 103.705 86.365 103.995 ;
        RECT 86.535 103.445 86.865 103.825 ;
        RECT 87.035 103.705 87.260 105.825 ;
        RECT 87.475 105.495 87.805 105.995 ;
        RECT 87.975 105.325 88.145 105.825 ;
        RECT 88.380 105.610 89.210 105.780 ;
        RECT 89.450 105.615 89.830 105.995 ;
        RECT 87.450 105.155 88.145 105.325 ;
        RECT 87.450 104.185 87.620 105.155 ;
        RECT 87.790 104.365 88.200 104.985 ;
        RECT 88.370 104.935 88.870 105.315 ;
        RECT 87.450 103.995 88.145 104.185 ;
        RECT 88.370 104.065 88.590 104.935 ;
        RECT 89.040 104.765 89.210 105.610 ;
        RECT 90.010 105.445 90.180 105.735 ;
        RECT 90.350 105.615 90.680 105.995 ;
        RECT 91.150 105.525 91.780 105.775 ;
        RECT 91.960 105.615 92.380 105.995 ;
        RECT 91.610 105.445 91.780 105.525 ;
        RECT 92.580 105.445 92.820 105.735 ;
        RECT 89.380 105.195 90.750 105.445 ;
        RECT 89.380 104.935 89.630 105.195 ;
        RECT 90.140 104.765 90.390 104.925 ;
        RECT 89.040 104.595 90.390 104.765 ;
        RECT 89.040 104.555 89.460 104.595 ;
        RECT 88.770 104.005 89.120 104.375 ;
        RECT 87.475 103.445 87.805 103.825 ;
        RECT 87.975 103.665 88.145 103.995 ;
        RECT 89.290 103.825 89.460 104.555 ;
        RECT 90.560 104.425 90.750 105.195 ;
        RECT 89.630 104.095 90.040 104.425 ;
        RECT 90.330 104.085 90.750 104.425 ;
        RECT 90.920 105.015 91.440 105.325 ;
        RECT 91.610 105.275 92.820 105.445 ;
        RECT 93.050 105.305 93.380 105.995 ;
        RECT 90.920 104.255 91.090 105.015 ;
        RECT 91.260 104.425 91.440 104.835 ;
        RECT 91.610 104.765 91.780 105.275 ;
        RECT 93.550 105.125 93.720 105.735 ;
        RECT 93.990 105.275 94.320 105.785 ;
        RECT 93.550 105.105 93.870 105.125 ;
        RECT 91.950 104.935 93.870 105.105 ;
        RECT 91.610 104.595 93.510 104.765 ;
        RECT 91.840 104.255 92.170 104.375 ;
        RECT 90.920 104.085 92.170 104.255 ;
        RECT 88.445 103.625 89.460 103.825 ;
        RECT 89.630 103.445 90.040 103.885 ;
        RECT 90.330 103.655 90.580 104.085 ;
        RECT 90.780 103.445 91.100 103.905 ;
        RECT 92.340 103.835 92.510 104.595 ;
        RECT 93.180 104.535 93.510 104.595 ;
        RECT 92.700 104.365 93.030 104.425 ;
        RECT 92.700 104.095 93.360 104.365 ;
        RECT 93.680 104.040 93.870 104.935 ;
        RECT 91.660 103.665 92.510 103.835 ;
        RECT 92.710 103.445 93.370 103.925 ;
        RECT 93.550 103.710 93.870 104.040 ;
        RECT 94.070 104.685 94.320 105.275 ;
        RECT 94.500 105.195 94.785 105.995 ;
        RECT 94.965 105.015 95.220 105.685 ;
        RECT 94.070 104.355 94.870 104.685 ;
        RECT 94.070 103.705 94.320 104.355 ;
        RECT 95.040 104.155 95.220 105.015 ;
        RECT 95.765 104.830 96.055 105.995 ;
        RECT 96.600 105.015 96.855 105.685 ;
        RECT 97.035 105.195 97.320 105.995 ;
        RECT 97.500 105.275 97.830 105.785 ;
        RECT 94.965 103.955 95.220 104.155 ;
        RECT 94.500 103.445 94.785 103.905 ;
        RECT 94.965 103.785 95.305 103.955 ;
        RECT 94.965 103.625 95.220 103.785 ;
        RECT 95.765 103.445 96.055 104.170 ;
        RECT 96.600 104.155 96.780 105.015 ;
        RECT 97.500 104.685 97.750 105.275 ;
        RECT 98.100 105.125 98.270 105.735 ;
        RECT 98.440 105.305 98.770 105.995 ;
        RECT 99.000 105.445 99.240 105.735 ;
        RECT 99.440 105.615 99.860 105.995 ;
        RECT 100.040 105.525 100.670 105.775 ;
        RECT 101.140 105.615 101.470 105.995 ;
        RECT 100.040 105.445 100.210 105.525 ;
        RECT 101.640 105.445 101.810 105.735 ;
        RECT 101.990 105.615 102.370 105.995 ;
        RECT 102.610 105.610 103.440 105.780 ;
        RECT 99.000 105.275 100.210 105.445 ;
        RECT 96.950 104.355 97.750 104.685 ;
        RECT 96.600 103.955 96.855 104.155 ;
        RECT 96.515 103.785 96.855 103.955 ;
        RECT 96.600 103.625 96.855 103.785 ;
        RECT 97.035 103.445 97.320 103.905 ;
        RECT 97.500 103.705 97.750 104.355 ;
        RECT 97.950 105.105 98.270 105.125 ;
        RECT 97.950 104.935 99.870 105.105 ;
        RECT 97.950 104.040 98.140 104.935 ;
        RECT 100.040 104.765 100.210 105.275 ;
        RECT 100.380 105.015 100.900 105.325 ;
        RECT 98.310 104.595 100.210 104.765 ;
        RECT 98.310 104.535 98.640 104.595 ;
        RECT 98.790 104.365 99.120 104.425 ;
        RECT 98.460 104.095 99.120 104.365 ;
        RECT 97.950 103.710 98.270 104.040 ;
        RECT 98.450 103.445 99.110 103.925 ;
        RECT 99.310 103.835 99.480 104.595 ;
        RECT 100.380 104.425 100.560 104.835 ;
        RECT 99.650 104.255 99.980 104.375 ;
        RECT 100.730 104.255 100.900 105.015 ;
        RECT 99.650 104.085 100.900 104.255 ;
        RECT 101.070 105.195 102.440 105.445 ;
        RECT 101.070 104.425 101.260 105.195 ;
        RECT 102.190 104.935 102.440 105.195 ;
        RECT 101.430 104.765 101.680 104.925 ;
        RECT 102.610 104.765 102.780 105.610 ;
        RECT 103.675 105.325 103.845 105.825 ;
        RECT 104.015 105.495 104.345 105.995 ;
        RECT 102.950 104.935 103.450 105.315 ;
        RECT 103.675 105.155 104.370 105.325 ;
        RECT 101.430 104.595 102.780 104.765 ;
        RECT 102.360 104.555 102.780 104.595 ;
        RECT 101.070 104.085 101.490 104.425 ;
        RECT 101.780 104.095 102.190 104.425 ;
        RECT 99.310 103.665 100.160 103.835 ;
        RECT 100.720 103.445 101.040 103.905 ;
        RECT 101.240 103.655 101.490 104.085 ;
        RECT 101.780 103.445 102.190 103.885 ;
        RECT 102.360 103.825 102.530 104.555 ;
        RECT 102.700 104.005 103.050 104.375 ;
        RECT 103.230 104.065 103.450 104.935 ;
        RECT 103.620 104.365 104.030 104.985 ;
        RECT 104.200 104.185 104.370 105.155 ;
        RECT 103.675 103.995 104.370 104.185 ;
        RECT 102.360 103.625 103.375 103.825 ;
        RECT 103.675 103.665 103.845 103.995 ;
        RECT 104.015 103.445 104.345 103.825 ;
        RECT 104.560 103.705 104.785 105.825 ;
        RECT 104.955 105.495 105.285 105.995 ;
        RECT 105.455 105.325 105.625 105.825 ;
        RECT 104.960 105.155 105.625 105.325 ;
        RECT 105.975 105.325 106.145 105.825 ;
        RECT 106.315 105.495 106.645 105.995 ;
        RECT 105.975 105.155 106.640 105.325 ;
        RECT 104.960 104.165 105.190 105.155 ;
        RECT 105.360 104.335 105.710 104.985 ;
        RECT 105.890 104.335 106.240 104.985 ;
        RECT 106.410 104.165 106.640 105.155 ;
        RECT 104.960 103.995 105.625 104.165 ;
        RECT 104.955 103.445 105.285 103.825 ;
        RECT 105.455 103.705 105.625 103.995 ;
        RECT 105.975 103.995 106.640 104.165 ;
        RECT 105.975 103.705 106.145 103.995 ;
        RECT 106.315 103.445 106.645 103.825 ;
        RECT 106.815 103.705 107.040 105.825 ;
        RECT 107.255 105.495 107.585 105.995 ;
        RECT 107.755 105.325 107.925 105.825 ;
        RECT 108.160 105.610 108.990 105.780 ;
        RECT 109.230 105.615 109.610 105.995 ;
        RECT 107.230 105.155 107.925 105.325 ;
        RECT 107.230 104.185 107.400 105.155 ;
        RECT 107.570 104.365 107.980 104.985 ;
        RECT 108.150 104.935 108.650 105.315 ;
        RECT 107.230 103.995 107.925 104.185 ;
        RECT 108.150 104.065 108.370 104.935 ;
        RECT 108.820 104.765 108.990 105.610 ;
        RECT 109.790 105.445 109.960 105.735 ;
        RECT 110.130 105.615 110.460 105.995 ;
        RECT 110.930 105.525 111.560 105.775 ;
        RECT 111.740 105.615 112.160 105.995 ;
        RECT 111.390 105.445 111.560 105.525 ;
        RECT 112.360 105.445 112.600 105.735 ;
        RECT 109.160 105.195 110.530 105.445 ;
        RECT 109.160 104.935 109.410 105.195 ;
        RECT 109.920 104.765 110.170 104.925 ;
        RECT 108.820 104.595 110.170 104.765 ;
        RECT 108.820 104.555 109.240 104.595 ;
        RECT 108.550 104.005 108.900 104.375 ;
        RECT 107.255 103.445 107.585 103.825 ;
        RECT 107.755 103.665 107.925 103.995 ;
        RECT 109.070 103.825 109.240 104.555 ;
        RECT 110.340 104.425 110.530 105.195 ;
        RECT 109.410 104.095 109.820 104.425 ;
        RECT 110.110 104.085 110.530 104.425 ;
        RECT 110.700 105.015 111.220 105.325 ;
        RECT 111.390 105.275 112.600 105.445 ;
        RECT 112.830 105.305 113.160 105.995 ;
        RECT 110.700 104.255 110.870 105.015 ;
        RECT 111.040 104.425 111.220 104.835 ;
        RECT 111.390 104.765 111.560 105.275 ;
        RECT 113.330 105.125 113.500 105.735 ;
        RECT 113.770 105.275 114.100 105.785 ;
        RECT 113.330 105.105 113.650 105.125 ;
        RECT 111.730 104.935 113.650 105.105 ;
        RECT 111.390 104.595 113.290 104.765 ;
        RECT 111.620 104.255 111.950 104.375 ;
        RECT 110.700 104.085 111.950 104.255 ;
        RECT 108.225 103.625 109.240 103.825 ;
        RECT 109.410 103.445 109.820 103.885 ;
        RECT 110.110 103.655 110.360 104.085 ;
        RECT 110.560 103.445 110.880 103.905 ;
        RECT 112.120 103.835 112.290 104.595 ;
        RECT 112.960 104.535 113.290 104.595 ;
        RECT 112.480 104.365 112.810 104.425 ;
        RECT 112.480 104.095 113.140 104.365 ;
        RECT 113.460 104.040 113.650 104.935 ;
        RECT 111.440 103.665 112.290 103.835 ;
        RECT 112.490 103.445 113.150 103.925 ;
        RECT 113.330 103.710 113.650 104.040 ;
        RECT 113.850 104.685 114.100 105.275 ;
        RECT 114.280 105.195 114.565 105.995 ;
        RECT 114.745 105.015 115.000 105.685 ;
        RECT 113.850 104.355 114.650 104.685 ;
        RECT 113.850 103.705 114.100 104.355 ;
        RECT 114.820 104.155 115.000 105.015 ;
        RECT 115.585 104.855 115.815 105.995 ;
        RECT 115.985 104.845 116.315 105.825 ;
        RECT 116.485 104.855 116.695 105.995 ;
        RECT 117.385 104.905 118.595 105.995 ;
        RECT 115.565 104.435 115.895 104.685 ;
        RECT 114.745 103.955 115.000 104.155 ;
        RECT 114.280 103.445 114.565 103.905 ;
        RECT 114.745 103.785 115.085 103.955 ;
        RECT 114.745 103.625 115.000 103.785 ;
        RECT 115.585 103.445 115.815 104.265 ;
        RECT 116.065 104.245 116.315 104.845 ;
        RECT 117.385 104.365 117.905 104.905 ;
        RECT 115.985 103.615 116.315 104.245 ;
        RECT 116.485 103.445 116.695 104.265 ;
        RECT 118.075 104.195 118.595 104.735 ;
        RECT 117.385 103.445 118.595 104.195 ;
        RECT 5.520 103.275 118.680 103.445 ;
        RECT 5.605 102.525 6.815 103.275 ;
        RECT 5.605 101.985 6.125 102.525 ;
        RECT 6.985 102.505 10.495 103.275 ;
        RECT 11.585 102.600 11.845 103.105 ;
        RECT 12.025 102.895 12.355 103.275 ;
        RECT 12.535 102.725 12.705 103.105 ;
        RECT 6.295 101.815 6.815 102.355 ;
        RECT 6.985 101.985 8.635 102.505 ;
        RECT 8.805 101.815 10.495 102.335 ;
        RECT 5.605 100.725 6.815 101.815 ;
        RECT 6.985 100.725 10.495 101.815 ;
        RECT 11.585 101.800 11.755 102.600 ;
        RECT 12.040 102.555 12.705 102.725 ;
        RECT 12.040 102.300 12.210 102.555 ;
        RECT 13.485 102.455 13.695 103.275 ;
        RECT 13.865 102.475 14.195 103.105 ;
        RECT 11.925 101.970 12.210 102.300 ;
        RECT 12.445 102.005 12.775 102.375 ;
        RECT 12.040 101.825 12.210 101.970 ;
        RECT 13.865 101.875 14.115 102.475 ;
        RECT 14.365 102.455 14.595 103.275 ;
        RECT 14.895 102.725 15.065 103.015 ;
        RECT 15.235 102.895 15.565 103.275 ;
        RECT 14.895 102.555 15.560 102.725 ;
        RECT 14.285 102.035 14.615 102.285 ;
        RECT 11.585 100.895 11.855 101.800 ;
        RECT 12.040 101.655 12.705 101.825 ;
        RECT 12.025 100.725 12.355 101.485 ;
        RECT 12.535 100.895 12.705 101.655 ;
        RECT 13.485 100.725 13.695 101.865 ;
        RECT 13.865 100.895 14.195 101.875 ;
        RECT 14.365 100.725 14.595 101.865 ;
        RECT 14.810 101.735 15.160 102.385 ;
        RECT 15.330 101.565 15.560 102.555 ;
        RECT 14.895 101.395 15.560 101.565 ;
        RECT 14.895 100.895 15.065 101.395 ;
        RECT 15.235 100.725 15.565 101.225 ;
        RECT 15.735 100.895 15.960 103.015 ;
        RECT 16.175 102.895 16.505 103.275 ;
        RECT 16.675 102.725 16.845 103.055 ;
        RECT 17.145 102.895 18.160 103.095 ;
        RECT 16.150 102.535 16.845 102.725 ;
        RECT 16.150 101.565 16.320 102.535 ;
        RECT 16.490 101.735 16.900 102.355 ;
        RECT 17.070 101.785 17.290 102.655 ;
        RECT 17.470 102.345 17.820 102.715 ;
        RECT 17.990 102.165 18.160 102.895 ;
        RECT 18.330 102.835 18.740 103.275 ;
        RECT 19.030 102.635 19.280 103.065 ;
        RECT 19.480 102.815 19.800 103.275 ;
        RECT 20.360 102.885 21.210 103.055 ;
        RECT 18.330 102.295 18.740 102.625 ;
        RECT 19.030 102.295 19.450 102.635 ;
        RECT 17.740 102.125 18.160 102.165 ;
        RECT 17.740 101.955 19.090 102.125 ;
        RECT 16.150 101.395 16.845 101.565 ;
        RECT 17.070 101.405 17.570 101.785 ;
        RECT 16.175 100.725 16.505 101.225 ;
        RECT 16.675 100.895 16.845 101.395 ;
        RECT 17.740 101.110 17.910 101.955 ;
        RECT 18.840 101.795 19.090 101.955 ;
        RECT 18.080 101.525 18.330 101.785 ;
        RECT 19.260 101.525 19.450 102.295 ;
        RECT 18.080 101.275 19.450 101.525 ;
        RECT 19.620 102.465 20.870 102.635 ;
        RECT 19.620 101.705 19.790 102.465 ;
        RECT 20.540 102.345 20.870 102.465 ;
        RECT 19.960 101.885 20.140 102.295 ;
        RECT 21.040 102.125 21.210 102.885 ;
        RECT 21.410 102.795 22.070 103.275 ;
        RECT 22.250 102.680 22.570 103.010 ;
        RECT 21.400 102.355 22.060 102.625 ;
        RECT 21.400 102.295 21.730 102.355 ;
        RECT 21.880 102.125 22.210 102.185 ;
        RECT 20.310 101.955 22.210 102.125 ;
        RECT 19.620 101.395 20.140 101.705 ;
        RECT 20.310 101.445 20.480 101.955 ;
        RECT 22.380 101.785 22.570 102.680 ;
        RECT 20.650 101.615 22.570 101.785 ;
        RECT 22.250 101.595 22.570 101.615 ;
        RECT 22.770 102.365 23.020 103.015 ;
        RECT 23.200 102.815 23.485 103.275 ;
        RECT 23.665 102.565 23.920 103.095 ;
        RECT 22.770 102.035 23.570 102.365 ;
        RECT 20.310 101.275 21.520 101.445 ;
        RECT 17.080 100.940 17.910 101.110 ;
        RECT 18.150 100.725 18.530 101.105 ;
        RECT 18.710 100.985 18.880 101.275 ;
        RECT 20.310 101.195 20.480 101.275 ;
        RECT 19.050 100.725 19.380 101.105 ;
        RECT 19.850 100.945 20.480 101.195 ;
        RECT 20.660 100.725 21.080 101.105 ;
        RECT 21.280 100.985 21.520 101.275 ;
        RECT 21.750 100.725 22.080 101.415 ;
        RECT 22.250 100.985 22.420 101.595 ;
        RECT 22.770 101.445 23.020 102.035 ;
        RECT 23.740 101.915 23.920 102.565 ;
        RECT 24.470 102.535 24.725 103.105 ;
        RECT 24.895 102.875 25.225 103.275 ;
        RECT 25.650 102.740 26.180 103.105 ;
        RECT 25.650 102.705 25.825 102.740 ;
        RECT 24.895 102.535 25.825 102.705 ;
        RECT 26.370 102.595 26.645 103.105 ;
        RECT 23.740 101.745 24.005 101.915 ;
        RECT 24.470 101.865 24.640 102.535 ;
        RECT 24.895 102.365 25.065 102.535 ;
        RECT 24.810 102.035 25.065 102.365 ;
        RECT 25.290 102.035 25.485 102.365 ;
        RECT 23.740 101.705 23.920 101.745 ;
        RECT 22.690 100.935 23.020 101.445 ;
        RECT 23.200 100.725 23.485 101.525 ;
        RECT 23.665 101.035 23.920 101.705 ;
        RECT 24.470 100.895 24.805 101.865 ;
        RECT 24.975 100.725 25.145 101.865 ;
        RECT 25.315 101.065 25.485 102.035 ;
        RECT 25.655 101.405 25.825 102.535 ;
        RECT 25.995 101.745 26.165 102.545 ;
        RECT 26.365 102.425 26.645 102.595 ;
        RECT 26.370 101.945 26.645 102.425 ;
        RECT 26.815 101.745 27.005 103.105 ;
        RECT 27.185 102.740 27.695 103.275 ;
        RECT 27.915 102.465 28.160 103.070 ;
        RECT 27.205 102.295 28.435 102.465 ;
        RECT 28.665 102.455 28.875 103.275 ;
        RECT 29.045 102.475 29.375 103.105 ;
        RECT 25.995 101.575 27.005 101.745 ;
        RECT 27.175 101.730 27.925 101.920 ;
        RECT 25.655 101.235 26.780 101.405 ;
        RECT 27.175 101.065 27.345 101.730 ;
        RECT 28.095 101.485 28.435 102.295 ;
        RECT 29.045 101.875 29.295 102.475 ;
        RECT 29.545 102.455 29.775 103.275 ;
        RECT 29.985 102.525 31.195 103.275 ;
        RECT 31.365 102.550 31.655 103.275 ;
        RECT 31.830 102.535 32.085 103.105 ;
        RECT 32.255 102.875 32.585 103.275 ;
        RECT 33.010 102.740 33.540 103.105 ;
        RECT 33.010 102.705 33.185 102.740 ;
        RECT 32.255 102.535 33.185 102.705 ;
        RECT 29.465 102.035 29.795 102.285 ;
        RECT 29.985 101.985 30.505 102.525 ;
        RECT 25.315 100.895 27.345 101.065 ;
        RECT 27.515 100.725 27.685 101.485 ;
        RECT 27.920 101.075 28.435 101.485 ;
        RECT 28.665 100.725 28.875 101.865 ;
        RECT 29.045 100.895 29.375 101.875 ;
        RECT 29.545 100.725 29.775 101.865 ;
        RECT 30.675 101.815 31.195 102.355 ;
        RECT 29.985 100.725 31.195 101.815 ;
        RECT 31.365 100.725 31.655 101.890 ;
        RECT 31.830 101.865 32.000 102.535 ;
        RECT 32.255 102.365 32.425 102.535 ;
        RECT 32.170 102.035 32.425 102.365 ;
        RECT 32.650 102.035 32.845 102.365 ;
        RECT 31.830 100.895 32.165 101.865 ;
        RECT 32.335 100.725 32.505 101.865 ;
        RECT 32.675 101.065 32.845 102.035 ;
        RECT 33.015 101.405 33.185 102.535 ;
        RECT 33.355 101.745 33.525 102.545 ;
        RECT 33.730 102.255 34.005 103.105 ;
        RECT 33.725 102.085 34.005 102.255 ;
        RECT 33.730 101.945 34.005 102.085 ;
        RECT 34.175 101.745 34.365 103.105 ;
        RECT 34.545 102.740 35.055 103.275 ;
        RECT 35.275 102.465 35.520 103.070 ;
        RECT 35.965 102.505 37.635 103.275 ;
        RECT 34.565 102.295 35.795 102.465 ;
        RECT 33.355 101.575 34.365 101.745 ;
        RECT 34.535 101.730 35.285 101.920 ;
        RECT 33.015 101.235 34.140 101.405 ;
        RECT 34.535 101.065 34.705 101.730 ;
        RECT 35.455 101.485 35.795 102.295 ;
        RECT 35.965 101.985 36.715 102.505 ;
        RECT 38.540 102.465 38.785 103.070 ;
        RECT 39.005 102.740 39.515 103.275 ;
        RECT 36.885 101.815 37.635 102.335 ;
        RECT 32.675 100.895 34.705 101.065 ;
        RECT 34.875 100.725 35.045 101.485 ;
        RECT 35.280 101.075 35.795 101.485 ;
        RECT 35.965 100.725 37.635 101.815 ;
        RECT 38.265 102.295 39.495 102.465 ;
        RECT 38.265 101.485 38.605 102.295 ;
        RECT 38.775 101.730 39.525 101.920 ;
        RECT 38.265 101.075 38.780 101.485 ;
        RECT 39.015 100.725 39.185 101.485 ;
        RECT 39.355 101.065 39.525 101.730 ;
        RECT 39.695 101.745 39.885 103.105 ;
        RECT 40.055 102.935 40.330 103.105 ;
        RECT 40.055 102.765 40.335 102.935 ;
        RECT 40.055 101.945 40.330 102.765 ;
        RECT 40.520 102.740 41.050 103.105 ;
        RECT 41.475 102.875 41.805 103.275 ;
        RECT 40.875 102.705 41.050 102.740 ;
        RECT 40.535 101.745 40.705 102.545 ;
        RECT 39.695 101.575 40.705 101.745 ;
        RECT 40.875 102.535 41.805 102.705 ;
        RECT 41.975 102.535 42.230 103.105 ;
        RECT 42.405 102.730 47.750 103.275 ;
        RECT 40.875 101.405 41.045 102.535 ;
        RECT 41.635 102.365 41.805 102.535 ;
        RECT 39.920 101.235 41.045 101.405 ;
        RECT 41.215 102.035 41.410 102.365 ;
        RECT 41.635 102.035 41.890 102.365 ;
        RECT 41.215 101.065 41.385 102.035 ;
        RECT 42.060 101.865 42.230 102.535 ;
        RECT 43.990 101.900 44.330 102.730 ;
        RECT 47.925 102.600 48.185 103.105 ;
        RECT 48.365 102.895 48.695 103.275 ;
        RECT 48.875 102.725 49.045 103.105 ;
        RECT 39.355 100.895 41.385 101.065 ;
        RECT 41.555 100.725 41.725 101.865 ;
        RECT 41.895 100.895 42.230 101.865 ;
        RECT 45.810 101.160 46.160 102.410 ;
        RECT 47.925 101.800 48.095 102.600 ;
        RECT 48.380 102.555 49.045 102.725 ;
        RECT 48.380 102.300 48.550 102.555 ;
        RECT 49.805 102.455 50.035 103.275 ;
        RECT 50.205 102.475 50.535 103.105 ;
        RECT 48.265 101.970 48.550 102.300 ;
        RECT 48.785 102.005 49.115 102.375 ;
        RECT 49.785 102.035 50.115 102.285 ;
        RECT 48.380 101.825 48.550 101.970 ;
        RECT 50.285 101.875 50.535 102.475 ;
        RECT 50.705 102.455 50.915 103.275 ;
        RECT 51.235 102.725 51.405 103.105 ;
        RECT 51.585 102.895 51.915 103.275 ;
        RECT 51.235 102.555 51.900 102.725 ;
        RECT 52.095 102.600 52.355 103.105 ;
        RECT 51.165 102.005 51.495 102.375 ;
        RECT 51.730 102.300 51.900 102.555 ;
        RECT 42.405 100.725 47.750 101.160 ;
        RECT 47.925 100.895 48.195 101.800 ;
        RECT 48.380 101.655 49.045 101.825 ;
        RECT 48.365 100.725 48.695 101.485 ;
        RECT 48.875 100.895 49.045 101.655 ;
        RECT 49.805 100.725 50.035 101.865 ;
        RECT 50.205 100.895 50.535 101.875 ;
        RECT 51.730 101.970 52.015 102.300 ;
        RECT 50.705 100.725 50.915 101.865 ;
        RECT 51.730 101.825 51.900 101.970 ;
        RECT 51.235 101.655 51.900 101.825 ;
        RECT 52.185 101.800 52.355 102.600 ;
        RECT 51.235 100.895 51.405 101.655 ;
        RECT 51.585 100.725 51.915 101.485 ;
        RECT 52.085 100.895 52.355 101.800 ;
        RECT 52.530 102.535 52.785 103.105 ;
        RECT 52.955 102.875 53.285 103.275 ;
        RECT 53.710 102.740 54.240 103.105 ;
        RECT 54.430 102.935 54.705 103.105 ;
        RECT 54.425 102.765 54.705 102.935 ;
        RECT 53.710 102.705 53.885 102.740 ;
        RECT 52.955 102.535 53.885 102.705 ;
        RECT 52.530 101.865 52.700 102.535 ;
        RECT 52.955 102.365 53.125 102.535 ;
        RECT 52.870 102.035 53.125 102.365 ;
        RECT 53.350 102.035 53.545 102.365 ;
        RECT 52.530 100.895 52.865 101.865 ;
        RECT 53.035 100.725 53.205 101.865 ;
        RECT 53.375 101.065 53.545 102.035 ;
        RECT 53.715 101.405 53.885 102.535 ;
        RECT 54.055 101.745 54.225 102.545 ;
        RECT 54.430 101.945 54.705 102.765 ;
        RECT 54.875 101.745 55.065 103.105 ;
        RECT 55.245 102.740 55.755 103.275 ;
        RECT 55.975 102.465 56.220 103.070 ;
        RECT 57.125 102.550 57.415 103.275 ;
        RECT 55.265 102.295 56.495 102.465 ;
        RECT 57.645 102.455 57.855 103.275 ;
        RECT 58.025 102.475 58.355 103.105 ;
        RECT 54.055 101.575 55.065 101.745 ;
        RECT 55.235 101.730 55.985 101.920 ;
        RECT 53.715 101.235 54.840 101.405 ;
        RECT 55.235 101.065 55.405 101.730 ;
        RECT 56.155 101.485 56.495 102.295 ;
        RECT 53.375 100.895 55.405 101.065 ;
        RECT 55.575 100.725 55.745 101.485 ;
        RECT 55.980 101.075 56.495 101.485 ;
        RECT 57.125 100.725 57.415 101.890 ;
        RECT 58.025 101.875 58.275 102.475 ;
        RECT 58.525 102.455 58.755 103.275 ;
        RECT 58.965 102.505 62.475 103.275 ;
        RECT 63.195 102.725 63.365 103.105 ;
        RECT 63.545 102.895 63.875 103.275 ;
        RECT 63.195 102.555 63.860 102.725 ;
        RECT 64.055 102.600 64.315 103.105 ;
        RECT 58.445 102.035 58.775 102.285 ;
        RECT 58.965 101.985 60.615 102.505 ;
        RECT 57.645 100.725 57.855 101.865 ;
        RECT 58.025 100.895 58.355 101.875 ;
        RECT 58.525 100.725 58.755 101.865 ;
        RECT 60.785 101.815 62.475 102.335 ;
        RECT 63.125 102.005 63.455 102.375 ;
        RECT 63.690 102.300 63.860 102.555 ;
        RECT 63.690 101.970 63.975 102.300 ;
        RECT 63.690 101.825 63.860 101.970 ;
        RECT 58.965 100.725 62.475 101.815 ;
        RECT 63.195 101.655 63.860 101.825 ;
        RECT 64.145 101.800 64.315 102.600 ;
        RECT 64.575 102.725 64.745 103.015 ;
        RECT 64.915 102.895 65.245 103.275 ;
        RECT 64.575 102.555 65.240 102.725 ;
        RECT 63.195 100.895 63.365 101.655 ;
        RECT 63.545 100.725 63.875 101.485 ;
        RECT 64.045 100.895 64.315 101.800 ;
        RECT 64.490 101.735 64.840 102.385 ;
        RECT 65.010 101.565 65.240 102.555 ;
        RECT 64.575 101.395 65.240 101.565 ;
        RECT 64.575 100.895 64.745 101.395 ;
        RECT 64.915 100.725 65.245 101.225 ;
        RECT 65.415 100.895 65.640 103.015 ;
        RECT 65.855 102.895 66.185 103.275 ;
        RECT 66.355 102.725 66.525 103.055 ;
        RECT 66.825 102.895 67.840 103.095 ;
        RECT 65.830 102.535 66.525 102.725 ;
        RECT 65.830 101.565 66.000 102.535 ;
        RECT 66.170 101.735 66.580 102.355 ;
        RECT 66.750 101.785 66.970 102.655 ;
        RECT 67.150 102.345 67.500 102.715 ;
        RECT 67.670 102.165 67.840 102.895 ;
        RECT 68.010 102.835 68.420 103.275 ;
        RECT 68.710 102.635 68.960 103.065 ;
        RECT 69.160 102.815 69.480 103.275 ;
        RECT 70.040 102.885 70.890 103.055 ;
        RECT 68.010 102.295 68.420 102.625 ;
        RECT 68.710 102.295 69.130 102.635 ;
        RECT 67.420 102.125 67.840 102.165 ;
        RECT 67.420 101.955 68.770 102.125 ;
        RECT 65.830 101.395 66.525 101.565 ;
        RECT 66.750 101.405 67.250 101.785 ;
        RECT 65.855 100.725 66.185 101.225 ;
        RECT 66.355 100.895 66.525 101.395 ;
        RECT 67.420 101.110 67.590 101.955 ;
        RECT 68.520 101.795 68.770 101.955 ;
        RECT 67.760 101.525 68.010 101.785 ;
        RECT 68.940 101.525 69.130 102.295 ;
        RECT 67.760 101.275 69.130 101.525 ;
        RECT 69.300 102.465 70.550 102.635 ;
        RECT 69.300 101.705 69.470 102.465 ;
        RECT 70.220 102.345 70.550 102.465 ;
        RECT 69.640 101.885 69.820 102.295 ;
        RECT 70.720 102.125 70.890 102.885 ;
        RECT 71.090 102.795 71.750 103.275 ;
        RECT 71.930 102.680 72.250 103.010 ;
        RECT 71.080 102.355 71.740 102.625 ;
        RECT 71.080 102.295 71.410 102.355 ;
        RECT 71.560 102.125 71.890 102.185 ;
        RECT 69.990 101.955 71.890 102.125 ;
        RECT 69.300 101.395 69.820 101.705 ;
        RECT 69.990 101.445 70.160 101.955 ;
        RECT 72.060 101.785 72.250 102.680 ;
        RECT 70.330 101.615 72.250 101.785 ;
        RECT 71.930 101.595 72.250 101.615 ;
        RECT 72.450 102.365 72.700 103.015 ;
        RECT 72.880 102.815 73.165 103.275 ;
        RECT 73.345 102.565 73.600 103.095 ;
        RECT 72.450 102.035 73.250 102.365 ;
        RECT 69.990 101.275 71.200 101.445 ;
        RECT 66.760 100.940 67.590 101.110 ;
        RECT 67.830 100.725 68.210 101.105 ;
        RECT 68.390 100.985 68.560 101.275 ;
        RECT 69.990 101.195 70.160 101.275 ;
        RECT 68.730 100.725 69.060 101.105 ;
        RECT 69.530 100.945 70.160 101.195 ;
        RECT 70.340 100.725 70.760 101.105 ;
        RECT 70.960 100.985 71.200 101.275 ;
        RECT 71.430 100.725 71.760 101.415 ;
        RECT 71.930 100.985 72.100 101.595 ;
        RECT 72.450 101.445 72.700 102.035 ;
        RECT 73.420 101.705 73.600 102.565 ;
        RECT 75.105 102.455 75.335 103.275 ;
        RECT 75.505 102.475 75.835 103.105 ;
        RECT 75.085 102.035 75.415 102.285 ;
        RECT 75.585 101.875 75.835 102.475 ;
        RECT 76.005 102.455 76.215 103.275 ;
        RECT 77.455 102.625 77.625 103.105 ;
        RECT 77.805 102.795 78.045 103.275 ;
        RECT 78.295 102.625 78.465 103.105 ;
        RECT 78.635 102.795 78.965 103.275 ;
        RECT 79.135 102.625 79.305 103.105 ;
        RECT 77.455 102.455 78.090 102.625 ;
        RECT 78.295 102.455 79.305 102.625 ;
        RECT 79.475 102.475 79.805 103.275 ;
        RECT 80.125 102.525 81.335 103.275 ;
        RECT 77.920 102.285 78.090 102.455 ;
        RECT 77.370 102.045 77.750 102.285 ;
        RECT 77.920 102.115 78.420 102.285 ;
        RECT 78.810 102.255 79.305 102.455 ;
        RECT 77.920 101.875 78.090 102.115 ;
        RECT 78.805 102.085 79.305 102.255 ;
        RECT 78.810 101.915 79.305 102.085 ;
        RECT 80.125 101.985 80.645 102.525 ;
        RECT 81.565 102.455 81.775 103.275 ;
        RECT 81.945 102.475 82.275 103.105 ;
        RECT 72.370 100.935 72.700 101.445 ;
        RECT 72.880 100.725 73.165 101.525 ;
        RECT 73.345 101.235 73.600 101.705 ;
        RECT 73.345 101.065 73.685 101.235 ;
        RECT 73.345 101.035 73.600 101.065 ;
        RECT 75.105 100.725 75.335 101.865 ;
        RECT 75.505 100.895 75.835 101.875 ;
        RECT 76.005 100.725 76.215 101.865 ;
        RECT 77.375 101.705 78.090 101.875 ;
        RECT 78.295 101.745 79.305 101.915 ;
        RECT 77.375 100.895 77.705 101.705 ;
        RECT 77.875 100.725 78.115 101.525 ;
        RECT 78.295 100.895 78.465 101.745 ;
        RECT 78.635 100.725 78.965 101.525 ;
        RECT 79.135 100.895 79.305 101.745 ;
        RECT 79.475 100.725 79.805 101.875 ;
        RECT 80.815 101.815 81.335 102.355 ;
        RECT 81.945 101.875 82.195 102.475 ;
        RECT 82.445 102.455 82.675 103.275 ;
        RECT 82.885 102.550 83.175 103.275 ;
        RECT 83.350 102.535 83.605 103.105 ;
        RECT 83.775 102.875 84.105 103.275 ;
        RECT 84.530 102.740 85.060 103.105 ;
        RECT 84.530 102.705 84.705 102.740 ;
        RECT 83.775 102.535 84.705 102.705 ;
        RECT 82.365 102.035 82.695 102.285 ;
        RECT 80.125 100.725 81.335 101.815 ;
        RECT 81.565 100.725 81.775 101.865 ;
        RECT 81.945 100.895 82.275 101.875 ;
        RECT 82.445 100.725 82.675 101.865 ;
        RECT 82.885 100.725 83.175 101.890 ;
        RECT 83.350 101.865 83.520 102.535 ;
        RECT 83.775 102.365 83.945 102.535 ;
        RECT 83.690 102.035 83.945 102.365 ;
        RECT 84.170 102.035 84.365 102.365 ;
        RECT 83.350 100.895 83.685 101.865 ;
        RECT 83.855 100.725 84.025 101.865 ;
        RECT 84.195 101.065 84.365 102.035 ;
        RECT 84.535 101.405 84.705 102.535 ;
        RECT 84.875 101.745 85.045 102.545 ;
        RECT 85.250 102.255 85.525 103.105 ;
        RECT 85.245 102.085 85.525 102.255 ;
        RECT 85.250 101.945 85.525 102.085 ;
        RECT 85.695 101.745 85.885 103.105 ;
        RECT 86.065 102.740 86.575 103.275 ;
        RECT 86.795 102.465 87.040 103.070 ;
        RECT 87.575 102.725 87.745 103.105 ;
        RECT 87.925 102.895 88.255 103.275 ;
        RECT 87.575 102.555 88.240 102.725 ;
        RECT 88.435 102.600 88.695 103.105 ;
        RECT 86.085 102.295 87.315 102.465 ;
        RECT 84.875 101.575 85.885 101.745 ;
        RECT 86.055 101.730 86.805 101.920 ;
        RECT 84.535 101.235 85.660 101.405 ;
        RECT 86.055 101.065 86.225 101.730 ;
        RECT 86.975 101.485 87.315 102.295 ;
        RECT 87.505 102.005 87.835 102.375 ;
        RECT 88.070 102.300 88.240 102.555 ;
        RECT 88.070 101.970 88.355 102.300 ;
        RECT 88.070 101.825 88.240 101.970 ;
        RECT 84.195 100.895 86.225 101.065 ;
        RECT 86.395 100.725 86.565 101.485 ;
        RECT 86.800 101.075 87.315 101.485 ;
        RECT 87.575 101.655 88.240 101.825 ;
        RECT 88.525 101.800 88.695 102.600 ;
        RECT 89.600 102.465 89.845 103.070 ;
        RECT 90.065 102.740 90.575 103.275 ;
        RECT 87.575 100.895 87.745 101.655 ;
        RECT 87.925 100.725 88.255 101.485 ;
        RECT 88.425 100.895 88.695 101.800 ;
        RECT 89.325 102.295 90.555 102.465 ;
        RECT 89.325 101.485 89.665 102.295 ;
        RECT 89.835 101.730 90.585 101.920 ;
        RECT 89.325 101.075 89.840 101.485 ;
        RECT 90.075 100.725 90.245 101.485 ;
        RECT 90.415 101.065 90.585 101.730 ;
        RECT 90.755 101.745 90.945 103.105 ;
        RECT 91.115 102.255 91.390 103.105 ;
        RECT 91.580 102.740 92.110 103.105 ;
        RECT 92.535 102.875 92.865 103.275 ;
        RECT 91.935 102.705 92.110 102.740 ;
        RECT 91.115 102.085 91.395 102.255 ;
        RECT 91.115 101.945 91.390 102.085 ;
        RECT 91.595 101.745 91.765 102.545 ;
        RECT 90.755 101.575 91.765 101.745 ;
        RECT 91.935 102.535 92.865 102.705 ;
        RECT 93.035 102.535 93.290 103.105 ;
        RECT 93.555 102.725 93.725 103.015 ;
        RECT 93.895 102.895 94.225 103.275 ;
        RECT 93.555 102.555 94.220 102.725 ;
        RECT 91.935 101.405 92.105 102.535 ;
        RECT 92.695 102.365 92.865 102.535 ;
        RECT 90.980 101.235 92.105 101.405 ;
        RECT 92.275 102.035 92.470 102.365 ;
        RECT 92.695 102.035 92.950 102.365 ;
        RECT 92.275 101.065 92.445 102.035 ;
        RECT 93.120 101.865 93.290 102.535 ;
        RECT 90.415 100.895 92.445 101.065 ;
        RECT 92.615 100.725 92.785 101.865 ;
        RECT 92.955 100.895 93.290 101.865 ;
        RECT 93.470 101.735 93.820 102.385 ;
        RECT 93.990 101.565 94.220 102.555 ;
        RECT 93.555 101.395 94.220 101.565 ;
        RECT 93.555 100.895 93.725 101.395 ;
        RECT 93.895 100.725 94.225 101.225 ;
        RECT 94.395 100.895 94.620 103.015 ;
        RECT 94.835 102.895 95.165 103.275 ;
        RECT 95.335 102.725 95.505 103.055 ;
        RECT 95.805 102.895 96.820 103.095 ;
        RECT 94.810 102.535 95.505 102.725 ;
        RECT 94.810 101.565 94.980 102.535 ;
        RECT 95.150 101.735 95.560 102.355 ;
        RECT 95.730 101.785 95.950 102.655 ;
        RECT 96.130 102.345 96.480 102.715 ;
        RECT 96.650 102.165 96.820 102.895 ;
        RECT 96.990 102.835 97.400 103.275 ;
        RECT 97.690 102.635 97.940 103.065 ;
        RECT 98.140 102.815 98.460 103.275 ;
        RECT 99.020 102.885 99.870 103.055 ;
        RECT 96.990 102.295 97.400 102.625 ;
        RECT 97.690 102.295 98.110 102.635 ;
        RECT 96.400 102.125 96.820 102.165 ;
        RECT 96.400 101.955 97.750 102.125 ;
        RECT 94.810 101.395 95.505 101.565 ;
        RECT 95.730 101.405 96.230 101.785 ;
        RECT 94.835 100.725 95.165 101.225 ;
        RECT 95.335 100.895 95.505 101.395 ;
        RECT 96.400 101.110 96.570 101.955 ;
        RECT 97.500 101.795 97.750 101.955 ;
        RECT 96.740 101.525 96.990 101.785 ;
        RECT 97.920 101.525 98.110 102.295 ;
        RECT 96.740 101.275 98.110 101.525 ;
        RECT 98.280 102.465 99.530 102.635 ;
        RECT 98.280 101.705 98.450 102.465 ;
        RECT 99.200 102.345 99.530 102.465 ;
        RECT 98.620 101.885 98.800 102.295 ;
        RECT 99.700 102.125 99.870 102.885 ;
        RECT 100.070 102.795 100.730 103.275 ;
        RECT 100.910 102.680 101.230 103.010 ;
        RECT 100.060 102.355 100.720 102.625 ;
        RECT 100.060 102.295 100.390 102.355 ;
        RECT 100.540 102.125 100.870 102.185 ;
        RECT 98.970 101.955 100.870 102.125 ;
        RECT 98.280 101.395 98.800 101.705 ;
        RECT 98.970 101.445 99.140 101.955 ;
        RECT 101.040 101.785 101.230 102.680 ;
        RECT 99.310 101.615 101.230 101.785 ;
        RECT 100.910 101.595 101.230 101.615 ;
        RECT 101.430 102.365 101.680 103.015 ;
        RECT 101.860 102.815 102.145 103.275 ;
        RECT 102.325 102.565 102.580 103.095 ;
        RECT 101.430 102.035 102.230 102.365 ;
        RECT 98.970 101.275 100.180 101.445 ;
        RECT 95.740 100.940 96.570 101.110 ;
        RECT 96.810 100.725 97.190 101.105 ;
        RECT 97.370 100.985 97.540 101.275 ;
        RECT 98.970 101.195 99.140 101.275 ;
        RECT 97.710 100.725 98.040 101.105 ;
        RECT 98.510 100.945 99.140 101.195 ;
        RECT 99.320 100.725 99.740 101.105 ;
        RECT 99.940 100.985 100.180 101.275 ;
        RECT 100.410 100.725 100.740 101.415 ;
        RECT 100.910 100.985 101.080 101.595 ;
        RECT 101.430 101.445 101.680 102.035 ;
        RECT 102.400 101.705 102.580 102.565 ;
        RECT 103.125 102.505 105.715 103.275 ;
        RECT 105.975 102.725 106.145 103.105 ;
        RECT 106.325 102.895 106.655 103.275 ;
        RECT 105.975 102.555 106.640 102.725 ;
        RECT 106.835 102.600 107.095 103.105 ;
        RECT 103.125 101.985 104.335 102.505 ;
        RECT 104.505 101.815 105.715 102.335 ;
        RECT 105.905 102.005 106.235 102.375 ;
        RECT 106.470 102.300 106.640 102.555 ;
        RECT 106.470 101.970 106.755 102.300 ;
        RECT 106.470 101.825 106.640 101.970 ;
        RECT 101.350 100.935 101.680 101.445 ;
        RECT 101.860 100.725 102.145 101.525 ;
        RECT 102.325 101.235 102.580 101.705 ;
        RECT 102.325 101.065 102.665 101.235 ;
        RECT 102.325 101.035 102.580 101.065 ;
        RECT 103.125 100.725 105.715 101.815 ;
        RECT 105.975 101.655 106.640 101.825 ;
        RECT 106.925 101.800 107.095 102.600 ;
        RECT 107.265 102.525 108.475 103.275 ;
        RECT 108.645 102.550 108.935 103.275 ;
        RECT 107.265 101.985 107.785 102.525 ;
        RECT 109.380 102.465 109.625 103.070 ;
        RECT 109.845 102.740 110.355 103.275 ;
        RECT 107.955 101.815 108.475 102.355 ;
        RECT 109.105 102.295 110.335 102.465 ;
        RECT 105.975 100.895 106.145 101.655 ;
        RECT 106.325 100.725 106.655 101.485 ;
        RECT 106.825 100.895 107.095 101.800 ;
        RECT 107.265 100.725 108.475 101.815 ;
        RECT 108.645 100.725 108.935 101.890 ;
        RECT 109.105 101.485 109.445 102.295 ;
        RECT 109.615 101.730 110.365 101.920 ;
        RECT 109.105 101.075 109.620 101.485 ;
        RECT 109.855 100.725 110.025 101.485 ;
        RECT 110.195 101.065 110.365 101.730 ;
        RECT 110.535 101.745 110.725 103.105 ;
        RECT 110.895 102.595 111.170 103.105 ;
        RECT 111.360 102.740 111.890 103.105 ;
        RECT 112.315 102.875 112.645 103.275 ;
        RECT 111.715 102.705 111.890 102.740 ;
        RECT 110.895 102.425 111.175 102.595 ;
        RECT 110.895 101.945 111.170 102.425 ;
        RECT 111.375 101.745 111.545 102.545 ;
        RECT 110.535 101.575 111.545 101.745 ;
        RECT 111.715 102.535 112.645 102.705 ;
        RECT 112.815 102.535 113.070 103.105 ;
        RECT 111.715 101.405 111.885 102.535 ;
        RECT 112.475 102.365 112.645 102.535 ;
        RECT 110.760 101.235 111.885 101.405 ;
        RECT 112.055 102.035 112.250 102.365 ;
        RECT 112.475 102.035 112.730 102.365 ;
        RECT 112.055 101.065 112.225 102.035 ;
        RECT 112.900 101.865 113.070 102.535 ;
        RECT 113.245 102.505 116.755 103.275 ;
        RECT 117.385 102.525 118.595 103.275 ;
        RECT 113.245 101.985 114.895 102.505 ;
        RECT 110.195 100.895 112.225 101.065 ;
        RECT 112.395 100.725 112.565 101.865 ;
        RECT 112.735 100.895 113.070 101.865 ;
        RECT 115.065 101.815 116.755 102.335 ;
        RECT 113.245 100.725 116.755 101.815 ;
        RECT 117.385 101.815 117.905 102.355 ;
        RECT 118.075 101.985 118.595 102.525 ;
        RECT 117.385 100.725 118.595 101.815 ;
        RECT 5.520 100.555 118.680 100.725 ;
        RECT 5.605 99.465 6.815 100.555 ;
        RECT 6.985 99.465 8.195 100.555 ;
        RECT 8.455 99.885 8.625 100.385 ;
        RECT 8.795 100.055 9.125 100.555 ;
        RECT 8.455 99.715 9.120 99.885 ;
        RECT 5.605 98.755 6.125 99.295 ;
        RECT 6.295 98.925 6.815 99.465 ;
        RECT 6.985 98.755 7.505 99.295 ;
        RECT 7.675 98.925 8.195 99.465 ;
        RECT 8.370 98.895 8.720 99.545 ;
        RECT 5.605 98.005 6.815 98.755 ;
        RECT 6.985 98.005 8.195 98.755 ;
        RECT 8.890 98.725 9.120 99.715 ;
        RECT 8.455 98.555 9.120 98.725 ;
        RECT 8.455 98.265 8.625 98.555 ;
        RECT 8.795 98.005 9.125 98.385 ;
        RECT 9.295 98.265 9.520 100.385 ;
        RECT 9.735 100.055 10.065 100.555 ;
        RECT 10.235 99.885 10.405 100.385 ;
        RECT 10.640 100.170 11.470 100.340 ;
        RECT 11.710 100.175 12.090 100.555 ;
        RECT 9.710 99.715 10.405 99.885 ;
        RECT 9.710 98.745 9.880 99.715 ;
        RECT 10.050 98.925 10.460 99.545 ;
        RECT 10.630 99.495 11.130 99.875 ;
        RECT 9.710 98.555 10.405 98.745 ;
        RECT 10.630 98.625 10.850 99.495 ;
        RECT 11.300 99.325 11.470 100.170 ;
        RECT 12.270 100.005 12.440 100.295 ;
        RECT 12.610 100.175 12.940 100.555 ;
        RECT 13.410 100.085 14.040 100.335 ;
        RECT 14.220 100.175 14.640 100.555 ;
        RECT 13.870 100.005 14.040 100.085 ;
        RECT 14.840 100.005 15.080 100.295 ;
        RECT 11.640 99.755 13.010 100.005 ;
        RECT 11.640 99.495 11.890 99.755 ;
        RECT 12.400 99.325 12.650 99.485 ;
        RECT 11.300 99.155 12.650 99.325 ;
        RECT 11.300 99.115 11.720 99.155 ;
        RECT 11.030 98.565 11.380 98.935 ;
        RECT 9.735 98.005 10.065 98.385 ;
        RECT 10.235 98.225 10.405 98.555 ;
        RECT 11.550 98.385 11.720 99.115 ;
        RECT 12.820 98.985 13.010 99.755 ;
        RECT 11.890 98.655 12.300 98.985 ;
        RECT 12.590 98.645 13.010 98.985 ;
        RECT 13.180 99.575 13.700 99.885 ;
        RECT 13.870 99.835 15.080 100.005 ;
        RECT 15.310 99.865 15.640 100.555 ;
        RECT 13.180 98.815 13.350 99.575 ;
        RECT 13.520 98.985 13.700 99.395 ;
        RECT 13.870 99.325 14.040 99.835 ;
        RECT 15.810 99.685 15.980 100.295 ;
        RECT 16.250 99.835 16.580 100.345 ;
        RECT 15.810 99.665 16.130 99.685 ;
        RECT 14.210 99.495 16.130 99.665 ;
        RECT 13.870 99.155 15.770 99.325 ;
        RECT 14.100 98.815 14.430 98.935 ;
        RECT 13.180 98.645 14.430 98.815 ;
        RECT 10.705 98.185 11.720 98.385 ;
        RECT 11.890 98.005 12.300 98.445 ;
        RECT 12.590 98.215 12.840 98.645 ;
        RECT 13.040 98.005 13.360 98.465 ;
        RECT 14.600 98.395 14.770 99.155 ;
        RECT 15.440 99.095 15.770 99.155 ;
        RECT 14.960 98.925 15.290 98.985 ;
        RECT 14.960 98.655 15.620 98.925 ;
        RECT 15.940 98.600 16.130 99.495 ;
        RECT 13.920 98.225 14.770 98.395 ;
        RECT 14.970 98.005 15.630 98.485 ;
        RECT 15.810 98.270 16.130 98.600 ;
        RECT 16.330 99.245 16.580 99.835 ;
        RECT 16.760 99.755 17.045 100.555 ;
        RECT 17.225 99.575 17.480 100.245 ;
        RECT 16.330 98.915 17.130 99.245 ;
        RECT 17.300 99.195 17.480 99.575 ;
        RECT 18.485 99.390 18.775 100.555 ;
        RECT 18.950 99.415 19.285 100.385 ;
        RECT 19.455 99.415 19.625 100.555 ;
        RECT 19.795 100.215 21.825 100.385 ;
        RECT 17.300 99.025 17.565 99.195 ;
        RECT 16.330 98.265 16.580 98.915 ;
        RECT 17.300 98.715 17.480 99.025 ;
        RECT 18.950 98.745 19.120 99.415 ;
        RECT 19.795 99.245 19.965 100.215 ;
        RECT 19.290 98.915 19.545 99.245 ;
        RECT 19.770 98.915 19.965 99.245 ;
        RECT 20.135 99.875 21.260 100.045 ;
        RECT 19.375 98.745 19.545 98.915 ;
        RECT 20.135 98.745 20.305 99.875 ;
        RECT 16.760 98.005 17.045 98.465 ;
        RECT 17.225 98.185 17.480 98.715 ;
        RECT 18.485 98.005 18.775 98.730 ;
        RECT 18.950 98.175 19.205 98.745 ;
        RECT 19.375 98.575 20.305 98.745 ;
        RECT 20.475 99.535 21.485 99.705 ;
        RECT 20.475 98.735 20.645 99.535 ;
        RECT 20.850 99.195 21.125 99.335 ;
        RECT 20.845 99.025 21.125 99.195 ;
        RECT 20.130 98.540 20.305 98.575 ;
        RECT 19.375 98.005 19.705 98.405 ;
        RECT 20.130 98.175 20.660 98.540 ;
        RECT 20.850 98.175 21.125 99.025 ;
        RECT 21.295 98.175 21.485 99.535 ;
        RECT 21.655 99.550 21.825 100.215 ;
        RECT 21.995 99.795 22.165 100.555 ;
        RECT 22.400 99.795 22.915 100.205 ;
        RECT 23.085 100.120 28.430 100.555 ;
        RECT 28.605 100.120 33.950 100.555 ;
        RECT 21.655 99.360 22.405 99.550 ;
        RECT 22.575 98.985 22.915 99.795 ;
        RECT 21.685 98.815 22.915 98.985 ;
        RECT 21.665 98.005 22.175 98.540 ;
        RECT 22.395 98.210 22.640 98.815 ;
        RECT 24.670 98.550 25.010 99.380 ;
        RECT 26.490 98.870 26.840 100.120 ;
        RECT 30.190 98.550 30.530 99.380 ;
        RECT 32.010 98.870 32.360 100.120 ;
        RECT 34.125 99.465 37.635 100.555 ;
        RECT 37.805 99.465 39.015 100.555 ;
        RECT 34.125 98.775 35.775 99.295 ;
        RECT 35.945 98.945 37.635 99.465 ;
        RECT 23.085 98.005 28.430 98.550 ;
        RECT 28.605 98.005 33.950 98.550 ;
        RECT 34.125 98.005 37.635 98.775 ;
        RECT 37.805 98.755 38.325 99.295 ;
        RECT 38.495 98.925 39.015 99.465 ;
        RECT 39.245 99.415 39.455 100.555 ;
        RECT 39.625 99.405 39.955 100.385 ;
        RECT 40.125 99.415 40.355 100.555 ;
        RECT 40.565 99.465 44.075 100.555 ;
        RECT 37.805 98.005 39.015 98.755 ;
        RECT 39.245 98.005 39.455 98.825 ;
        RECT 39.625 98.805 39.875 99.405 ;
        RECT 40.045 98.995 40.375 99.245 ;
        RECT 39.625 98.175 39.955 98.805 ;
        RECT 40.125 98.005 40.355 98.825 ;
        RECT 40.565 98.775 42.215 99.295 ;
        RECT 42.385 98.945 44.075 99.465 ;
        RECT 44.245 99.390 44.535 100.555 ;
        RECT 44.705 99.465 48.215 100.555 ;
        RECT 44.705 98.775 46.355 99.295 ;
        RECT 46.525 98.945 48.215 99.465 ;
        RECT 48.385 99.480 48.655 100.385 ;
        RECT 48.825 99.795 49.155 100.555 ;
        RECT 49.335 99.625 49.505 100.385 ;
        RECT 40.565 98.005 44.075 98.775 ;
        RECT 44.245 98.005 44.535 98.730 ;
        RECT 44.705 98.005 48.215 98.775 ;
        RECT 48.385 98.680 48.555 99.480 ;
        RECT 48.840 99.455 49.505 99.625 ;
        RECT 48.840 99.310 49.010 99.455 ;
        RECT 50.265 99.415 50.495 100.555 ;
        RECT 50.665 99.405 50.995 100.385 ;
        RECT 51.165 99.415 51.375 100.555 ;
        RECT 51.605 100.120 56.950 100.555 ;
        RECT 57.125 100.120 62.470 100.555 ;
        RECT 48.725 98.980 49.010 99.310 ;
        RECT 48.840 98.725 49.010 98.980 ;
        RECT 49.245 98.905 49.575 99.275 ;
        RECT 50.245 98.995 50.575 99.245 ;
        RECT 48.385 98.175 48.645 98.680 ;
        RECT 48.840 98.555 49.505 98.725 ;
        RECT 48.825 98.005 49.155 98.385 ;
        RECT 49.335 98.175 49.505 98.555 ;
        RECT 50.265 98.005 50.495 98.825 ;
        RECT 50.745 98.805 50.995 99.405 ;
        RECT 50.665 98.175 50.995 98.805 ;
        RECT 51.165 98.005 51.375 98.825 ;
        RECT 53.190 98.550 53.530 99.380 ;
        RECT 55.010 98.870 55.360 100.120 ;
        RECT 58.710 98.550 59.050 99.380 ;
        RECT 60.530 98.870 60.880 100.120 ;
        RECT 62.645 99.465 65.235 100.555 ;
        RECT 62.645 98.775 63.855 99.295 ;
        RECT 64.025 98.945 65.235 99.465 ;
        RECT 65.410 99.415 65.745 100.385 ;
        RECT 65.915 99.415 66.085 100.555 ;
        RECT 66.255 100.215 68.285 100.385 ;
        RECT 51.605 98.005 56.950 98.550 ;
        RECT 57.125 98.005 62.470 98.550 ;
        RECT 62.645 98.005 65.235 98.775 ;
        RECT 65.410 98.745 65.580 99.415 ;
        RECT 66.255 99.245 66.425 100.215 ;
        RECT 65.750 98.915 66.005 99.245 ;
        RECT 66.230 98.915 66.425 99.245 ;
        RECT 66.595 99.875 67.720 100.045 ;
        RECT 65.835 98.745 66.005 98.915 ;
        RECT 66.595 98.745 66.765 99.875 ;
        RECT 65.410 98.175 65.665 98.745 ;
        RECT 65.835 98.575 66.765 98.745 ;
        RECT 66.935 99.535 67.945 99.705 ;
        RECT 66.935 98.735 67.105 99.535 ;
        RECT 66.590 98.540 66.765 98.575 ;
        RECT 65.835 98.005 66.165 98.405 ;
        RECT 66.590 98.175 67.120 98.540 ;
        RECT 67.310 98.515 67.585 99.335 ;
        RECT 67.305 98.345 67.585 98.515 ;
        RECT 67.310 98.175 67.585 98.345 ;
        RECT 67.755 98.175 67.945 99.535 ;
        RECT 68.115 99.550 68.285 100.215 ;
        RECT 68.455 99.795 68.625 100.555 ;
        RECT 68.860 99.795 69.375 100.205 ;
        RECT 68.115 99.360 68.865 99.550 ;
        RECT 69.035 98.985 69.375 99.795 ;
        RECT 70.005 99.390 70.295 100.555 ;
        RECT 71.015 99.885 71.185 100.385 ;
        RECT 71.355 100.055 71.685 100.555 ;
        RECT 71.015 99.715 71.680 99.885 ;
        RECT 68.145 98.815 69.375 98.985 ;
        RECT 70.930 98.895 71.280 99.545 ;
        RECT 68.125 98.005 68.635 98.540 ;
        RECT 68.855 98.210 69.100 98.815 ;
        RECT 70.005 98.005 70.295 98.730 ;
        RECT 71.450 98.725 71.680 99.715 ;
        RECT 71.015 98.555 71.680 98.725 ;
        RECT 71.015 98.265 71.185 98.555 ;
        RECT 71.355 98.005 71.685 98.385 ;
        RECT 71.855 98.265 72.080 100.385 ;
        RECT 72.295 100.055 72.625 100.555 ;
        RECT 72.795 99.885 72.965 100.385 ;
        RECT 73.200 100.170 74.030 100.340 ;
        RECT 74.270 100.175 74.650 100.555 ;
        RECT 72.270 99.715 72.965 99.885 ;
        RECT 72.270 98.745 72.440 99.715 ;
        RECT 72.610 98.925 73.020 99.545 ;
        RECT 73.190 99.495 73.690 99.875 ;
        RECT 72.270 98.555 72.965 98.745 ;
        RECT 73.190 98.625 73.410 99.495 ;
        RECT 73.860 99.325 74.030 100.170 ;
        RECT 74.830 100.005 75.000 100.295 ;
        RECT 75.170 100.175 75.500 100.555 ;
        RECT 75.970 100.085 76.600 100.335 ;
        RECT 76.780 100.175 77.200 100.555 ;
        RECT 76.430 100.005 76.600 100.085 ;
        RECT 77.400 100.005 77.640 100.295 ;
        RECT 74.200 99.755 75.570 100.005 ;
        RECT 74.200 99.495 74.450 99.755 ;
        RECT 74.960 99.325 75.210 99.485 ;
        RECT 73.860 99.155 75.210 99.325 ;
        RECT 73.860 99.115 74.280 99.155 ;
        RECT 73.590 98.565 73.940 98.935 ;
        RECT 72.295 98.005 72.625 98.385 ;
        RECT 72.795 98.225 72.965 98.555 ;
        RECT 74.110 98.385 74.280 99.115 ;
        RECT 75.380 98.985 75.570 99.755 ;
        RECT 74.450 98.655 74.860 98.985 ;
        RECT 75.150 98.645 75.570 98.985 ;
        RECT 75.740 99.575 76.260 99.885 ;
        RECT 76.430 99.835 77.640 100.005 ;
        RECT 77.870 99.865 78.200 100.555 ;
        RECT 75.740 98.815 75.910 99.575 ;
        RECT 76.080 98.985 76.260 99.395 ;
        RECT 76.430 99.325 76.600 99.835 ;
        RECT 78.370 99.685 78.540 100.295 ;
        RECT 78.810 99.835 79.140 100.345 ;
        RECT 78.370 99.665 78.690 99.685 ;
        RECT 76.770 99.495 78.690 99.665 ;
        RECT 76.430 99.155 78.330 99.325 ;
        RECT 76.660 98.815 76.990 98.935 ;
        RECT 75.740 98.645 76.990 98.815 ;
        RECT 73.265 98.185 74.280 98.385 ;
        RECT 74.450 98.005 74.860 98.445 ;
        RECT 75.150 98.215 75.400 98.645 ;
        RECT 75.600 98.005 75.920 98.465 ;
        RECT 77.160 98.395 77.330 99.155 ;
        RECT 78.000 99.095 78.330 99.155 ;
        RECT 77.520 98.925 77.850 98.985 ;
        RECT 77.520 98.655 78.180 98.925 ;
        RECT 78.500 98.600 78.690 99.495 ;
        RECT 76.480 98.225 77.330 98.395 ;
        RECT 77.530 98.005 78.190 98.485 ;
        RECT 78.370 98.270 78.690 98.600 ;
        RECT 78.890 99.245 79.140 99.835 ;
        RECT 79.320 99.755 79.605 100.555 ;
        RECT 79.785 99.575 80.040 100.245 ;
        RECT 80.585 100.120 85.930 100.555 ;
        RECT 86.105 100.120 91.450 100.555 ;
        RECT 78.890 98.915 79.690 99.245 ;
        RECT 78.890 98.265 79.140 98.915 ;
        RECT 79.860 98.715 80.040 99.575 ;
        RECT 79.785 98.515 80.040 98.715 ;
        RECT 82.170 98.550 82.510 99.380 ;
        RECT 83.990 98.870 84.340 100.120 ;
        RECT 87.690 98.550 88.030 99.380 ;
        RECT 89.510 98.870 89.860 100.120 ;
        RECT 91.625 99.465 95.135 100.555 ;
        RECT 91.625 98.775 93.275 99.295 ;
        RECT 93.445 98.945 95.135 99.465 ;
        RECT 95.765 99.390 96.055 100.555 ;
        RECT 96.230 99.415 96.565 100.385 ;
        RECT 96.735 99.415 96.905 100.555 ;
        RECT 97.075 100.215 99.105 100.385 ;
        RECT 79.320 98.005 79.605 98.465 ;
        RECT 79.785 98.345 80.125 98.515 ;
        RECT 79.785 98.185 80.040 98.345 ;
        RECT 80.585 98.005 85.930 98.550 ;
        RECT 86.105 98.005 91.450 98.550 ;
        RECT 91.625 98.005 95.135 98.775 ;
        RECT 96.230 98.745 96.400 99.415 ;
        RECT 97.075 99.245 97.245 100.215 ;
        RECT 96.570 98.915 96.825 99.245 ;
        RECT 97.050 98.915 97.245 99.245 ;
        RECT 97.415 99.875 98.540 100.045 ;
        RECT 96.655 98.745 96.825 98.915 ;
        RECT 97.415 98.745 97.585 99.875 ;
        RECT 95.765 98.005 96.055 98.730 ;
        RECT 96.230 98.175 96.485 98.745 ;
        RECT 96.655 98.575 97.585 98.745 ;
        RECT 97.755 99.535 98.765 99.705 ;
        RECT 97.755 98.735 97.925 99.535 ;
        RECT 98.130 99.195 98.405 99.335 ;
        RECT 98.125 99.025 98.405 99.195 ;
        RECT 97.410 98.540 97.585 98.575 ;
        RECT 96.655 98.005 96.985 98.405 ;
        RECT 97.410 98.175 97.940 98.540 ;
        RECT 98.130 98.175 98.405 99.025 ;
        RECT 98.575 98.175 98.765 99.535 ;
        RECT 98.935 99.550 99.105 100.215 ;
        RECT 99.275 99.795 99.445 100.555 ;
        RECT 99.680 99.795 100.195 100.205 ;
        RECT 100.365 100.120 105.710 100.555 ;
        RECT 98.935 99.360 99.685 99.550 ;
        RECT 99.855 98.985 100.195 99.795 ;
        RECT 98.965 98.815 100.195 98.985 ;
        RECT 98.945 98.005 99.455 98.540 ;
        RECT 99.675 98.210 99.920 98.815 ;
        RECT 101.950 98.550 102.290 99.380 ;
        RECT 103.770 98.870 104.120 100.120 ;
        RECT 106.350 99.415 106.685 100.385 ;
        RECT 106.855 99.415 107.025 100.555 ;
        RECT 107.195 100.215 109.225 100.385 ;
        RECT 106.350 98.745 106.520 99.415 ;
        RECT 107.195 99.245 107.365 100.215 ;
        RECT 106.690 98.915 106.945 99.245 ;
        RECT 107.170 98.915 107.365 99.245 ;
        RECT 107.535 99.875 108.660 100.045 ;
        RECT 106.775 98.745 106.945 98.915 ;
        RECT 107.535 98.745 107.705 99.875 ;
        RECT 100.365 98.005 105.710 98.550 ;
        RECT 106.350 98.175 106.605 98.745 ;
        RECT 106.775 98.575 107.705 98.745 ;
        RECT 107.875 99.535 108.885 99.705 ;
        RECT 107.875 98.735 108.045 99.535 ;
        RECT 107.530 98.540 107.705 98.575 ;
        RECT 106.775 98.005 107.105 98.405 ;
        RECT 107.530 98.175 108.060 98.540 ;
        RECT 108.250 98.515 108.525 99.335 ;
        RECT 108.245 98.345 108.525 98.515 ;
        RECT 108.250 98.175 108.525 98.345 ;
        RECT 108.695 98.175 108.885 99.535 ;
        RECT 109.055 99.550 109.225 100.215 ;
        RECT 109.395 99.795 109.565 100.555 ;
        RECT 109.800 99.795 110.315 100.205 ;
        RECT 110.485 100.120 115.830 100.555 ;
        RECT 109.055 99.360 109.805 99.550 ;
        RECT 109.975 98.985 110.315 99.795 ;
        RECT 109.085 98.815 110.315 98.985 ;
        RECT 109.065 98.005 109.575 98.540 ;
        RECT 109.795 98.210 110.040 98.815 ;
        RECT 112.070 98.550 112.410 99.380 ;
        RECT 113.890 98.870 114.240 100.120 ;
        RECT 116.005 99.465 117.215 100.555 ;
        RECT 116.005 98.755 116.525 99.295 ;
        RECT 116.695 98.925 117.215 99.465 ;
        RECT 117.385 99.465 118.595 100.555 ;
        RECT 117.385 98.925 117.905 99.465 ;
        RECT 118.075 98.755 118.595 99.295 ;
        RECT 110.485 98.005 115.830 98.550 ;
        RECT 116.005 98.005 117.215 98.755 ;
        RECT 117.385 98.005 118.595 98.755 ;
        RECT 5.520 97.835 118.680 98.005 ;
        RECT 5.605 97.085 6.815 97.835 ;
        RECT 6.985 97.085 8.195 97.835 ;
        RECT 8.455 97.285 8.625 97.575 ;
        RECT 8.795 97.455 9.125 97.835 ;
        RECT 8.455 97.115 9.120 97.285 ;
        RECT 5.605 96.545 6.125 97.085 ;
        RECT 6.295 96.375 6.815 96.915 ;
        RECT 6.985 96.545 7.505 97.085 ;
        RECT 7.675 96.375 8.195 96.915 ;
        RECT 5.605 95.285 6.815 96.375 ;
        RECT 6.985 95.285 8.195 96.375 ;
        RECT 8.370 96.295 8.720 96.945 ;
        RECT 8.890 96.125 9.120 97.115 ;
        RECT 8.455 95.955 9.120 96.125 ;
        RECT 8.455 95.455 8.625 95.955 ;
        RECT 8.795 95.285 9.125 95.785 ;
        RECT 9.295 95.455 9.520 97.575 ;
        RECT 9.735 97.455 10.065 97.835 ;
        RECT 10.235 97.285 10.405 97.615 ;
        RECT 10.705 97.455 11.720 97.655 ;
        RECT 9.710 97.095 10.405 97.285 ;
        RECT 9.710 96.125 9.880 97.095 ;
        RECT 10.050 96.295 10.460 96.915 ;
        RECT 10.630 96.345 10.850 97.215 ;
        RECT 11.030 96.905 11.380 97.275 ;
        RECT 11.550 96.725 11.720 97.455 ;
        RECT 11.890 97.395 12.300 97.835 ;
        RECT 12.590 97.195 12.840 97.625 ;
        RECT 13.040 97.375 13.360 97.835 ;
        RECT 13.920 97.445 14.770 97.615 ;
        RECT 11.890 96.855 12.300 97.185 ;
        RECT 12.590 96.855 13.010 97.195 ;
        RECT 11.300 96.685 11.720 96.725 ;
        RECT 11.300 96.515 12.650 96.685 ;
        RECT 9.710 95.955 10.405 96.125 ;
        RECT 10.630 95.965 11.130 96.345 ;
        RECT 9.735 95.285 10.065 95.785 ;
        RECT 10.235 95.455 10.405 95.955 ;
        RECT 11.300 95.670 11.470 96.515 ;
        RECT 12.400 96.355 12.650 96.515 ;
        RECT 11.640 96.085 11.890 96.345 ;
        RECT 12.820 96.085 13.010 96.855 ;
        RECT 11.640 95.835 13.010 96.085 ;
        RECT 13.180 97.025 14.430 97.195 ;
        RECT 13.180 96.265 13.350 97.025 ;
        RECT 14.100 96.905 14.430 97.025 ;
        RECT 13.520 96.445 13.700 96.855 ;
        RECT 14.600 96.685 14.770 97.445 ;
        RECT 14.970 97.355 15.630 97.835 ;
        RECT 15.810 97.240 16.130 97.570 ;
        RECT 14.960 96.915 15.620 97.185 ;
        RECT 14.960 96.855 15.290 96.915 ;
        RECT 15.440 96.685 15.770 96.745 ;
        RECT 13.870 96.515 15.770 96.685 ;
        RECT 13.180 95.955 13.700 96.265 ;
        RECT 13.870 96.005 14.040 96.515 ;
        RECT 15.940 96.345 16.130 97.240 ;
        RECT 14.210 96.175 16.130 96.345 ;
        RECT 15.810 96.155 16.130 96.175 ;
        RECT 16.330 96.925 16.580 97.575 ;
        RECT 16.760 97.375 17.045 97.835 ;
        RECT 17.225 97.495 17.480 97.655 ;
        RECT 17.225 97.325 17.565 97.495 ;
        RECT 17.225 97.125 17.480 97.325 ;
        RECT 16.330 96.595 17.130 96.925 ;
        RECT 13.870 95.835 15.080 96.005 ;
        RECT 10.640 95.500 11.470 95.670 ;
        RECT 11.710 95.285 12.090 95.665 ;
        RECT 12.270 95.545 12.440 95.835 ;
        RECT 13.870 95.755 14.040 95.835 ;
        RECT 12.610 95.285 12.940 95.665 ;
        RECT 13.410 95.505 14.040 95.755 ;
        RECT 14.220 95.285 14.640 95.665 ;
        RECT 14.840 95.545 15.080 95.835 ;
        RECT 15.310 95.285 15.640 95.975 ;
        RECT 15.810 95.545 15.980 96.155 ;
        RECT 16.330 96.005 16.580 96.595 ;
        RECT 17.300 96.265 17.480 97.125 ;
        RECT 16.250 95.495 16.580 96.005 ;
        RECT 16.760 95.285 17.045 96.085 ;
        RECT 17.225 95.595 17.480 96.265 ;
        RECT 18.030 97.095 18.285 97.665 ;
        RECT 18.455 97.435 18.785 97.835 ;
        RECT 19.210 97.300 19.740 97.665 ;
        RECT 19.930 97.495 20.205 97.665 ;
        RECT 19.925 97.325 20.205 97.495 ;
        RECT 19.210 97.265 19.385 97.300 ;
        RECT 18.455 97.095 19.385 97.265 ;
        RECT 18.030 96.425 18.200 97.095 ;
        RECT 18.455 96.925 18.625 97.095 ;
        RECT 18.370 96.595 18.625 96.925 ;
        RECT 18.850 96.595 19.045 96.925 ;
        RECT 18.030 95.455 18.365 96.425 ;
        RECT 18.535 95.285 18.705 96.425 ;
        RECT 18.875 95.625 19.045 96.595 ;
        RECT 19.215 95.965 19.385 97.095 ;
        RECT 19.555 96.305 19.725 97.105 ;
        RECT 19.930 96.505 20.205 97.325 ;
        RECT 20.375 96.305 20.565 97.665 ;
        RECT 20.745 97.300 21.255 97.835 ;
        RECT 21.475 97.025 21.720 97.630 ;
        RECT 22.165 97.290 27.510 97.835 ;
        RECT 20.765 96.855 21.995 97.025 ;
        RECT 19.555 96.135 20.565 96.305 ;
        RECT 20.735 96.290 21.485 96.480 ;
        RECT 19.215 95.795 20.340 95.965 ;
        RECT 20.735 95.625 20.905 96.290 ;
        RECT 21.655 96.045 21.995 96.855 ;
        RECT 23.750 96.460 24.090 97.290 ;
        RECT 27.685 97.065 31.195 97.835 ;
        RECT 31.365 97.110 31.655 97.835 ;
        RECT 31.825 97.375 32.385 97.665 ;
        RECT 32.555 97.375 32.805 97.835 ;
        RECT 18.875 95.455 20.905 95.625 ;
        RECT 21.075 95.285 21.245 96.045 ;
        RECT 21.480 95.635 21.995 96.045 ;
        RECT 25.570 95.720 25.920 96.970 ;
        RECT 27.685 96.545 29.335 97.065 ;
        RECT 29.505 96.375 31.195 96.895 ;
        RECT 22.165 95.285 27.510 95.720 ;
        RECT 27.685 95.285 31.195 96.375 ;
        RECT 31.365 95.285 31.655 96.450 ;
        RECT 31.825 96.005 32.075 97.375 ;
        RECT 33.425 97.205 33.755 97.565 ;
        RECT 32.365 97.015 33.755 97.205 ;
        RECT 34.500 97.125 34.755 97.655 ;
        RECT 34.935 97.375 35.220 97.835 ;
        RECT 32.365 96.925 32.535 97.015 ;
        RECT 32.245 96.595 32.535 96.925 ;
        RECT 32.705 96.595 33.045 96.845 ;
        RECT 33.265 96.595 33.940 96.845 ;
        RECT 32.365 96.345 32.535 96.595 ;
        RECT 32.365 96.175 33.305 96.345 ;
        RECT 33.675 96.235 33.940 96.595 ;
        RECT 34.500 96.265 34.680 97.125 ;
        RECT 35.400 96.925 35.650 97.575 ;
        RECT 34.850 96.595 35.650 96.925 ;
        RECT 31.825 95.455 32.285 96.005 ;
        RECT 32.475 95.285 32.805 96.005 ;
        RECT 33.005 95.625 33.305 96.175 ;
        RECT 33.475 95.285 33.755 95.955 ;
        RECT 34.500 95.795 34.755 96.265 ;
        RECT 34.415 95.625 34.755 95.795 ;
        RECT 34.500 95.595 34.755 95.625 ;
        RECT 34.935 95.285 35.220 96.085 ;
        RECT 35.400 96.005 35.650 96.595 ;
        RECT 35.850 97.240 36.170 97.570 ;
        RECT 36.350 97.355 37.010 97.835 ;
        RECT 37.210 97.445 38.060 97.615 ;
        RECT 35.850 96.345 36.040 97.240 ;
        RECT 36.360 96.915 37.020 97.185 ;
        RECT 36.690 96.855 37.020 96.915 ;
        RECT 36.210 96.685 36.540 96.745 ;
        RECT 37.210 96.685 37.380 97.445 ;
        RECT 38.620 97.375 38.940 97.835 ;
        RECT 39.140 97.195 39.390 97.625 ;
        RECT 39.680 97.395 40.090 97.835 ;
        RECT 40.260 97.455 41.275 97.655 ;
        RECT 37.550 97.025 38.800 97.195 ;
        RECT 37.550 96.905 37.880 97.025 ;
        RECT 36.210 96.515 38.110 96.685 ;
        RECT 35.850 96.175 37.770 96.345 ;
        RECT 35.850 96.155 36.170 96.175 ;
        RECT 35.400 95.495 35.730 96.005 ;
        RECT 36.000 95.545 36.170 96.155 ;
        RECT 37.940 96.005 38.110 96.515 ;
        RECT 38.280 96.445 38.460 96.855 ;
        RECT 38.630 96.265 38.800 97.025 ;
        RECT 36.340 95.285 36.670 95.975 ;
        RECT 36.900 95.835 38.110 96.005 ;
        RECT 38.280 95.955 38.800 96.265 ;
        RECT 38.970 96.855 39.390 97.195 ;
        RECT 39.680 96.855 40.090 97.185 ;
        RECT 38.970 96.085 39.160 96.855 ;
        RECT 40.260 96.725 40.430 97.455 ;
        RECT 41.575 97.285 41.745 97.615 ;
        RECT 41.915 97.455 42.245 97.835 ;
        RECT 40.600 96.905 40.950 97.275 ;
        RECT 40.260 96.685 40.680 96.725 ;
        RECT 39.330 96.515 40.680 96.685 ;
        RECT 39.330 96.355 39.580 96.515 ;
        RECT 40.090 96.085 40.340 96.345 ;
        RECT 38.970 95.835 40.340 96.085 ;
        RECT 36.900 95.545 37.140 95.835 ;
        RECT 37.940 95.755 38.110 95.835 ;
        RECT 37.340 95.285 37.760 95.665 ;
        RECT 37.940 95.505 38.570 95.755 ;
        RECT 39.040 95.285 39.370 95.665 ;
        RECT 39.540 95.545 39.710 95.835 ;
        RECT 40.510 95.670 40.680 96.515 ;
        RECT 41.130 96.345 41.350 97.215 ;
        RECT 41.575 97.095 42.270 97.285 ;
        RECT 40.850 95.965 41.350 96.345 ;
        RECT 41.520 96.295 41.930 96.915 ;
        RECT 42.100 96.125 42.270 97.095 ;
        RECT 41.575 95.955 42.270 96.125 ;
        RECT 39.890 95.285 40.270 95.665 ;
        RECT 40.510 95.500 41.340 95.670 ;
        RECT 41.575 95.455 41.745 95.955 ;
        RECT 41.915 95.285 42.245 95.785 ;
        RECT 42.460 95.455 42.685 97.575 ;
        RECT 42.855 97.455 43.185 97.835 ;
        RECT 43.355 97.285 43.525 97.575 ;
        RECT 42.860 97.115 43.525 97.285 ;
        RECT 42.860 96.125 43.090 97.115 ;
        RECT 43.785 97.065 45.455 97.835 ;
        RECT 45.715 97.285 45.885 97.575 ;
        RECT 46.055 97.455 46.385 97.835 ;
        RECT 45.715 97.115 46.380 97.285 ;
        RECT 43.260 96.295 43.610 96.945 ;
        RECT 43.785 96.545 44.535 97.065 ;
        RECT 44.705 96.375 45.455 96.895 ;
        RECT 42.860 95.955 43.525 96.125 ;
        RECT 42.855 95.285 43.185 95.785 ;
        RECT 43.355 95.455 43.525 95.955 ;
        RECT 43.785 95.285 45.455 96.375 ;
        RECT 45.630 96.295 45.980 96.945 ;
        RECT 46.150 96.125 46.380 97.115 ;
        RECT 45.715 95.955 46.380 96.125 ;
        RECT 45.715 95.455 45.885 95.955 ;
        RECT 46.055 95.285 46.385 95.785 ;
        RECT 46.555 95.455 46.780 97.575 ;
        RECT 46.995 97.455 47.325 97.835 ;
        RECT 47.495 97.285 47.665 97.615 ;
        RECT 47.965 97.455 48.980 97.655 ;
        RECT 46.970 97.095 47.665 97.285 ;
        RECT 46.970 96.125 47.140 97.095 ;
        RECT 47.310 96.295 47.720 96.915 ;
        RECT 47.890 96.345 48.110 97.215 ;
        RECT 48.290 96.905 48.640 97.275 ;
        RECT 48.810 96.725 48.980 97.455 ;
        RECT 49.150 97.395 49.560 97.835 ;
        RECT 49.850 97.195 50.100 97.625 ;
        RECT 50.300 97.375 50.620 97.835 ;
        RECT 51.180 97.445 52.030 97.615 ;
        RECT 49.150 96.855 49.560 97.185 ;
        RECT 49.850 96.855 50.270 97.195 ;
        RECT 48.560 96.685 48.980 96.725 ;
        RECT 48.560 96.515 49.910 96.685 ;
        RECT 46.970 95.955 47.665 96.125 ;
        RECT 47.890 95.965 48.390 96.345 ;
        RECT 46.995 95.285 47.325 95.785 ;
        RECT 47.495 95.455 47.665 95.955 ;
        RECT 48.560 95.670 48.730 96.515 ;
        RECT 49.660 96.355 49.910 96.515 ;
        RECT 48.900 96.085 49.150 96.345 ;
        RECT 50.080 96.085 50.270 96.855 ;
        RECT 48.900 95.835 50.270 96.085 ;
        RECT 50.440 97.025 51.690 97.195 ;
        RECT 50.440 96.265 50.610 97.025 ;
        RECT 51.360 96.905 51.690 97.025 ;
        RECT 50.780 96.445 50.960 96.855 ;
        RECT 51.860 96.685 52.030 97.445 ;
        RECT 52.230 97.355 52.890 97.835 ;
        RECT 53.070 97.240 53.390 97.570 ;
        RECT 52.220 96.915 52.880 97.185 ;
        RECT 52.220 96.855 52.550 96.915 ;
        RECT 52.700 96.685 53.030 96.745 ;
        RECT 51.130 96.515 53.030 96.685 ;
        RECT 50.440 95.955 50.960 96.265 ;
        RECT 51.130 96.005 51.300 96.515 ;
        RECT 53.200 96.345 53.390 97.240 ;
        RECT 51.470 96.175 53.390 96.345 ;
        RECT 53.070 96.155 53.390 96.175 ;
        RECT 53.590 96.925 53.840 97.575 ;
        RECT 54.020 97.375 54.305 97.835 ;
        RECT 54.485 97.125 54.740 97.655 ;
        RECT 53.590 96.595 54.390 96.925 ;
        RECT 51.130 95.835 52.340 96.005 ;
        RECT 47.900 95.500 48.730 95.670 ;
        RECT 48.970 95.285 49.350 95.665 ;
        RECT 49.530 95.545 49.700 95.835 ;
        RECT 51.130 95.755 51.300 95.835 ;
        RECT 49.870 95.285 50.200 95.665 ;
        RECT 50.670 95.505 51.300 95.755 ;
        RECT 51.480 95.285 51.900 95.665 ;
        RECT 52.100 95.545 52.340 95.835 ;
        RECT 52.570 95.285 52.900 95.975 ;
        RECT 53.070 95.545 53.240 96.155 ;
        RECT 53.590 96.005 53.840 96.595 ;
        RECT 54.560 96.265 54.740 97.125 ;
        RECT 55.285 97.065 56.955 97.835 ;
        RECT 57.125 97.110 57.415 97.835 ;
        RECT 58.105 97.355 58.385 97.835 ;
        RECT 58.555 97.185 58.815 97.575 ;
        RECT 58.990 97.355 59.245 97.835 ;
        RECT 59.415 97.185 59.710 97.575 ;
        RECT 59.890 97.355 60.165 97.835 ;
        RECT 60.335 97.335 60.635 97.665 ;
        RECT 55.285 96.545 56.035 97.065 ;
        RECT 58.060 97.015 59.710 97.185 ;
        RECT 56.205 96.375 56.955 96.895 ;
        RECT 58.060 96.505 58.465 97.015 ;
        RECT 58.635 96.675 59.775 96.845 ;
        RECT 53.510 95.495 53.840 96.005 ;
        RECT 54.020 95.285 54.305 96.085 ;
        RECT 54.485 95.795 54.740 96.265 ;
        RECT 54.485 95.625 54.825 95.795 ;
        RECT 54.485 95.595 54.740 95.625 ;
        RECT 55.285 95.285 56.955 96.375 ;
        RECT 57.125 95.285 57.415 96.450 ;
        RECT 58.060 96.335 58.815 96.505 ;
        RECT 58.100 95.285 58.385 96.155 ;
        RECT 58.555 96.085 58.815 96.335 ;
        RECT 59.605 96.425 59.775 96.675 ;
        RECT 59.945 96.595 60.295 97.165 ;
        RECT 60.465 96.425 60.635 97.335 ;
        RECT 59.605 96.255 60.635 96.425 ;
        RECT 58.555 95.915 59.675 96.085 ;
        RECT 58.555 95.455 58.815 95.915 ;
        RECT 58.990 95.285 59.245 95.745 ;
        RECT 59.415 95.455 59.675 95.915 ;
        RECT 59.845 95.285 60.155 96.085 ;
        RECT 60.325 95.455 60.635 96.255 ;
        RECT 61.725 97.160 61.985 97.665 ;
        RECT 62.165 97.455 62.495 97.835 ;
        RECT 62.675 97.285 62.845 97.665 ;
        RECT 61.725 96.360 61.895 97.160 ;
        RECT 62.180 97.115 62.845 97.285 ;
        RECT 62.180 96.860 62.350 97.115 ;
        RECT 63.605 97.015 63.835 97.835 ;
        RECT 64.005 97.035 64.335 97.665 ;
        RECT 62.065 96.530 62.350 96.860 ;
        RECT 62.585 96.565 62.915 96.935 ;
        RECT 63.585 96.595 63.915 96.845 ;
        RECT 62.180 96.385 62.350 96.530 ;
        RECT 64.085 96.435 64.335 97.035 ;
        RECT 64.505 97.015 64.715 97.835 ;
        RECT 64.945 97.065 68.455 97.835 ;
        RECT 68.625 97.085 69.835 97.835 ;
        RECT 70.010 97.095 70.265 97.665 ;
        RECT 70.435 97.435 70.765 97.835 ;
        RECT 71.190 97.300 71.720 97.665 ;
        RECT 71.190 97.265 71.365 97.300 ;
        RECT 70.435 97.095 71.365 97.265 ;
        RECT 64.945 96.545 66.595 97.065 ;
        RECT 61.725 95.455 61.995 96.360 ;
        RECT 62.180 96.215 62.845 96.385 ;
        RECT 62.165 95.285 62.495 96.045 ;
        RECT 62.675 95.455 62.845 96.215 ;
        RECT 63.605 95.285 63.835 96.425 ;
        RECT 64.005 95.455 64.335 96.435 ;
        RECT 64.505 95.285 64.715 96.425 ;
        RECT 66.765 96.375 68.455 96.895 ;
        RECT 68.625 96.545 69.145 97.085 ;
        RECT 69.315 96.375 69.835 96.915 ;
        RECT 64.945 95.285 68.455 96.375 ;
        RECT 68.625 95.285 69.835 96.375 ;
        RECT 70.010 96.425 70.180 97.095 ;
        RECT 70.435 96.925 70.605 97.095 ;
        RECT 70.350 96.595 70.605 96.925 ;
        RECT 70.830 96.595 71.025 96.925 ;
        RECT 70.010 95.455 70.345 96.425 ;
        RECT 70.515 95.285 70.685 96.425 ;
        RECT 70.855 95.625 71.025 96.595 ;
        RECT 71.195 95.965 71.365 97.095 ;
        RECT 71.535 96.305 71.705 97.105 ;
        RECT 71.910 96.815 72.185 97.665 ;
        RECT 71.905 96.645 72.185 96.815 ;
        RECT 71.910 96.505 72.185 96.645 ;
        RECT 72.355 96.305 72.545 97.665 ;
        RECT 72.725 97.300 73.235 97.835 ;
        RECT 73.455 97.025 73.700 97.630 ;
        RECT 74.145 97.160 74.405 97.665 ;
        RECT 74.585 97.455 74.915 97.835 ;
        RECT 75.095 97.285 75.265 97.665 ;
        RECT 75.525 97.290 80.870 97.835 ;
        RECT 72.745 96.855 73.975 97.025 ;
        RECT 71.535 96.135 72.545 96.305 ;
        RECT 72.715 96.290 73.465 96.480 ;
        RECT 71.195 95.795 72.320 95.965 ;
        RECT 72.715 95.625 72.885 96.290 ;
        RECT 73.635 96.045 73.975 96.855 ;
        RECT 70.855 95.455 72.885 95.625 ;
        RECT 73.055 95.285 73.225 96.045 ;
        RECT 73.460 95.635 73.975 96.045 ;
        RECT 74.145 96.360 74.315 97.160 ;
        RECT 74.600 97.115 75.265 97.285 ;
        RECT 74.600 96.860 74.770 97.115 ;
        RECT 74.485 96.530 74.770 96.860 ;
        RECT 75.005 96.565 75.335 96.935 ;
        RECT 74.600 96.385 74.770 96.530 ;
        RECT 77.110 96.460 77.450 97.290 ;
        RECT 81.045 97.065 82.715 97.835 ;
        RECT 82.885 97.110 83.175 97.835 ;
        RECT 83.345 97.335 83.645 97.665 ;
        RECT 83.815 97.355 84.090 97.835 ;
        RECT 74.145 95.455 74.415 96.360 ;
        RECT 74.600 96.215 75.265 96.385 ;
        RECT 74.585 95.285 74.915 96.045 ;
        RECT 75.095 95.455 75.265 96.215 ;
        RECT 78.930 95.720 79.280 96.970 ;
        RECT 81.045 96.545 81.795 97.065 ;
        RECT 81.965 96.375 82.715 96.895 ;
        RECT 75.525 95.285 80.870 95.720 ;
        RECT 81.045 95.285 82.715 96.375 ;
        RECT 82.885 95.285 83.175 96.450 ;
        RECT 83.345 96.425 83.515 97.335 ;
        RECT 84.270 97.185 84.565 97.575 ;
        RECT 84.735 97.355 84.990 97.835 ;
        RECT 85.165 97.185 85.425 97.575 ;
        RECT 85.595 97.355 85.875 97.835 ;
        RECT 86.305 97.205 86.635 97.565 ;
        RECT 87.255 97.375 87.505 97.835 ;
        RECT 87.675 97.375 88.235 97.665 ;
        RECT 83.685 96.595 84.035 97.165 ;
        RECT 84.270 97.015 85.920 97.185 ;
        RECT 86.305 97.015 87.695 97.205 ;
        RECT 84.205 96.675 85.345 96.845 ;
        RECT 84.205 96.425 84.375 96.675 ;
        RECT 85.515 96.505 85.920 97.015 ;
        RECT 87.525 96.925 87.695 97.015 ;
        RECT 83.345 96.255 84.375 96.425 ;
        RECT 85.165 96.335 85.920 96.505 ;
        RECT 86.120 96.595 86.795 96.845 ;
        RECT 87.015 96.595 87.355 96.845 ;
        RECT 87.525 96.595 87.815 96.925 ;
        RECT 83.345 95.455 83.655 96.255 ;
        RECT 85.165 96.085 85.425 96.335 ;
        RECT 86.120 96.235 86.385 96.595 ;
        RECT 87.525 96.345 87.695 96.595 ;
        RECT 86.755 96.175 87.695 96.345 ;
        RECT 83.825 95.285 84.135 96.085 ;
        RECT 84.305 95.915 85.425 96.085 ;
        RECT 84.305 95.455 84.565 95.915 ;
        RECT 84.735 95.285 84.990 95.745 ;
        RECT 85.165 95.455 85.425 95.915 ;
        RECT 85.595 95.285 85.880 96.155 ;
        RECT 86.305 95.285 86.585 95.955 ;
        RECT 86.755 95.625 87.055 96.175 ;
        RECT 87.985 96.005 88.235 97.375 ;
        RECT 87.255 95.285 87.585 96.005 ;
        RECT 87.775 95.455 88.235 96.005 ;
        RECT 88.405 97.375 88.965 97.665 ;
        RECT 89.135 97.375 89.385 97.835 ;
        RECT 88.405 96.005 88.655 97.375 ;
        RECT 90.005 97.205 90.335 97.565 ;
        RECT 88.945 97.015 90.335 97.205 ;
        RECT 90.905 97.205 91.235 97.565 ;
        RECT 91.855 97.375 92.105 97.835 ;
        RECT 92.275 97.375 92.835 97.665 ;
        RECT 90.905 97.015 92.295 97.205 ;
        RECT 88.945 96.925 89.115 97.015 ;
        RECT 88.825 96.595 89.115 96.925 ;
        RECT 92.125 96.925 92.295 97.015 ;
        RECT 89.285 96.595 89.625 96.845 ;
        RECT 89.845 96.595 90.520 96.845 ;
        RECT 88.945 96.345 89.115 96.595 ;
        RECT 88.945 96.175 89.885 96.345 ;
        RECT 90.255 96.235 90.520 96.595 ;
        RECT 90.720 96.595 91.395 96.845 ;
        RECT 91.615 96.595 91.955 96.845 ;
        RECT 92.125 96.595 92.415 96.925 ;
        RECT 90.720 96.235 90.985 96.595 ;
        RECT 92.125 96.345 92.295 96.595 ;
        RECT 88.405 95.455 88.865 96.005 ;
        RECT 89.055 95.285 89.385 96.005 ;
        RECT 89.585 95.625 89.885 96.175 ;
        RECT 91.355 96.175 92.295 96.345 ;
        RECT 90.055 95.285 90.335 95.955 ;
        RECT 90.905 95.285 91.185 95.955 ;
        RECT 91.355 95.625 91.655 96.175 ;
        RECT 92.585 96.005 92.835 97.375 ;
        RECT 93.005 97.085 94.215 97.835 ;
        RECT 94.385 97.375 94.945 97.665 ;
        RECT 95.115 97.375 95.365 97.835 ;
        RECT 93.005 96.545 93.525 97.085 ;
        RECT 93.695 96.375 94.215 96.915 ;
        RECT 91.855 95.285 92.185 96.005 ;
        RECT 92.375 95.455 92.835 96.005 ;
        RECT 93.005 95.285 94.215 96.375 ;
        RECT 94.385 96.005 94.635 97.375 ;
        RECT 95.985 97.205 96.315 97.565 ;
        RECT 96.685 97.290 102.030 97.835 ;
        RECT 102.205 97.290 107.550 97.835 ;
        RECT 94.925 97.015 96.315 97.205 ;
        RECT 94.925 96.925 95.095 97.015 ;
        RECT 94.805 96.595 95.095 96.925 ;
        RECT 95.265 96.595 95.605 96.845 ;
        RECT 95.825 96.595 96.500 96.845 ;
        RECT 94.925 96.345 95.095 96.595 ;
        RECT 94.925 96.175 95.865 96.345 ;
        RECT 96.235 96.235 96.500 96.595 ;
        RECT 98.270 96.460 98.610 97.290 ;
        RECT 94.385 95.455 94.845 96.005 ;
        RECT 95.035 95.285 95.365 96.005 ;
        RECT 95.565 95.625 95.865 96.175 ;
        RECT 96.035 95.285 96.315 95.955 ;
        RECT 100.090 95.720 100.440 96.970 ;
        RECT 103.790 96.460 104.130 97.290 ;
        RECT 108.645 97.110 108.935 97.835 ;
        RECT 109.105 97.160 109.365 97.665 ;
        RECT 109.545 97.455 109.875 97.835 ;
        RECT 110.055 97.285 110.225 97.665 ;
        RECT 105.610 95.720 105.960 96.970 ;
        RECT 96.685 95.285 102.030 95.720 ;
        RECT 102.205 95.285 107.550 95.720 ;
        RECT 108.645 95.285 108.935 96.450 ;
        RECT 109.105 96.360 109.275 97.160 ;
        RECT 109.560 97.115 110.225 97.285 ;
        RECT 109.560 96.860 109.730 97.115 ;
        RECT 110.985 97.015 111.215 97.835 ;
        RECT 111.385 97.035 111.715 97.665 ;
        RECT 109.445 96.530 109.730 96.860 ;
        RECT 109.965 96.565 110.295 96.935 ;
        RECT 110.965 96.595 111.295 96.845 ;
        RECT 109.560 96.385 109.730 96.530 ;
        RECT 111.465 96.435 111.715 97.035 ;
        RECT 111.885 97.015 112.095 97.835 ;
        RECT 112.325 97.065 115.835 97.835 ;
        RECT 116.005 97.085 117.215 97.835 ;
        RECT 117.385 97.085 118.595 97.835 ;
        RECT 112.325 96.545 113.975 97.065 ;
        RECT 109.105 95.455 109.375 96.360 ;
        RECT 109.560 96.215 110.225 96.385 ;
        RECT 109.545 95.285 109.875 96.045 ;
        RECT 110.055 95.455 110.225 96.215 ;
        RECT 110.985 95.285 111.215 96.425 ;
        RECT 111.385 95.455 111.715 96.435 ;
        RECT 111.885 95.285 112.095 96.425 ;
        RECT 114.145 96.375 115.835 96.895 ;
        RECT 116.005 96.545 116.525 97.085 ;
        RECT 116.695 96.375 117.215 96.915 ;
        RECT 112.325 95.285 115.835 96.375 ;
        RECT 116.005 95.285 117.215 96.375 ;
        RECT 117.385 96.375 117.905 96.915 ;
        RECT 118.075 96.545 118.595 97.085 ;
        RECT 117.385 95.285 118.595 96.375 ;
        RECT 5.520 95.115 118.680 95.285 ;
        RECT 5.605 94.025 6.815 95.115 ;
        RECT 6.985 94.680 12.330 95.115 ;
        RECT 5.605 93.315 6.125 93.855 ;
        RECT 6.295 93.485 6.815 94.025 ;
        RECT 5.605 92.565 6.815 93.315 ;
        RECT 8.570 93.110 8.910 93.940 ;
        RECT 10.390 93.430 10.740 94.680 ;
        RECT 12.505 94.040 12.775 94.945 ;
        RECT 12.945 94.355 13.275 95.115 ;
        RECT 13.455 94.185 13.625 94.945 ;
        RECT 12.505 93.240 12.675 94.040 ;
        RECT 12.960 94.015 13.625 94.185 ;
        RECT 12.960 93.870 13.130 94.015 ;
        RECT 13.945 93.975 14.155 95.115 ;
        RECT 12.845 93.540 13.130 93.870 ;
        RECT 14.325 93.965 14.655 94.945 ;
        RECT 14.825 93.975 15.055 95.115 ;
        RECT 15.265 94.025 17.855 95.115 ;
        RECT 12.960 93.285 13.130 93.540 ;
        RECT 13.365 93.465 13.695 93.835 ;
        RECT 6.985 92.565 12.330 93.110 ;
        RECT 12.505 92.735 12.765 93.240 ;
        RECT 12.960 93.115 13.625 93.285 ;
        RECT 12.945 92.565 13.275 92.945 ;
        RECT 13.455 92.735 13.625 93.115 ;
        RECT 13.945 92.565 14.155 93.385 ;
        RECT 14.325 93.365 14.575 93.965 ;
        RECT 14.745 93.555 15.075 93.805 ;
        RECT 14.325 92.735 14.655 93.365 ;
        RECT 14.825 92.565 15.055 93.385 ;
        RECT 15.265 93.335 16.475 93.855 ;
        RECT 16.645 93.505 17.855 94.025 ;
        RECT 18.485 93.950 18.775 95.115 ;
        RECT 19.605 94.445 19.885 95.115 ;
        RECT 20.055 94.225 20.355 94.775 ;
        RECT 20.555 94.395 20.885 95.115 ;
        RECT 21.075 94.395 21.535 94.945 ;
        RECT 19.420 93.805 19.685 94.165 ;
        RECT 20.055 94.055 20.995 94.225 ;
        RECT 20.825 93.805 20.995 94.055 ;
        RECT 19.420 93.555 20.095 93.805 ;
        RECT 20.315 93.555 20.655 93.805 ;
        RECT 20.825 93.475 21.115 93.805 ;
        RECT 20.825 93.385 20.995 93.475 ;
        RECT 15.265 92.565 17.855 93.335 ;
        RECT 18.485 92.565 18.775 93.290 ;
        RECT 19.605 93.195 20.995 93.385 ;
        RECT 19.605 92.835 19.935 93.195 ;
        RECT 21.285 93.025 21.535 94.395 ;
        RECT 20.555 92.565 20.805 93.025 ;
        RECT 20.975 92.735 21.535 93.025 ;
        RECT 21.705 94.395 22.165 94.945 ;
        RECT 22.355 94.395 22.685 95.115 ;
        RECT 21.705 93.025 21.955 94.395 ;
        RECT 22.885 94.225 23.185 94.775 ;
        RECT 23.355 94.445 23.635 95.115 ;
        RECT 24.205 94.445 24.485 95.115 ;
        RECT 22.245 94.055 23.185 94.225 ;
        RECT 24.655 94.225 24.955 94.775 ;
        RECT 25.155 94.395 25.485 95.115 ;
        RECT 25.675 94.395 26.135 94.945 ;
        RECT 26.505 94.445 26.785 95.115 ;
        RECT 22.245 93.805 22.415 94.055 ;
        RECT 23.555 93.805 23.820 94.165 ;
        RECT 22.125 93.475 22.415 93.805 ;
        RECT 22.585 93.555 22.925 93.805 ;
        RECT 23.145 93.555 23.820 93.805 ;
        RECT 24.020 93.805 24.285 94.165 ;
        RECT 24.655 94.055 25.595 94.225 ;
        RECT 25.425 93.805 25.595 94.055 ;
        RECT 24.020 93.555 24.695 93.805 ;
        RECT 24.915 93.555 25.255 93.805 ;
        RECT 22.245 93.385 22.415 93.475 ;
        RECT 25.425 93.475 25.715 93.805 ;
        RECT 25.425 93.385 25.595 93.475 ;
        RECT 22.245 93.195 23.635 93.385 ;
        RECT 21.705 92.735 22.265 93.025 ;
        RECT 22.435 92.565 22.685 93.025 ;
        RECT 23.305 92.835 23.635 93.195 ;
        RECT 24.205 93.195 25.595 93.385 ;
        RECT 24.205 92.835 24.535 93.195 ;
        RECT 25.885 93.025 26.135 94.395 ;
        RECT 26.955 94.225 27.255 94.775 ;
        RECT 27.455 94.395 27.785 95.115 ;
        RECT 27.975 94.395 28.435 94.945 ;
        RECT 26.320 93.805 26.585 94.165 ;
        RECT 26.955 94.055 27.895 94.225 ;
        RECT 27.725 93.805 27.895 94.055 ;
        RECT 26.320 93.555 26.995 93.805 ;
        RECT 27.215 93.555 27.555 93.805 ;
        RECT 27.725 93.475 28.015 93.805 ;
        RECT 27.725 93.385 27.895 93.475 ;
        RECT 25.155 92.565 25.405 93.025 ;
        RECT 25.575 92.735 26.135 93.025 ;
        RECT 26.505 93.195 27.895 93.385 ;
        RECT 26.505 92.835 26.835 93.195 ;
        RECT 28.185 93.025 28.435 94.395 ;
        RECT 28.695 94.370 28.965 95.115 ;
        RECT 29.595 95.110 35.870 95.115 ;
        RECT 29.135 94.200 29.425 94.940 ;
        RECT 29.595 94.385 29.850 95.110 ;
        RECT 30.035 94.215 30.295 94.940 ;
        RECT 30.465 94.385 30.710 95.110 ;
        RECT 30.895 94.215 31.155 94.940 ;
        RECT 31.325 94.385 31.570 95.110 ;
        RECT 31.755 94.215 32.015 94.940 ;
        RECT 32.185 94.385 32.430 95.110 ;
        RECT 32.600 94.215 32.860 94.940 ;
        RECT 33.030 94.385 33.290 95.110 ;
        RECT 33.460 94.215 33.720 94.940 ;
        RECT 33.890 94.385 34.150 95.110 ;
        RECT 34.320 94.215 34.580 94.940 ;
        RECT 34.750 94.385 35.010 95.110 ;
        RECT 35.180 94.215 35.440 94.940 ;
        RECT 35.610 94.315 35.870 95.110 ;
        RECT 30.035 94.200 35.440 94.215 ;
        RECT 28.695 93.975 35.440 94.200 ;
        RECT 28.695 93.385 29.860 93.975 ;
        RECT 36.040 93.805 36.290 94.940 ;
        RECT 36.470 94.305 36.730 95.115 ;
        RECT 36.905 93.805 37.150 94.945 ;
        RECT 37.330 94.305 37.625 95.115 ;
        RECT 37.805 94.040 38.075 94.945 ;
        RECT 38.245 94.355 38.575 95.115 ;
        RECT 38.755 94.185 38.925 94.945 ;
        RECT 30.030 93.555 37.150 93.805 ;
        RECT 28.695 93.215 35.440 93.385 ;
        RECT 27.455 92.565 27.705 93.025 ;
        RECT 27.875 92.735 28.435 93.025 ;
        RECT 28.695 92.565 28.995 93.045 ;
        RECT 29.165 92.760 29.425 93.215 ;
        RECT 29.595 92.565 29.855 93.045 ;
        RECT 30.035 92.760 30.295 93.215 ;
        RECT 30.465 92.565 30.715 93.045 ;
        RECT 30.895 92.760 31.155 93.215 ;
        RECT 31.325 92.565 31.575 93.045 ;
        RECT 31.755 92.760 32.015 93.215 ;
        RECT 32.185 92.565 32.430 93.045 ;
        RECT 32.600 92.760 32.875 93.215 ;
        RECT 33.045 92.565 33.290 93.045 ;
        RECT 33.460 92.760 33.720 93.215 ;
        RECT 33.890 92.565 34.150 93.045 ;
        RECT 34.320 92.760 34.580 93.215 ;
        RECT 34.750 92.565 35.010 93.045 ;
        RECT 35.180 92.760 35.440 93.215 ;
        RECT 35.610 92.565 35.870 93.125 ;
        RECT 36.040 92.745 36.290 93.555 ;
        RECT 36.470 92.565 36.730 93.090 ;
        RECT 36.900 92.745 37.150 93.555 ;
        RECT 37.320 93.245 37.635 93.805 ;
        RECT 37.805 93.240 37.975 94.040 ;
        RECT 38.260 94.015 38.925 94.185 ;
        RECT 39.645 94.355 40.160 94.765 ;
        RECT 40.395 94.355 40.565 95.115 ;
        RECT 40.735 94.775 42.765 94.945 ;
        RECT 38.260 93.870 38.430 94.015 ;
        RECT 38.145 93.540 38.430 93.870 ;
        RECT 38.260 93.285 38.430 93.540 ;
        RECT 38.665 93.465 38.995 93.835 ;
        RECT 39.645 93.545 39.985 94.355 ;
        RECT 40.735 94.110 40.905 94.775 ;
        RECT 41.300 94.435 42.425 94.605 ;
        RECT 40.155 93.920 40.905 94.110 ;
        RECT 41.075 94.095 42.085 94.265 ;
        RECT 39.645 93.375 40.875 93.545 ;
        RECT 37.330 92.565 37.635 93.075 ;
        RECT 37.805 92.735 38.065 93.240 ;
        RECT 38.260 93.115 38.925 93.285 ;
        RECT 38.245 92.565 38.575 92.945 ;
        RECT 38.755 92.735 38.925 93.115 ;
        RECT 39.920 92.770 40.165 93.375 ;
        RECT 40.385 92.565 40.895 93.100 ;
        RECT 41.075 92.735 41.265 94.095 ;
        RECT 41.435 93.755 41.710 93.895 ;
        RECT 41.435 93.585 41.715 93.755 ;
        RECT 41.435 92.735 41.710 93.585 ;
        RECT 41.915 93.295 42.085 94.095 ;
        RECT 42.255 93.305 42.425 94.435 ;
        RECT 42.595 93.805 42.765 94.775 ;
        RECT 42.935 93.975 43.105 95.115 ;
        RECT 43.275 93.975 43.610 94.945 ;
        RECT 42.595 93.475 42.790 93.805 ;
        RECT 43.015 93.475 43.270 93.805 ;
        RECT 43.015 93.305 43.185 93.475 ;
        RECT 43.440 93.305 43.610 93.975 ;
        RECT 44.245 93.950 44.535 95.115 ;
        RECT 44.705 94.040 44.975 94.945 ;
        RECT 45.145 94.355 45.475 95.115 ;
        RECT 45.655 94.185 45.825 94.945 ;
        RECT 42.255 93.135 43.185 93.305 ;
        RECT 42.255 93.100 42.430 93.135 ;
        RECT 41.900 92.735 42.430 93.100 ;
        RECT 42.855 92.565 43.185 92.965 ;
        RECT 43.355 92.735 43.610 93.305 ;
        RECT 44.245 92.565 44.535 93.290 ;
        RECT 44.705 93.240 44.875 94.040 ;
        RECT 45.160 94.015 45.825 94.185 ;
        RECT 46.085 94.025 47.755 95.115 ;
        RECT 48.125 94.445 48.405 95.115 ;
        RECT 48.575 94.225 48.875 94.775 ;
        RECT 49.075 94.395 49.405 95.115 ;
        RECT 49.595 94.395 50.055 94.945 ;
        RECT 45.160 93.870 45.330 94.015 ;
        RECT 45.045 93.540 45.330 93.870 ;
        RECT 45.160 93.285 45.330 93.540 ;
        RECT 45.565 93.465 45.895 93.835 ;
        RECT 46.085 93.335 46.835 93.855 ;
        RECT 47.005 93.505 47.755 94.025 ;
        RECT 47.940 93.805 48.205 94.165 ;
        RECT 48.575 94.055 49.515 94.225 ;
        RECT 49.345 93.805 49.515 94.055 ;
        RECT 47.940 93.555 48.615 93.805 ;
        RECT 48.835 93.555 49.175 93.805 ;
        RECT 49.345 93.475 49.635 93.805 ;
        RECT 49.345 93.385 49.515 93.475 ;
        RECT 44.705 92.735 44.965 93.240 ;
        RECT 45.160 93.115 45.825 93.285 ;
        RECT 45.145 92.565 45.475 92.945 ;
        RECT 45.655 92.735 45.825 93.115 ;
        RECT 46.085 92.565 47.755 93.335 ;
        RECT 48.125 93.195 49.515 93.385 ;
        RECT 48.125 92.835 48.455 93.195 ;
        RECT 49.805 93.025 50.055 94.395 ;
        RECT 49.075 92.565 49.325 93.025 ;
        RECT 49.495 92.735 50.055 93.025 ;
        RECT 50.230 93.975 50.565 94.945 ;
        RECT 50.735 93.975 50.905 95.115 ;
        RECT 51.075 94.775 53.105 94.945 ;
        RECT 50.230 93.305 50.400 93.975 ;
        RECT 51.075 93.805 51.245 94.775 ;
        RECT 50.570 93.475 50.825 93.805 ;
        RECT 51.050 93.475 51.245 93.805 ;
        RECT 51.415 94.435 52.540 94.605 ;
        RECT 50.655 93.305 50.825 93.475 ;
        RECT 51.415 93.305 51.585 94.435 ;
        RECT 50.230 92.735 50.485 93.305 ;
        RECT 50.655 93.135 51.585 93.305 ;
        RECT 51.755 94.095 52.765 94.265 ;
        RECT 51.755 93.295 51.925 94.095 ;
        RECT 52.130 93.755 52.405 93.895 ;
        RECT 52.125 93.585 52.405 93.755 ;
        RECT 51.410 93.100 51.585 93.135 ;
        RECT 50.655 92.565 50.985 92.965 ;
        RECT 51.410 92.735 51.940 93.100 ;
        RECT 52.130 92.735 52.405 93.585 ;
        RECT 52.575 92.735 52.765 94.095 ;
        RECT 52.935 94.110 53.105 94.775 ;
        RECT 53.275 94.355 53.445 95.115 ;
        RECT 53.680 94.355 54.195 94.765 ;
        RECT 52.935 93.920 53.685 94.110 ;
        RECT 53.855 93.545 54.195 94.355 ;
        RECT 52.965 93.375 54.195 93.545 ;
        RECT 54.365 94.395 54.825 94.945 ;
        RECT 55.015 94.395 55.345 95.115 ;
        RECT 52.945 92.565 53.455 93.100 ;
        RECT 53.675 92.770 53.920 93.375 ;
        RECT 54.365 93.025 54.615 94.395 ;
        RECT 55.545 94.225 55.845 94.775 ;
        RECT 56.015 94.445 56.295 95.115 ;
        RECT 54.905 94.055 55.845 94.225 ;
        RECT 56.665 94.395 57.125 94.945 ;
        RECT 57.315 94.395 57.645 95.115 ;
        RECT 54.905 93.805 55.075 94.055 ;
        RECT 56.215 93.805 56.480 94.165 ;
        RECT 54.785 93.475 55.075 93.805 ;
        RECT 55.245 93.555 55.585 93.805 ;
        RECT 55.805 93.555 56.480 93.805 ;
        RECT 54.905 93.385 55.075 93.475 ;
        RECT 54.905 93.195 56.295 93.385 ;
        RECT 54.365 92.735 54.925 93.025 ;
        RECT 55.095 92.565 55.345 93.025 ;
        RECT 55.965 92.835 56.295 93.195 ;
        RECT 56.665 93.025 56.915 94.395 ;
        RECT 57.845 94.225 58.145 94.775 ;
        RECT 58.315 94.445 58.595 95.115 ;
        RECT 59.055 94.445 59.225 94.945 ;
        RECT 59.395 94.615 59.725 95.115 ;
        RECT 59.055 94.275 59.720 94.445 ;
        RECT 57.205 94.055 58.145 94.225 ;
        RECT 57.205 93.805 57.375 94.055 ;
        RECT 58.515 93.805 58.780 94.165 ;
        RECT 57.085 93.475 57.375 93.805 ;
        RECT 57.545 93.555 57.885 93.805 ;
        RECT 58.105 93.555 58.780 93.805 ;
        RECT 57.205 93.385 57.375 93.475 ;
        RECT 58.970 93.455 59.320 94.105 ;
        RECT 57.205 93.195 58.595 93.385 ;
        RECT 59.490 93.285 59.720 94.275 ;
        RECT 56.665 92.735 57.225 93.025 ;
        RECT 57.395 92.565 57.645 93.025 ;
        RECT 58.265 92.835 58.595 93.195 ;
        RECT 59.055 93.115 59.720 93.285 ;
        RECT 59.055 92.825 59.225 93.115 ;
        RECT 59.395 92.565 59.725 92.945 ;
        RECT 59.895 92.825 60.120 94.945 ;
        RECT 60.335 94.615 60.665 95.115 ;
        RECT 60.835 94.445 61.005 94.945 ;
        RECT 61.240 94.730 62.070 94.900 ;
        RECT 62.310 94.735 62.690 95.115 ;
        RECT 60.310 94.275 61.005 94.445 ;
        RECT 60.310 93.305 60.480 94.275 ;
        RECT 60.650 93.485 61.060 94.105 ;
        RECT 61.230 94.055 61.730 94.435 ;
        RECT 60.310 93.115 61.005 93.305 ;
        RECT 61.230 93.185 61.450 94.055 ;
        RECT 61.900 93.885 62.070 94.730 ;
        RECT 62.870 94.565 63.040 94.855 ;
        RECT 63.210 94.735 63.540 95.115 ;
        RECT 64.010 94.645 64.640 94.895 ;
        RECT 64.820 94.735 65.240 95.115 ;
        RECT 64.470 94.565 64.640 94.645 ;
        RECT 65.440 94.565 65.680 94.855 ;
        RECT 62.240 94.315 63.610 94.565 ;
        RECT 62.240 94.055 62.490 94.315 ;
        RECT 63.000 93.885 63.250 94.045 ;
        RECT 61.900 93.715 63.250 93.885 ;
        RECT 61.900 93.675 62.320 93.715 ;
        RECT 61.630 93.125 61.980 93.495 ;
        RECT 60.335 92.565 60.665 92.945 ;
        RECT 60.835 92.785 61.005 93.115 ;
        RECT 62.150 92.945 62.320 93.675 ;
        RECT 63.420 93.545 63.610 94.315 ;
        RECT 62.490 93.215 62.900 93.545 ;
        RECT 63.190 93.205 63.610 93.545 ;
        RECT 63.780 94.135 64.300 94.445 ;
        RECT 64.470 94.395 65.680 94.565 ;
        RECT 65.910 94.425 66.240 95.115 ;
        RECT 63.780 93.375 63.950 94.135 ;
        RECT 64.120 93.545 64.300 93.955 ;
        RECT 64.470 93.885 64.640 94.395 ;
        RECT 66.410 94.245 66.580 94.855 ;
        RECT 66.850 94.395 67.180 94.905 ;
        RECT 66.410 94.225 66.730 94.245 ;
        RECT 64.810 94.055 66.730 94.225 ;
        RECT 64.470 93.715 66.370 93.885 ;
        RECT 64.700 93.375 65.030 93.495 ;
        RECT 63.780 93.205 65.030 93.375 ;
        RECT 61.305 92.745 62.320 92.945 ;
        RECT 62.490 92.565 62.900 93.005 ;
        RECT 63.190 92.775 63.440 93.205 ;
        RECT 63.640 92.565 63.960 93.025 ;
        RECT 65.200 92.955 65.370 93.715 ;
        RECT 66.040 93.655 66.370 93.715 ;
        RECT 65.560 93.485 65.890 93.545 ;
        RECT 65.560 93.215 66.220 93.485 ;
        RECT 66.540 93.160 66.730 94.055 ;
        RECT 64.520 92.785 65.370 92.955 ;
        RECT 65.570 92.565 66.230 93.045 ;
        RECT 66.410 92.830 66.730 93.160 ;
        RECT 66.930 93.805 67.180 94.395 ;
        RECT 67.360 94.315 67.645 95.115 ;
        RECT 67.825 94.135 68.080 94.805 ;
        RECT 66.930 93.475 67.730 93.805 ;
        RECT 66.930 92.825 67.180 93.475 ;
        RECT 67.900 93.275 68.080 94.135 ;
        RECT 68.625 94.025 69.835 95.115 ;
        RECT 67.825 93.075 68.080 93.275 ;
        RECT 68.625 93.315 69.145 93.855 ;
        RECT 69.315 93.485 69.835 94.025 ;
        RECT 70.005 93.950 70.295 95.115 ;
        RECT 70.465 94.025 73.975 95.115 ;
        RECT 70.465 93.335 72.115 93.855 ;
        RECT 72.285 93.505 73.975 94.025 ;
        RECT 74.610 93.975 74.945 94.945 ;
        RECT 75.115 93.975 75.285 95.115 ;
        RECT 75.455 94.775 77.485 94.945 ;
        RECT 67.360 92.565 67.645 93.025 ;
        RECT 67.825 92.905 68.165 93.075 ;
        RECT 67.825 92.745 68.080 92.905 ;
        RECT 68.625 92.565 69.835 93.315 ;
        RECT 70.005 92.565 70.295 93.290 ;
        RECT 70.465 92.565 73.975 93.335 ;
        RECT 74.610 93.305 74.780 93.975 ;
        RECT 75.455 93.805 75.625 94.775 ;
        RECT 74.950 93.475 75.205 93.805 ;
        RECT 75.430 93.475 75.625 93.805 ;
        RECT 75.795 94.435 76.920 94.605 ;
        RECT 75.035 93.305 75.205 93.475 ;
        RECT 75.795 93.305 75.965 94.435 ;
        RECT 74.610 92.735 74.865 93.305 ;
        RECT 75.035 93.135 75.965 93.305 ;
        RECT 76.135 94.095 77.145 94.265 ;
        RECT 76.135 93.295 76.305 94.095 ;
        RECT 75.790 93.100 75.965 93.135 ;
        RECT 75.035 92.565 75.365 92.965 ;
        RECT 75.790 92.735 76.320 93.100 ;
        RECT 76.510 93.075 76.785 93.895 ;
        RECT 76.505 92.905 76.785 93.075 ;
        RECT 76.510 92.735 76.785 92.905 ;
        RECT 76.955 92.735 77.145 94.095 ;
        RECT 77.315 94.110 77.485 94.775 ;
        RECT 77.655 94.355 77.825 95.115 ;
        RECT 78.060 94.355 78.575 94.765 ;
        RECT 77.315 93.920 78.065 94.110 ;
        RECT 78.235 93.545 78.575 94.355 ;
        RECT 78.745 94.025 82.255 95.115 ;
        RECT 82.425 94.025 83.635 95.115 ;
        RECT 77.345 93.375 78.575 93.545 ;
        RECT 77.325 92.565 77.835 93.100 ;
        RECT 78.055 92.770 78.300 93.375 ;
        RECT 78.745 93.335 80.395 93.855 ;
        RECT 80.565 93.505 82.255 94.025 ;
        RECT 78.745 92.565 82.255 93.335 ;
        RECT 82.425 93.315 82.945 93.855 ;
        RECT 83.115 93.485 83.635 94.025 ;
        RECT 83.805 94.395 84.265 94.945 ;
        RECT 84.455 94.395 84.785 95.115 ;
        RECT 82.425 92.565 83.635 93.315 ;
        RECT 83.805 93.025 84.055 94.395 ;
        RECT 84.985 94.225 85.285 94.775 ;
        RECT 85.455 94.445 85.735 95.115 ;
        RECT 84.345 94.055 85.285 94.225 ;
        RECT 84.345 93.805 84.515 94.055 ;
        RECT 85.655 93.805 85.920 94.165 ;
        RECT 86.115 93.975 86.445 95.115 ;
        RECT 84.225 93.475 84.515 93.805 ;
        RECT 84.685 93.555 85.025 93.805 ;
        RECT 85.245 93.555 85.920 93.805 ;
        RECT 84.345 93.385 84.515 93.475 ;
        RECT 84.345 93.195 85.735 93.385 ;
        RECT 86.105 93.225 86.445 93.805 ;
        RECT 86.615 93.775 86.975 94.945 ;
        RECT 87.175 93.945 87.505 95.115 ;
        RECT 87.705 93.775 88.035 94.945 ;
        RECT 88.235 93.945 88.565 95.115 ;
        RECT 88.865 94.395 89.325 94.945 ;
        RECT 89.515 94.395 89.845 95.115 ;
        RECT 86.615 93.495 88.035 93.775 ;
        RECT 83.805 92.735 84.365 93.025 ;
        RECT 84.535 92.565 84.785 93.025 ;
        RECT 85.405 92.835 85.735 93.195 ;
        RECT 86.615 93.160 86.975 93.495 ;
        RECT 86.115 92.565 86.445 93.055 ;
        RECT 86.615 92.735 87.235 93.160 ;
        RECT 87.695 92.565 88.025 93.255 ;
        RECT 88.865 93.025 89.115 94.395 ;
        RECT 90.045 94.225 90.345 94.775 ;
        RECT 90.515 94.445 90.795 95.115 ;
        RECT 89.405 94.055 90.345 94.225 ;
        RECT 91.165 94.395 91.625 94.945 ;
        RECT 91.815 94.395 92.145 95.115 ;
        RECT 89.405 93.805 89.575 94.055 ;
        RECT 90.715 93.805 90.980 94.165 ;
        RECT 89.285 93.475 89.575 93.805 ;
        RECT 89.745 93.555 90.085 93.805 ;
        RECT 90.305 93.555 90.980 93.805 ;
        RECT 89.405 93.385 89.575 93.475 ;
        RECT 89.405 93.195 90.795 93.385 ;
        RECT 88.865 92.735 89.425 93.025 ;
        RECT 89.595 92.565 89.845 93.025 ;
        RECT 90.465 92.835 90.795 93.195 ;
        RECT 91.165 93.025 91.415 94.395 ;
        RECT 92.345 94.225 92.645 94.775 ;
        RECT 92.815 94.445 93.095 95.115 ;
        RECT 91.705 94.055 92.645 94.225 ;
        RECT 93.555 94.185 93.725 94.945 ;
        RECT 93.905 94.355 94.235 95.115 ;
        RECT 91.705 93.805 91.875 94.055 ;
        RECT 93.015 93.805 93.280 94.165 ;
        RECT 93.555 94.015 94.220 94.185 ;
        RECT 94.405 94.040 94.675 94.945 ;
        RECT 94.050 93.870 94.220 94.015 ;
        RECT 91.585 93.475 91.875 93.805 ;
        RECT 92.045 93.555 92.385 93.805 ;
        RECT 92.605 93.555 93.280 93.805 ;
        RECT 91.705 93.385 91.875 93.475 ;
        RECT 93.485 93.465 93.815 93.835 ;
        RECT 94.050 93.540 94.335 93.870 ;
        RECT 91.705 93.195 93.095 93.385 ;
        RECT 94.050 93.285 94.220 93.540 ;
        RECT 91.165 92.735 91.725 93.025 ;
        RECT 91.895 92.565 92.145 93.025 ;
        RECT 92.765 92.835 93.095 93.195 ;
        RECT 93.555 93.115 94.220 93.285 ;
        RECT 94.505 93.240 94.675 94.040 ;
        RECT 95.765 93.950 96.055 95.115 ;
        RECT 96.225 94.025 97.895 95.115 ;
        RECT 96.225 93.335 96.975 93.855 ;
        RECT 97.145 93.505 97.895 94.025 ;
        RECT 98.585 93.975 98.795 95.115 ;
        RECT 98.965 93.965 99.295 94.945 ;
        RECT 99.465 93.975 99.695 95.115 ;
        RECT 99.905 94.680 105.250 95.115 ;
        RECT 93.555 92.735 93.725 93.115 ;
        RECT 93.905 92.565 94.235 92.945 ;
        RECT 94.415 92.735 94.675 93.240 ;
        RECT 95.765 92.565 96.055 93.290 ;
        RECT 96.225 92.565 97.895 93.335 ;
        RECT 98.585 92.565 98.795 93.385 ;
        RECT 98.965 93.365 99.215 93.965 ;
        RECT 99.385 93.555 99.715 93.805 ;
        RECT 98.965 92.735 99.295 93.365 ;
        RECT 99.465 92.565 99.695 93.385 ;
        RECT 101.490 93.110 101.830 93.940 ;
        RECT 103.310 93.430 103.660 94.680 ;
        RECT 106.435 94.445 106.605 94.945 ;
        RECT 106.775 94.615 107.105 95.115 ;
        RECT 106.435 94.275 107.100 94.445 ;
        RECT 106.350 93.455 106.700 94.105 ;
        RECT 106.870 93.285 107.100 94.275 ;
        RECT 106.435 93.115 107.100 93.285 ;
        RECT 99.905 92.565 105.250 93.110 ;
        RECT 106.435 92.825 106.605 93.115 ;
        RECT 106.775 92.565 107.105 92.945 ;
        RECT 107.275 92.825 107.500 94.945 ;
        RECT 107.715 94.615 108.045 95.115 ;
        RECT 108.215 94.445 108.385 94.945 ;
        RECT 108.620 94.730 109.450 94.900 ;
        RECT 109.690 94.735 110.070 95.115 ;
        RECT 107.690 94.275 108.385 94.445 ;
        RECT 107.690 93.305 107.860 94.275 ;
        RECT 108.030 93.485 108.440 94.105 ;
        RECT 108.610 94.055 109.110 94.435 ;
        RECT 107.690 93.115 108.385 93.305 ;
        RECT 108.610 93.185 108.830 94.055 ;
        RECT 109.280 93.885 109.450 94.730 ;
        RECT 110.250 94.565 110.420 94.855 ;
        RECT 110.590 94.735 110.920 95.115 ;
        RECT 111.390 94.645 112.020 94.895 ;
        RECT 112.200 94.735 112.620 95.115 ;
        RECT 111.850 94.565 112.020 94.645 ;
        RECT 112.820 94.565 113.060 94.855 ;
        RECT 109.620 94.315 110.990 94.565 ;
        RECT 109.620 94.055 109.870 94.315 ;
        RECT 110.380 93.885 110.630 94.045 ;
        RECT 109.280 93.715 110.630 93.885 ;
        RECT 109.280 93.675 109.700 93.715 ;
        RECT 109.010 93.125 109.360 93.495 ;
        RECT 107.715 92.565 108.045 92.945 ;
        RECT 108.215 92.785 108.385 93.115 ;
        RECT 109.530 92.945 109.700 93.675 ;
        RECT 110.800 93.545 110.990 94.315 ;
        RECT 109.870 93.215 110.280 93.545 ;
        RECT 110.570 93.205 110.990 93.545 ;
        RECT 111.160 94.135 111.680 94.445 ;
        RECT 111.850 94.395 113.060 94.565 ;
        RECT 113.290 94.425 113.620 95.115 ;
        RECT 111.160 93.375 111.330 94.135 ;
        RECT 111.500 93.545 111.680 93.955 ;
        RECT 111.850 93.885 112.020 94.395 ;
        RECT 113.790 94.245 113.960 94.855 ;
        RECT 114.230 94.395 114.560 94.905 ;
        RECT 113.790 94.225 114.110 94.245 ;
        RECT 112.190 94.055 114.110 94.225 ;
        RECT 111.850 93.715 113.750 93.885 ;
        RECT 112.080 93.375 112.410 93.495 ;
        RECT 111.160 93.205 112.410 93.375 ;
        RECT 108.685 92.745 109.700 92.945 ;
        RECT 109.870 92.565 110.280 93.005 ;
        RECT 110.570 92.775 110.820 93.205 ;
        RECT 111.020 92.565 111.340 93.025 ;
        RECT 112.580 92.955 112.750 93.715 ;
        RECT 113.420 93.655 113.750 93.715 ;
        RECT 112.940 93.485 113.270 93.545 ;
        RECT 112.940 93.215 113.600 93.485 ;
        RECT 113.920 93.160 114.110 94.055 ;
        RECT 111.900 92.785 112.750 92.955 ;
        RECT 112.950 92.565 113.610 93.045 ;
        RECT 113.790 92.830 114.110 93.160 ;
        RECT 114.310 93.805 114.560 94.395 ;
        RECT 114.740 94.315 115.025 95.115 ;
        RECT 115.205 94.135 115.460 94.805 ;
        RECT 114.310 93.475 115.110 93.805 ;
        RECT 114.310 92.825 114.560 93.475 ;
        RECT 115.280 93.275 115.460 94.135 ;
        RECT 116.005 94.025 117.215 95.115 ;
        RECT 115.205 93.075 115.460 93.275 ;
        RECT 116.005 93.315 116.525 93.855 ;
        RECT 116.695 93.485 117.215 94.025 ;
        RECT 117.385 94.025 118.595 95.115 ;
        RECT 117.385 93.485 117.905 94.025 ;
        RECT 118.075 93.315 118.595 93.855 ;
        RECT 114.740 92.565 115.025 93.025 ;
        RECT 115.205 92.905 115.545 93.075 ;
        RECT 115.205 92.745 115.460 92.905 ;
        RECT 116.005 92.565 117.215 93.315 ;
        RECT 117.385 92.565 118.595 93.315 ;
        RECT 5.520 92.395 118.680 92.565 ;
        RECT 5.605 91.645 6.815 92.395 ;
        RECT 6.985 91.850 12.330 92.395 ;
        RECT 12.505 91.850 17.850 92.395 ;
        RECT 5.605 91.105 6.125 91.645 ;
        RECT 6.295 90.935 6.815 91.475 ;
        RECT 8.570 91.020 8.910 91.850 ;
        RECT 5.605 89.845 6.815 90.935 ;
        RECT 10.390 90.280 10.740 91.530 ;
        RECT 14.090 91.020 14.430 91.850 ;
        RECT 18.025 91.625 20.615 92.395 ;
        RECT 21.445 91.765 21.775 92.125 ;
        RECT 22.395 91.935 22.645 92.395 ;
        RECT 22.815 91.935 23.375 92.225 ;
        RECT 15.910 90.280 16.260 91.530 ;
        RECT 18.025 91.105 19.235 91.625 ;
        RECT 21.445 91.575 22.835 91.765 ;
        RECT 22.665 91.485 22.835 91.575 ;
        RECT 19.405 90.935 20.615 91.455 ;
        RECT 6.985 89.845 12.330 90.280 ;
        RECT 12.505 89.845 17.850 90.280 ;
        RECT 18.025 89.845 20.615 90.935 ;
        RECT 21.260 91.155 21.935 91.405 ;
        RECT 22.155 91.155 22.495 91.405 ;
        RECT 22.665 91.155 22.955 91.485 ;
        RECT 21.260 90.795 21.525 91.155 ;
        RECT 22.665 90.905 22.835 91.155 ;
        RECT 21.895 90.735 22.835 90.905 ;
        RECT 21.445 89.845 21.725 90.515 ;
        RECT 21.895 90.185 22.195 90.735 ;
        RECT 23.125 90.565 23.375 91.935 ;
        RECT 23.545 91.850 28.890 92.395 ;
        RECT 25.130 91.020 25.470 91.850 ;
        RECT 29.065 91.625 30.735 92.395 ;
        RECT 31.365 91.670 31.655 92.395 ;
        RECT 31.835 91.745 32.165 92.220 ;
        RECT 32.335 91.915 32.505 92.395 ;
        RECT 32.675 91.745 33.005 92.220 ;
        RECT 33.175 91.915 33.345 92.395 ;
        RECT 33.515 91.745 33.845 92.220 ;
        RECT 34.015 91.915 34.185 92.395 ;
        RECT 34.355 91.745 34.685 92.220 ;
        RECT 34.855 91.915 35.025 92.395 ;
        RECT 35.195 91.745 35.525 92.220 ;
        RECT 35.695 91.915 35.865 92.395 ;
        RECT 36.035 92.220 36.285 92.225 ;
        RECT 36.035 91.745 36.365 92.220 ;
        RECT 36.535 91.915 36.705 92.395 ;
        RECT 36.955 92.220 37.125 92.225 ;
        RECT 36.875 91.745 37.205 92.220 ;
        RECT 37.375 91.915 37.545 92.395 ;
        RECT 37.795 92.220 37.965 92.225 ;
        RECT 37.715 91.745 38.045 92.220 ;
        RECT 38.215 91.915 38.385 92.395 ;
        RECT 38.555 91.745 38.885 92.220 ;
        RECT 39.055 91.915 39.225 92.395 ;
        RECT 39.395 91.745 39.725 92.220 ;
        RECT 39.895 91.915 40.065 92.395 ;
        RECT 40.235 91.745 40.565 92.220 ;
        RECT 40.735 91.915 40.905 92.395 ;
        RECT 41.075 91.745 41.405 92.220 ;
        RECT 41.575 91.915 41.745 92.395 ;
        RECT 41.915 91.745 42.245 92.220 ;
        RECT 42.415 91.915 42.585 92.395 ;
        RECT 22.395 89.845 22.725 90.565 ;
        RECT 22.915 90.015 23.375 90.565 ;
        RECT 26.950 90.280 27.300 91.530 ;
        RECT 29.065 91.105 29.815 91.625 ;
        RECT 31.835 91.575 33.345 91.745 ;
        RECT 33.515 91.575 35.865 91.745 ;
        RECT 36.035 91.575 42.695 91.745 ;
        RECT 42.925 91.575 43.135 92.395 ;
        RECT 43.305 91.595 43.635 92.225 ;
        RECT 29.985 90.935 30.735 91.455 ;
        RECT 33.175 91.405 33.345 91.575 ;
        RECT 35.690 91.405 35.865 91.575 ;
        RECT 31.830 91.205 33.005 91.405 ;
        RECT 33.175 91.205 35.485 91.405 ;
        RECT 35.690 91.205 42.250 91.405 ;
        RECT 33.175 91.035 33.345 91.205 ;
        RECT 35.690 91.035 35.865 91.205 ;
        RECT 42.420 91.035 42.695 91.575 ;
        RECT 23.545 89.845 28.890 90.280 ;
        RECT 29.065 89.845 30.735 90.935 ;
        RECT 31.365 89.845 31.655 91.010 ;
        RECT 31.835 90.865 33.345 91.035 ;
        RECT 33.515 90.865 35.865 91.035 ;
        RECT 36.035 90.865 42.695 91.035 ;
        RECT 43.305 90.995 43.555 91.595 ;
        RECT 43.805 91.575 44.035 92.395 ;
        RECT 44.245 91.850 49.590 92.395 ;
        RECT 43.725 91.155 44.055 91.405 ;
        RECT 45.830 91.020 46.170 91.850 ;
        RECT 49.765 91.625 52.355 92.395 ;
        RECT 52.725 91.765 53.055 92.125 ;
        RECT 53.675 91.935 53.925 92.395 ;
        RECT 54.095 91.935 54.655 92.225 ;
        RECT 31.835 90.015 32.165 90.865 ;
        RECT 32.335 89.845 32.505 90.695 ;
        RECT 32.675 90.015 33.005 90.865 ;
        RECT 33.175 89.845 33.345 90.695 ;
        RECT 33.515 90.015 33.845 90.865 ;
        RECT 34.015 89.845 34.185 90.645 ;
        RECT 34.355 90.015 34.685 90.865 ;
        RECT 34.855 89.845 35.025 90.645 ;
        RECT 35.195 90.015 35.525 90.865 ;
        RECT 35.695 89.845 35.865 90.645 ;
        RECT 36.035 90.015 36.365 90.865 ;
        RECT 36.535 89.845 36.705 90.645 ;
        RECT 36.875 90.015 37.205 90.865 ;
        RECT 37.375 89.845 37.545 90.645 ;
        RECT 37.715 90.015 38.045 90.865 ;
        RECT 38.215 89.845 38.385 90.645 ;
        RECT 38.555 90.015 38.885 90.865 ;
        RECT 39.055 89.845 39.225 90.645 ;
        RECT 39.395 90.015 39.725 90.865 ;
        RECT 39.895 89.845 40.065 90.645 ;
        RECT 40.235 90.015 40.565 90.865 ;
        RECT 40.735 89.845 40.905 90.645 ;
        RECT 41.075 90.015 41.405 90.865 ;
        RECT 41.575 89.845 41.745 90.645 ;
        RECT 41.915 90.015 42.245 90.865 ;
        RECT 42.415 89.845 42.585 90.645 ;
        RECT 42.925 89.845 43.135 90.985 ;
        RECT 43.305 90.015 43.635 90.995 ;
        RECT 43.805 89.845 44.035 90.985 ;
        RECT 47.650 90.280 48.000 91.530 ;
        RECT 49.765 91.105 50.975 91.625 ;
        RECT 52.725 91.575 54.115 91.765 ;
        RECT 53.945 91.485 54.115 91.575 ;
        RECT 51.145 90.935 52.355 91.455 ;
        RECT 44.245 89.845 49.590 90.280 ;
        RECT 49.765 89.845 52.355 90.935 ;
        RECT 52.540 91.155 53.215 91.405 ;
        RECT 53.435 91.155 53.775 91.405 ;
        RECT 53.945 91.155 54.235 91.485 ;
        RECT 52.540 90.795 52.805 91.155 ;
        RECT 53.945 90.905 54.115 91.155 ;
        RECT 53.175 90.735 54.115 90.905 ;
        RECT 52.725 89.845 53.005 90.515 ;
        RECT 53.175 90.185 53.475 90.735 ;
        RECT 54.405 90.565 54.655 91.935 ;
        RECT 54.825 91.625 56.495 92.395 ;
        RECT 57.125 91.670 57.415 92.395 ;
        RECT 57.590 91.995 57.925 92.395 ;
        RECT 58.095 91.825 58.300 92.225 ;
        RECT 58.510 91.915 58.785 92.395 ;
        RECT 58.995 91.895 59.255 92.225 ;
        RECT 57.615 91.655 58.300 91.825 ;
        RECT 54.825 91.105 55.575 91.625 ;
        RECT 55.745 90.935 56.495 91.455 ;
        RECT 53.675 89.845 54.005 90.565 ;
        RECT 54.195 90.015 54.655 90.565 ;
        RECT 54.825 89.845 56.495 90.935 ;
        RECT 57.125 89.845 57.415 91.010 ;
        RECT 57.615 90.625 57.955 91.655 ;
        RECT 58.125 90.985 58.375 91.485 ;
        RECT 58.555 91.155 58.915 91.735 ;
        RECT 59.085 90.985 59.255 91.895 ;
        RECT 59.625 91.765 59.955 92.125 ;
        RECT 60.575 91.935 60.825 92.395 ;
        RECT 60.995 91.935 61.555 92.225 ;
        RECT 59.625 91.575 61.015 91.765 ;
        RECT 60.845 91.485 61.015 91.575 ;
        RECT 58.125 90.815 59.255 90.985 ;
        RECT 57.615 90.450 58.280 90.625 ;
        RECT 57.590 89.845 57.925 90.270 ;
        RECT 58.095 90.045 58.280 90.450 ;
        RECT 58.485 89.845 58.815 90.625 ;
        RECT 58.985 90.045 59.255 90.815 ;
        RECT 59.440 91.155 60.115 91.405 ;
        RECT 60.335 91.155 60.675 91.405 ;
        RECT 60.845 91.155 61.135 91.485 ;
        RECT 59.440 90.795 59.705 91.155 ;
        RECT 60.845 90.905 61.015 91.155 ;
        RECT 60.075 90.735 61.015 90.905 ;
        RECT 59.625 89.845 59.905 90.515 ;
        RECT 60.075 90.185 60.375 90.735 ;
        RECT 61.305 90.565 61.555 91.935 ;
        RECT 60.575 89.845 60.905 90.565 ;
        RECT 61.095 90.015 61.555 90.565 ;
        RECT 61.725 91.895 61.985 92.225 ;
        RECT 62.195 91.915 62.470 92.395 ;
        RECT 61.725 90.985 61.895 91.895 ;
        RECT 62.680 91.825 62.885 92.225 ;
        RECT 63.055 91.995 63.390 92.395 ;
        RECT 62.065 91.155 62.425 91.735 ;
        RECT 62.680 91.655 63.365 91.825 ;
        RECT 62.605 90.985 62.855 91.485 ;
        RECT 61.725 90.815 62.855 90.985 ;
        RECT 61.725 90.045 61.995 90.815 ;
        RECT 63.025 90.625 63.365 91.655 ;
        RECT 62.165 89.845 62.495 90.625 ;
        RECT 62.700 90.450 63.365 90.625 ;
        RECT 63.570 91.655 63.825 92.225 ;
        RECT 63.995 91.995 64.325 92.395 ;
        RECT 64.750 91.860 65.280 92.225 ;
        RECT 64.750 91.825 64.925 91.860 ;
        RECT 63.995 91.655 64.925 91.825 ;
        RECT 65.470 91.715 65.745 92.225 ;
        RECT 63.570 90.985 63.740 91.655 ;
        RECT 63.995 91.485 64.165 91.655 ;
        RECT 63.910 91.155 64.165 91.485 ;
        RECT 64.390 91.155 64.585 91.485 ;
        RECT 62.700 90.045 62.885 90.450 ;
        RECT 63.055 89.845 63.390 90.270 ;
        RECT 63.570 90.015 63.905 90.985 ;
        RECT 64.075 89.845 64.245 90.985 ;
        RECT 64.415 90.185 64.585 91.155 ;
        RECT 64.755 90.525 64.925 91.655 ;
        RECT 65.095 90.865 65.265 91.665 ;
        RECT 65.465 91.545 65.745 91.715 ;
        RECT 65.470 91.065 65.745 91.545 ;
        RECT 65.915 90.865 66.105 92.225 ;
        RECT 66.285 91.860 66.795 92.395 ;
        RECT 67.015 91.585 67.260 92.190 ;
        RECT 67.705 91.850 73.050 92.395 ;
        RECT 73.225 91.850 78.570 92.395 ;
        RECT 66.305 91.415 67.535 91.585 ;
        RECT 65.095 90.695 66.105 90.865 ;
        RECT 66.275 90.850 67.025 91.040 ;
        RECT 64.755 90.355 65.880 90.525 ;
        RECT 66.275 90.185 66.445 90.850 ;
        RECT 67.195 90.605 67.535 91.415 ;
        RECT 69.290 91.020 69.630 91.850 ;
        RECT 64.415 90.015 66.445 90.185 ;
        RECT 66.615 89.845 66.785 90.605 ;
        RECT 67.020 90.195 67.535 90.605 ;
        RECT 71.110 90.280 71.460 91.530 ;
        RECT 74.810 91.020 75.150 91.850 ;
        RECT 78.745 91.625 82.255 92.395 ;
        RECT 82.885 91.670 83.175 92.395 ;
        RECT 84.265 91.885 84.570 92.395 ;
        RECT 76.630 90.280 76.980 91.530 ;
        RECT 78.745 91.105 80.395 91.625 ;
        RECT 80.565 90.935 82.255 91.455 ;
        RECT 84.265 91.155 84.580 91.715 ;
        RECT 84.750 91.405 85.000 92.215 ;
        RECT 85.170 91.870 85.430 92.395 ;
        RECT 85.610 91.405 85.860 92.215 ;
        RECT 86.030 91.835 86.290 92.395 ;
        RECT 86.460 91.745 86.720 92.200 ;
        RECT 86.890 91.915 87.150 92.395 ;
        RECT 87.320 91.745 87.580 92.200 ;
        RECT 87.750 91.915 88.010 92.395 ;
        RECT 88.180 91.745 88.440 92.200 ;
        RECT 88.610 91.915 88.855 92.395 ;
        RECT 89.025 91.745 89.300 92.200 ;
        RECT 89.470 91.915 89.715 92.395 ;
        RECT 89.885 91.745 90.145 92.200 ;
        RECT 90.325 91.915 90.575 92.395 ;
        RECT 90.745 91.745 91.005 92.200 ;
        RECT 91.185 91.915 91.435 92.395 ;
        RECT 91.605 91.745 91.865 92.200 ;
        RECT 92.045 91.915 92.305 92.395 ;
        RECT 92.475 91.745 92.735 92.200 ;
        RECT 92.905 91.915 93.205 92.395 ;
        RECT 93.555 91.845 93.725 92.135 ;
        RECT 93.895 92.015 94.225 92.395 ;
        RECT 86.460 91.575 93.205 91.745 ;
        RECT 93.555 91.675 94.220 91.845 ;
        RECT 84.750 91.155 91.870 91.405 ;
        RECT 67.705 89.845 73.050 90.280 ;
        RECT 73.225 89.845 78.570 90.280 ;
        RECT 78.745 89.845 82.255 90.935 ;
        RECT 82.885 89.845 83.175 91.010 ;
        RECT 84.275 89.845 84.570 90.655 ;
        RECT 84.750 90.015 84.995 91.155 ;
        RECT 85.170 89.845 85.430 90.655 ;
        RECT 85.610 90.020 85.860 91.155 ;
        RECT 92.040 90.985 93.205 91.575 ;
        RECT 86.460 90.760 93.205 90.985 ;
        RECT 93.470 90.855 93.820 91.505 ;
        RECT 86.460 90.745 91.865 90.760 ;
        RECT 86.030 89.850 86.290 90.645 ;
        RECT 86.460 90.020 86.720 90.745 ;
        RECT 86.890 89.850 87.150 90.575 ;
        RECT 87.320 90.020 87.580 90.745 ;
        RECT 87.750 89.850 88.010 90.575 ;
        RECT 88.180 90.020 88.440 90.745 ;
        RECT 88.610 89.850 88.870 90.575 ;
        RECT 89.040 90.020 89.300 90.745 ;
        RECT 89.470 89.850 89.715 90.575 ;
        RECT 89.885 90.020 90.145 90.745 ;
        RECT 90.330 89.850 90.575 90.575 ;
        RECT 90.745 90.020 91.005 90.745 ;
        RECT 91.190 89.850 91.435 90.575 ;
        RECT 91.605 90.020 91.865 90.745 ;
        RECT 92.050 89.850 92.305 90.575 ;
        RECT 92.475 90.020 92.765 90.760 ;
        RECT 93.990 90.685 94.220 91.675 ;
        RECT 86.030 89.845 92.305 89.850 ;
        RECT 92.935 89.845 93.205 90.590 ;
        RECT 93.555 90.515 94.220 90.685 ;
        RECT 93.555 90.015 93.725 90.515 ;
        RECT 93.895 89.845 94.225 90.345 ;
        RECT 94.395 90.015 94.620 92.135 ;
        RECT 94.835 92.015 95.165 92.395 ;
        RECT 95.335 91.845 95.505 92.175 ;
        RECT 95.805 92.015 96.820 92.215 ;
        RECT 94.810 91.655 95.505 91.845 ;
        RECT 94.810 90.685 94.980 91.655 ;
        RECT 95.150 90.855 95.560 91.475 ;
        RECT 95.730 90.905 95.950 91.775 ;
        RECT 96.130 91.465 96.480 91.835 ;
        RECT 96.650 91.285 96.820 92.015 ;
        RECT 96.990 91.955 97.400 92.395 ;
        RECT 97.690 91.755 97.940 92.185 ;
        RECT 98.140 91.935 98.460 92.395 ;
        RECT 99.020 92.005 99.870 92.175 ;
        RECT 96.990 91.415 97.400 91.745 ;
        RECT 97.690 91.415 98.110 91.755 ;
        RECT 96.400 91.245 96.820 91.285 ;
        RECT 96.400 91.075 97.750 91.245 ;
        RECT 94.810 90.515 95.505 90.685 ;
        RECT 95.730 90.525 96.230 90.905 ;
        RECT 94.835 89.845 95.165 90.345 ;
        RECT 95.335 90.015 95.505 90.515 ;
        RECT 96.400 90.230 96.570 91.075 ;
        RECT 97.500 90.915 97.750 91.075 ;
        RECT 96.740 90.645 96.990 90.905 ;
        RECT 97.920 90.645 98.110 91.415 ;
        RECT 96.740 90.395 98.110 90.645 ;
        RECT 98.280 91.585 99.530 91.755 ;
        RECT 98.280 90.825 98.450 91.585 ;
        RECT 99.200 91.465 99.530 91.585 ;
        RECT 98.620 91.005 98.800 91.415 ;
        RECT 99.700 91.245 99.870 92.005 ;
        RECT 100.070 91.915 100.730 92.395 ;
        RECT 100.910 91.800 101.230 92.130 ;
        RECT 100.060 91.475 100.720 91.745 ;
        RECT 100.060 91.415 100.390 91.475 ;
        RECT 100.540 91.245 100.870 91.305 ;
        RECT 98.970 91.075 100.870 91.245 ;
        RECT 98.280 90.515 98.800 90.825 ;
        RECT 98.970 90.565 99.140 91.075 ;
        RECT 101.040 90.905 101.230 91.800 ;
        RECT 99.310 90.735 101.230 90.905 ;
        RECT 100.910 90.715 101.230 90.735 ;
        RECT 101.430 91.485 101.680 92.135 ;
        RECT 101.860 91.935 102.145 92.395 ;
        RECT 102.325 91.685 102.580 92.215 ;
        RECT 101.430 91.155 102.230 91.485 ;
        RECT 98.970 90.395 100.180 90.565 ;
        RECT 95.740 90.060 96.570 90.230 ;
        RECT 96.810 89.845 97.190 90.225 ;
        RECT 97.370 90.105 97.540 90.395 ;
        RECT 98.970 90.315 99.140 90.395 ;
        RECT 97.710 89.845 98.040 90.225 ;
        RECT 98.510 90.065 99.140 90.315 ;
        RECT 99.320 89.845 99.740 90.225 ;
        RECT 99.940 90.105 100.180 90.395 ;
        RECT 100.410 89.845 100.740 90.535 ;
        RECT 100.910 90.105 101.080 90.715 ;
        RECT 101.430 90.565 101.680 91.155 ;
        RECT 102.400 90.825 102.580 91.685 ;
        RECT 103.215 91.845 103.385 92.225 ;
        RECT 103.565 92.015 103.895 92.395 ;
        RECT 103.215 91.675 103.880 91.845 ;
        RECT 104.075 91.720 104.335 92.225 ;
        RECT 103.145 91.125 103.475 91.495 ;
        RECT 103.710 91.420 103.880 91.675 ;
        RECT 103.710 91.090 103.995 91.420 ;
        RECT 103.710 90.945 103.880 91.090 ;
        RECT 101.350 90.055 101.680 90.565 ;
        RECT 101.860 89.845 102.145 90.645 ;
        RECT 102.325 90.355 102.580 90.825 ;
        RECT 103.215 90.775 103.880 90.945 ;
        RECT 104.165 90.920 104.335 91.720 ;
        RECT 104.505 91.625 108.015 92.395 ;
        RECT 108.645 91.670 108.935 92.395 ;
        RECT 109.110 91.655 109.365 92.225 ;
        RECT 109.535 91.995 109.865 92.395 ;
        RECT 110.290 91.860 110.820 92.225 ;
        RECT 110.290 91.825 110.465 91.860 ;
        RECT 109.535 91.655 110.465 91.825 ;
        RECT 111.010 91.715 111.285 92.225 ;
        RECT 104.505 91.105 106.155 91.625 ;
        RECT 106.325 90.935 108.015 91.455 ;
        RECT 102.325 90.185 102.665 90.355 ;
        RECT 102.325 90.155 102.580 90.185 ;
        RECT 103.215 90.015 103.385 90.775 ;
        RECT 103.565 89.845 103.895 90.605 ;
        RECT 104.065 90.015 104.335 90.920 ;
        RECT 104.505 89.845 108.015 90.935 ;
        RECT 108.645 89.845 108.935 91.010 ;
        RECT 109.110 90.985 109.280 91.655 ;
        RECT 109.535 91.485 109.705 91.655 ;
        RECT 109.450 91.155 109.705 91.485 ;
        RECT 109.930 91.155 110.125 91.485 ;
        RECT 109.110 90.015 109.445 90.985 ;
        RECT 109.615 89.845 109.785 90.985 ;
        RECT 109.955 90.185 110.125 91.155 ;
        RECT 110.295 90.525 110.465 91.655 ;
        RECT 110.635 90.865 110.805 91.665 ;
        RECT 111.005 91.545 111.285 91.715 ;
        RECT 111.010 91.065 111.285 91.545 ;
        RECT 111.455 90.865 111.645 92.225 ;
        RECT 111.825 91.860 112.335 92.395 ;
        RECT 112.555 91.585 112.800 92.190 ;
        RECT 113.245 91.625 116.755 92.395 ;
        RECT 117.385 91.645 118.595 92.395 ;
        RECT 111.845 91.415 113.075 91.585 ;
        RECT 110.635 90.695 111.645 90.865 ;
        RECT 111.815 90.850 112.565 91.040 ;
        RECT 110.295 90.355 111.420 90.525 ;
        RECT 111.815 90.185 111.985 90.850 ;
        RECT 112.735 90.605 113.075 91.415 ;
        RECT 113.245 91.105 114.895 91.625 ;
        RECT 115.065 90.935 116.755 91.455 ;
        RECT 109.955 90.015 111.985 90.185 ;
        RECT 112.155 89.845 112.325 90.605 ;
        RECT 112.560 90.195 113.075 90.605 ;
        RECT 113.245 89.845 116.755 90.935 ;
        RECT 117.385 90.935 117.905 91.475 ;
        RECT 118.075 91.105 118.595 91.645 ;
        RECT 117.385 89.845 118.595 90.935 ;
        RECT 5.520 89.675 118.680 89.845 ;
        RECT 5.605 88.585 6.815 89.675 ;
        RECT 6.985 89.240 12.330 89.675 ;
        RECT 5.605 87.875 6.125 88.415 ;
        RECT 6.295 88.045 6.815 88.585 ;
        RECT 5.605 87.125 6.815 87.875 ;
        RECT 8.570 87.670 8.910 88.500 ;
        RECT 10.390 87.990 10.740 89.240 ;
        RECT 12.965 88.600 13.235 89.505 ;
        RECT 13.405 88.915 13.735 89.675 ;
        RECT 13.915 88.745 14.085 89.505 ;
        RECT 12.965 87.800 13.135 88.600 ;
        RECT 13.420 88.575 14.085 88.745 ;
        RECT 14.345 88.585 17.855 89.675 ;
        RECT 13.420 88.430 13.590 88.575 ;
        RECT 13.305 88.100 13.590 88.430 ;
        RECT 13.420 87.845 13.590 88.100 ;
        RECT 13.825 88.025 14.155 88.395 ;
        RECT 14.345 87.895 15.995 88.415 ;
        RECT 16.165 88.065 17.855 88.585 ;
        RECT 18.485 88.510 18.775 89.675 ;
        RECT 18.945 88.585 20.615 89.675 ;
        RECT 20.790 89.165 22.445 89.455 ;
        RECT 18.945 87.895 19.695 88.415 ;
        RECT 19.865 88.065 20.615 88.585 ;
        RECT 20.790 88.825 22.380 88.995 ;
        RECT 22.615 88.875 22.895 89.675 ;
        RECT 20.790 88.535 21.110 88.825 ;
        RECT 22.210 88.705 22.380 88.825 ;
        RECT 6.985 87.125 12.330 87.670 ;
        RECT 12.965 87.295 13.225 87.800 ;
        RECT 13.420 87.675 14.085 87.845 ;
        RECT 13.405 87.125 13.735 87.505 ;
        RECT 13.915 87.295 14.085 87.675 ;
        RECT 14.345 87.125 17.855 87.895 ;
        RECT 18.485 87.125 18.775 87.850 ;
        RECT 18.945 87.125 20.615 87.895 ;
        RECT 20.790 87.795 21.140 88.365 ;
        RECT 21.310 88.035 22.020 88.655 ;
        RECT 22.210 88.535 22.935 88.705 ;
        RECT 23.105 88.535 23.375 89.505 ;
        RECT 23.750 88.705 24.080 89.505 ;
        RECT 24.250 88.875 24.580 89.675 ;
        RECT 24.880 88.705 25.210 89.505 ;
        RECT 25.855 88.875 26.105 89.675 ;
        RECT 23.750 88.535 26.185 88.705 ;
        RECT 26.375 88.535 26.545 89.675 ;
        RECT 26.715 88.535 27.055 89.505 ;
        RECT 27.230 89.165 28.885 89.455 ;
        RECT 27.230 88.825 28.820 88.995 ;
        RECT 29.055 88.875 29.335 89.675 ;
        RECT 27.230 88.535 27.550 88.825 ;
        RECT 28.650 88.705 28.820 88.825 ;
        RECT 22.765 88.365 22.935 88.535 ;
        RECT 22.190 88.035 22.595 88.365 ;
        RECT 22.765 88.035 23.035 88.365 ;
        RECT 22.765 87.865 22.935 88.035 ;
        RECT 21.325 87.695 22.935 87.865 ;
        RECT 23.205 87.800 23.375 88.535 ;
        RECT 23.545 88.115 23.895 88.365 ;
        RECT 24.080 87.905 24.250 88.535 ;
        RECT 24.420 88.115 24.750 88.315 ;
        RECT 24.920 88.115 25.250 88.315 ;
        RECT 25.420 88.115 25.840 88.315 ;
        RECT 26.015 88.285 26.185 88.535 ;
        RECT 26.015 88.115 26.710 88.285 ;
        RECT 26.880 87.975 27.055 88.535 ;
        RECT 20.795 87.125 21.125 87.625 ;
        RECT 21.325 87.345 21.495 87.695 ;
        RECT 21.695 87.125 22.025 87.525 ;
        RECT 22.195 87.345 22.365 87.695 ;
        RECT 22.535 87.125 22.915 87.525 ;
        RECT 23.105 87.455 23.375 87.800 ;
        RECT 23.750 87.295 24.250 87.905 ;
        RECT 24.880 87.775 26.105 87.945 ;
        RECT 26.825 87.925 27.055 87.975 ;
        RECT 24.880 87.295 25.210 87.775 ;
        RECT 25.380 87.125 25.605 87.585 ;
        RECT 25.775 87.295 26.105 87.775 ;
        RECT 26.295 87.125 26.545 87.925 ;
        RECT 26.715 87.295 27.055 87.925 ;
        RECT 27.230 87.795 27.580 88.365 ;
        RECT 27.750 88.035 28.460 88.655 ;
        RECT 28.650 88.535 29.375 88.705 ;
        RECT 29.545 88.535 29.815 89.505 ;
        RECT 30.485 88.535 30.715 89.675 ;
        RECT 29.205 88.365 29.375 88.535 ;
        RECT 28.630 88.035 29.035 88.365 ;
        RECT 29.205 88.035 29.475 88.365 ;
        RECT 29.205 87.865 29.375 88.035 ;
        RECT 27.765 87.695 29.375 87.865 ;
        RECT 29.645 87.800 29.815 88.535 ;
        RECT 30.885 88.525 31.215 89.505 ;
        RECT 31.385 88.535 31.595 89.675 ;
        RECT 31.830 89.165 33.485 89.455 ;
        RECT 31.830 88.825 33.420 88.995 ;
        RECT 33.655 88.875 33.935 89.675 ;
        RECT 31.830 88.535 32.150 88.825 ;
        RECT 33.250 88.705 33.420 88.825 ;
        RECT 30.465 88.115 30.795 88.365 ;
        RECT 27.235 87.125 27.565 87.625 ;
        RECT 27.765 87.345 27.935 87.695 ;
        RECT 28.135 87.125 28.465 87.525 ;
        RECT 28.635 87.345 28.805 87.695 ;
        RECT 28.975 87.125 29.355 87.525 ;
        RECT 29.545 87.455 29.815 87.800 ;
        RECT 30.485 87.125 30.715 87.945 ;
        RECT 30.965 87.925 31.215 88.525 ;
        RECT 32.345 88.485 33.060 88.655 ;
        RECT 33.250 88.535 33.975 88.705 ;
        RECT 34.145 88.535 34.415 89.505 ;
        RECT 34.675 89.005 34.845 89.505 ;
        RECT 35.015 89.175 35.345 89.675 ;
        RECT 34.675 88.835 35.340 89.005 ;
        RECT 30.885 87.295 31.215 87.925 ;
        RECT 31.385 87.125 31.595 87.945 ;
        RECT 31.830 87.795 32.180 88.365 ;
        RECT 32.350 88.035 33.060 88.485 ;
        RECT 33.805 88.365 33.975 88.535 ;
        RECT 33.230 88.035 33.635 88.365 ;
        RECT 33.805 88.035 34.075 88.365 ;
        RECT 33.805 87.865 33.975 88.035 ;
        RECT 32.365 87.695 33.975 87.865 ;
        RECT 34.245 87.800 34.415 88.535 ;
        RECT 34.590 88.015 34.940 88.665 ;
        RECT 35.110 87.845 35.340 88.835 ;
        RECT 31.835 87.125 32.165 87.625 ;
        RECT 32.365 87.345 32.535 87.695 ;
        RECT 32.735 87.125 33.065 87.525 ;
        RECT 33.235 87.345 33.405 87.695 ;
        RECT 33.575 87.125 33.955 87.525 ;
        RECT 34.145 87.455 34.415 87.800 ;
        RECT 34.675 87.675 35.340 87.845 ;
        RECT 34.675 87.385 34.845 87.675 ;
        RECT 35.015 87.125 35.345 87.505 ;
        RECT 35.515 87.385 35.740 89.505 ;
        RECT 35.955 89.175 36.285 89.675 ;
        RECT 36.455 89.005 36.625 89.505 ;
        RECT 36.860 89.290 37.690 89.460 ;
        RECT 37.930 89.295 38.310 89.675 ;
        RECT 35.930 88.835 36.625 89.005 ;
        RECT 35.930 87.865 36.100 88.835 ;
        RECT 36.270 88.045 36.680 88.665 ;
        RECT 36.850 88.615 37.350 88.995 ;
        RECT 35.930 87.675 36.625 87.865 ;
        RECT 36.850 87.745 37.070 88.615 ;
        RECT 37.520 88.445 37.690 89.290 ;
        RECT 38.490 89.125 38.660 89.415 ;
        RECT 38.830 89.295 39.160 89.675 ;
        RECT 39.630 89.205 40.260 89.455 ;
        RECT 40.440 89.295 40.860 89.675 ;
        RECT 40.090 89.125 40.260 89.205 ;
        RECT 41.060 89.125 41.300 89.415 ;
        RECT 37.860 88.875 39.230 89.125 ;
        RECT 37.860 88.615 38.110 88.875 ;
        RECT 38.620 88.445 38.870 88.605 ;
        RECT 37.520 88.275 38.870 88.445 ;
        RECT 37.520 88.235 37.940 88.275 ;
        RECT 37.250 87.685 37.600 88.055 ;
        RECT 35.955 87.125 36.285 87.505 ;
        RECT 36.455 87.345 36.625 87.675 ;
        RECT 37.770 87.505 37.940 88.235 ;
        RECT 39.040 88.105 39.230 88.875 ;
        RECT 38.110 87.775 38.520 88.105 ;
        RECT 38.810 87.765 39.230 88.105 ;
        RECT 39.400 88.695 39.920 89.005 ;
        RECT 40.090 88.955 41.300 89.125 ;
        RECT 41.530 88.985 41.860 89.675 ;
        RECT 39.400 87.935 39.570 88.695 ;
        RECT 39.740 88.105 39.920 88.515 ;
        RECT 40.090 88.445 40.260 88.955 ;
        RECT 42.030 88.805 42.200 89.415 ;
        RECT 42.470 88.955 42.800 89.465 ;
        RECT 42.030 88.785 42.350 88.805 ;
        RECT 40.430 88.615 42.350 88.785 ;
        RECT 40.090 88.275 41.990 88.445 ;
        RECT 40.320 87.935 40.650 88.055 ;
        RECT 39.400 87.765 40.650 87.935 ;
        RECT 36.925 87.305 37.940 87.505 ;
        RECT 38.110 87.125 38.520 87.565 ;
        RECT 38.810 87.335 39.060 87.765 ;
        RECT 39.260 87.125 39.580 87.585 ;
        RECT 40.820 87.515 40.990 88.275 ;
        RECT 41.660 88.215 41.990 88.275 ;
        RECT 41.180 88.045 41.510 88.105 ;
        RECT 41.180 87.775 41.840 88.045 ;
        RECT 42.160 87.720 42.350 88.615 ;
        RECT 40.140 87.345 40.990 87.515 ;
        RECT 41.190 87.125 41.850 87.605 ;
        RECT 42.030 87.390 42.350 87.720 ;
        RECT 42.550 88.365 42.800 88.955 ;
        RECT 42.980 88.875 43.265 89.675 ;
        RECT 43.445 88.695 43.700 89.365 ;
        RECT 43.520 88.655 43.700 88.695 ;
        RECT 43.520 88.485 43.785 88.655 ;
        RECT 44.245 88.510 44.535 89.675 ;
        RECT 44.745 88.535 44.975 89.675 ;
        RECT 45.145 88.525 45.475 89.505 ;
        RECT 45.645 88.535 45.855 89.675 ;
        RECT 46.085 89.240 51.430 89.675 ;
        RECT 42.550 88.035 43.350 88.365 ;
        RECT 42.550 87.385 42.800 88.035 ;
        RECT 43.520 87.835 43.700 88.485 ;
        RECT 44.725 88.115 45.055 88.365 ;
        RECT 42.980 87.125 43.265 87.585 ;
        RECT 43.445 87.305 43.700 87.835 ;
        RECT 44.245 87.125 44.535 87.850 ;
        RECT 44.745 87.125 44.975 87.945 ;
        RECT 45.225 87.925 45.475 88.525 ;
        RECT 45.145 87.295 45.475 87.925 ;
        RECT 45.645 87.125 45.855 87.945 ;
        RECT 47.670 87.670 48.010 88.500 ;
        RECT 49.490 87.990 49.840 89.240 ;
        RECT 51.605 88.535 51.875 89.505 ;
        RECT 52.085 88.875 52.365 89.675 ;
        RECT 52.535 89.165 54.190 89.455 ;
        RECT 54.365 89.240 59.710 89.675 ;
        RECT 59.885 89.240 65.230 89.675 ;
        RECT 52.600 88.825 54.190 88.995 ;
        RECT 52.600 88.705 52.770 88.825 ;
        RECT 52.045 88.535 52.770 88.705 ;
        RECT 51.605 87.800 51.775 88.535 ;
        RECT 52.045 88.365 52.215 88.535 ;
        RECT 51.945 88.035 52.215 88.365 ;
        RECT 52.385 88.035 52.790 88.365 ;
        RECT 52.960 88.035 53.670 88.655 ;
        RECT 53.870 88.535 54.190 88.825 ;
        RECT 52.045 87.865 52.215 88.035 ;
        RECT 46.085 87.125 51.430 87.670 ;
        RECT 51.605 87.455 51.875 87.800 ;
        RECT 52.045 87.695 53.655 87.865 ;
        RECT 53.840 87.795 54.190 88.365 ;
        RECT 52.065 87.125 52.445 87.525 ;
        RECT 52.615 87.345 52.785 87.695 ;
        RECT 52.955 87.125 53.285 87.525 ;
        RECT 53.485 87.345 53.655 87.695 ;
        RECT 55.950 87.670 56.290 88.500 ;
        RECT 57.770 87.990 58.120 89.240 ;
        RECT 61.470 87.670 61.810 88.500 ;
        RECT 63.290 87.990 63.640 89.240 ;
        RECT 66.530 88.705 66.860 89.505 ;
        RECT 67.030 88.875 67.360 89.675 ;
        RECT 67.660 88.705 67.990 89.505 ;
        RECT 68.635 88.875 68.885 89.675 ;
        RECT 66.530 88.535 68.965 88.705 ;
        RECT 69.155 88.535 69.325 89.675 ;
        RECT 69.495 88.535 69.835 89.505 ;
        RECT 66.325 88.115 66.675 88.365 ;
        RECT 66.860 87.905 67.030 88.535 ;
        RECT 67.200 88.115 67.530 88.315 ;
        RECT 67.700 88.115 68.030 88.315 ;
        RECT 68.200 88.115 68.620 88.315 ;
        RECT 68.795 88.285 68.965 88.535 ;
        RECT 69.605 88.485 69.835 88.535 ;
        RECT 70.005 88.510 70.295 89.675 ;
        RECT 71.475 89.005 71.645 89.505 ;
        RECT 71.815 89.175 72.145 89.675 ;
        RECT 71.475 88.835 72.140 89.005 ;
        RECT 68.795 88.115 69.490 88.285 ;
        RECT 53.855 87.125 54.185 87.625 ;
        RECT 54.365 87.125 59.710 87.670 ;
        RECT 59.885 87.125 65.230 87.670 ;
        RECT 66.530 87.295 67.030 87.905 ;
        RECT 67.660 87.775 68.885 87.945 ;
        RECT 69.660 87.925 69.835 88.485 ;
        RECT 71.390 88.015 71.740 88.665 ;
        RECT 67.660 87.295 67.990 87.775 ;
        RECT 68.160 87.125 68.385 87.585 ;
        RECT 68.555 87.295 68.885 87.775 ;
        RECT 69.075 87.125 69.325 87.925 ;
        RECT 69.495 87.295 69.835 87.925 ;
        RECT 70.005 87.125 70.295 87.850 ;
        RECT 71.910 87.845 72.140 88.835 ;
        RECT 71.475 87.675 72.140 87.845 ;
        RECT 71.475 87.385 71.645 87.675 ;
        RECT 71.815 87.125 72.145 87.505 ;
        RECT 72.315 87.385 72.540 89.505 ;
        RECT 72.755 89.175 73.085 89.675 ;
        RECT 73.255 89.005 73.425 89.505 ;
        RECT 73.660 89.290 74.490 89.460 ;
        RECT 74.730 89.295 75.110 89.675 ;
        RECT 72.730 88.835 73.425 89.005 ;
        RECT 72.730 87.865 72.900 88.835 ;
        RECT 73.070 88.045 73.480 88.665 ;
        RECT 73.650 88.615 74.150 88.995 ;
        RECT 72.730 87.675 73.425 87.865 ;
        RECT 73.650 87.745 73.870 88.615 ;
        RECT 74.320 88.445 74.490 89.290 ;
        RECT 75.290 89.125 75.460 89.415 ;
        RECT 75.630 89.295 75.960 89.675 ;
        RECT 76.430 89.205 77.060 89.455 ;
        RECT 77.240 89.295 77.660 89.675 ;
        RECT 76.890 89.125 77.060 89.205 ;
        RECT 77.860 89.125 78.100 89.415 ;
        RECT 74.660 88.875 76.030 89.125 ;
        RECT 74.660 88.615 74.910 88.875 ;
        RECT 75.420 88.445 75.670 88.605 ;
        RECT 74.320 88.275 75.670 88.445 ;
        RECT 74.320 88.235 74.740 88.275 ;
        RECT 74.050 87.685 74.400 88.055 ;
        RECT 72.755 87.125 73.085 87.505 ;
        RECT 73.255 87.345 73.425 87.675 ;
        RECT 74.570 87.505 74.740 88.235 ;
        RECT 75.840 88.105 76.030 88.875 ;
        RECT 74.910 87.775 75.320 88.105 ;
        RECT 75.610 87.765 76.030 88.105 ;
        RECT 76.200 88.695 76.720 89.005 ;
        RECT 76.890 88.955 78.100 89.125 ;
        RECT 78.330 88.985 78.660 89.675 ;
        RECT 76.200 87.935 76.370 88.695 ;
        RECT 76.540 88.105 76.720 88.515 ;
        RECT 76.890 88.445 77.060 88.955 ;
        RECT 78.830 88.805 79.000 89.415 ;
        RECT 79.270 88.955 79.600 89.465 ;
        RECT 78.830 88.785 79.150 88.805 ;
        RECT 77.230 88.615 79.150 88.785 ;
        RECT 76.890 88.275 78.790 88.445 ;
        RECT 77.120 87.935 77.450 88.055 ;
        RECT 76.200 87.765 77.450 87.935 ;
        RECT 73.725 87.305 74.740 87.505 ;
        RECT 74.910 87.125 75.320 87.565 ;
        RECT 75.610 87.335 75.860 87.765 ;
        RECT 76.060 87.125 76.380 87.585 ;
        RECT 77.620 87.515 77.790 88.275 ;
        RECT 78.460 88.215 78.790 88.275 ;
        RECT 77.980 88.045 78.310 88.105 ;
        RECT 77.980 87.775 78.640 88.045 ;
        RECT 78.960 87.720 79.150 88.615 ;
        RECT 76.940 87.345 77.790 87.515 ;
        RECT 77.990 87.125 78.650 87.605 ;
        RECT 78.830 87.390 79.150 87.720 ;
        RECT 79.350 88.365 79.600 88.955 ;
        RECT 79.780 88.875 80.065 89.675 ;
        RECT 80.245 88.695 80.500 89.365 ;
        RECT 79.350 88.035 80.150 88.365 ;
        RECT 79.350 87.385 79.600 88.035 ;
        RECT 80.320 87.835 80.500 88.695 ;
        RECT 81.250 88.705 81.580 89.505 ;
        RECT 81.750 88.875 82.080 89.675 ;
        RECT 82.380 88.705 82.710 89.505 ;
        RECT 83.355 88.875 83.605 89.675 ;
        RECT 81.250 88.535 83.685 88.705 ;
        RECT 83.875 88.535 84.045 89.675 ;
        RECT 84.215 88.535 84.555 89.505 ;
        RECT 84.930 88.705 85.260 89.505 ;
        RECT 85.430 88.875 85.760 89.675 ;
        RECT 86.060 88.705 86.390 89.505 ;
        RECT 87.035 88.875 87.285 89.675 ;
        RECT 84.930 88.535 87.365 88.705 ;
        RECT 87.555 88.535 87.725 89.675 ;
        RECT 87.895 88.535 88.235 89.505 ;
        RECT 81.045 88.115 81.395 88.365 ;
        RECT 81.580 87.905 81.750 88.535 ;
        RECT 81.920 88.115 82.250 88.315 ;
        RECT 82.420 88.115 82.750 88.315 ;
        RECT 82.920 88.115 83.340 88.315 ;
        RECT 83.515 88.285 83.685 88.535 ;
        RECT 83.515 88.115 84.210 88.285 ;
        RECT 84.380 87.975 84.555 88.535 ;
        RECT 84.725 88.115 85.075 88.365 ;
        RECT 80.245 87.635 80.500 87.835 ;
        RECT 79.780 87.125 80.065 87.585 ;
        RECT 80.245 87.465 80.585 87.635 ;
        RECT 80.245 87.305 80.500 87.465 ;
        RECT 81.250 87.295 81.750 87.905 ;
        RECT 82.380 87.775 83.605 87.945 ;
        RECT 84.325 87.925 84.555 87.975 ;
        RECT 82.380 87.295 82.710 87.775 ;
        RECT 82.880 87.125 83.105 87.585 ;
        RECT 83.275 87.295 83.605 87.775 ;
        RECT 83.795 87.125 84.045 87.925 ;
        RECT 84.215 87.295 84.555 87.925 ;
        RECT 85.260 87.905 85.430 88.535 ;
        RECT 85.600 88.115 85.930 88.315 ;
        RECT 86.100 88.115 86.430 88.315 ;
        RECT 86.600 88.115 87.020 88.315 ;
        RECT 87.195 88.285 87.365 88.535 ;
        RECT 88.005 88.485 88.235 88.535 ;
        RECT 87.195 88.115 87.890 88.285 ;
        RECT 84.930 87.295 85.430 87.905 ;
        RECT 86.060 87.775 87.285 87.945 ;
        RECT 88.060 87.925 88.235 88.485 ;
        RECT 86.060 87.295 86.390 87.775 ;
        RECT 86.560 87.125 86.785 87.585 ;
        RECT 86.955 87.295 87.285 87.775 ;
        RECT 87.475 87.125 87.725 87.925 ;
        RECT 87.895 87.295 88.235 87.925 ;
        RECT 88.405 88.535 88.675 89.505 ;
        RECT 88.885 88.875 89.165 89.675 ;
        RECT 89.335 89.165 90.990 89.455 ;
        RECT 89.400 88.825 90.990 88.995 ;
        RECT 89.400 88.705 89.570 88.825 ;
        RECT 88.845 88.535 89.570 88.705 ;
        RECT 88.405 87.800 88.575 88.535 ;
        RECT 88.845 88.365 89.015 88.535 ;
        RECT 88.745 88.035 89.015 88.365 ;
        RECT 89.185 88.035 89.590 88.365 ;
        RECT 89.760 88.035 90.470 88.655 ;
        RECT 90.670 88.535 90.990 88.825 ;
        RECT 91.165 88.535 91.435 89.505 ;
        RECT 91.645 88.875 91.925 89.675 ;
        RECT 92.095 89.165 93.750 89.455 ;
        RECT 92.160 88.825 93.750 88.995 ;
        RECT 92.160 88.705 92.330 88.825 ;
        RECT 91.605 88.535 92.330 88.705 ;
        RECT 88.845 87.865 89.015 88.035 ;
        RECT 88.405 87.455 88.675 87.800 ;
        RECT 88.845 87.695 90.455 87.865 ;
        RECT 90.640 87.795 90.990 88.365 ;
        RECT 91.165 87.800 91.335 88.535 ;
        RECT 91.605 88.365 91.775 88.535 ;
        RECT 91.505 88.035 91.775 88.365 ;
        RECT 91.945 88.035 92.350 88.365 ;
        RECT 92.520 88.035 93.230 88.655 ;
        RECT 93.430 88.535 93.750 88.825 ;
        RECT 93.925 88.585 95.595 89.675 ;
        RECT 91.605 87.865 91.775 88.035 ;
        RECT 88.865 87.125 89.245 87.525 ;
        RECT 89.415 87.345 89.585 87.695 ;
        RECT 89.755 87.125 90.085 87.525 ;
        RECT 90.285 87.345 90.455 87.695 ;
        RECT 90.655 87.125 90.985 87.625 ;
        RECT 91.165 87.455 91.435 87.800 ;
        RECT 91.605 87.695 93.215 87.865 ;
        RECT 93.400 87.795 93.750 88.365 ;
        RECT 93.925 87.895 94.675 88.415 ;
        RECT 94.845 88.065 95.595 88.585 ;
        RECT 95.765 88.510 96.055 89.675 ;
        RECT 96.230 88.535 96.565 89.505 ;
        RECT 96.735 88.535 96.905 89.675 ;
        RECT 97.075 89.335 99.105 89.505 ;
        RECT 91.625 87.125 92.005 87.525 ;
        RECT 92.175 87.345 92.345 87.695 ;
        RECT 92.515 87.125 92.845 87.525 ;
        RECT 93.045 87.345 93.215 87.695 ;
        RECT 93.415 87.125 93.745 87.625 ;
        RECT 93.925 87.125 95.595 87.895 ;
        RECT 96.230 87.865 96.400 88.535 ;
        RECT 97.075 88.365 97.245 89.335 ;
        RECT 96.570 88.035 96.825 88.365 ;
        RECT 97.050 88.035 97.245 88.365 ;
        RECT 97.415 88.995 98.540 89.165 ;
        RECT 96.655 87.865 96.825 88.035 ;
        RECT 97.415 87.865 97.585 88.995 ;
        RECT 95.765 87.125 96.055 87.850 ;
        RECT 96.230 87.295 96.485 87.865 ;
        RECT 96.655 87.695 97.585 87.865 ;
        RECT 97.755 88.655 98.765 88.825 ;
        RECT 97.755 87.855 97.925 88.655 ;
        RECT 98.130 88.315 98.405 88.455 ;
        RECT 98.125 88.145 98.405 88.315 ;
        RECT 97.410 87.660 97.585 87.695 ;
        RECT 96.655 87.125 96.985 87.525 ;
        RECT 97.410 87.295 97.940 87.660 ;
        RECT 98.130 87.295 98.405 88.145 ;
        RECT 98.575 87.295 98.765 88.655 ;
        RECT 98.935 88.670 99.105 89.335 ;
        RECT 99.275 88.915 99.445 89.675 ;
        RECT 99.680 88.915 100.195 89.325 ;
        RECT 98.935 88.480 99.685 88.670 ;
        RECT 99.855 88.105 100.195 88.915 ;
        RECT 98.965 87.935 100.195 88.105 ;
        RECT 100.365 88.955 100.825 89.505 ;
        RECT 101.015 88.955 101.345 89.675 ;
        RECT 98.945 87.125 99.455 87.660 ;
        RECT 99.675 87.330 99.920 87.935 ;
        RECT 100.365 87.585 100.615 88.955 ;
        RECT 101.545 88.785 101.845 89.335 ;
        RECT 102.015 89.005 102.295 89.675 ;
        RECT 103.215 89.005 103.385 89.505 ;
        RECT 103.555 89.175 103.885 89.675 ;
        RECT 103.215 88.835 103.880 89.005 ;
        RECT 100.905 88.615 101.845 88.785 ;
        RECT 100.905 88.365 101.075 88.615 ;
        RECT 102.215 88.365 102.480 88.725 ;
        RECT 100.785 88.035 101.075 88.365 ;
        RECT 101.245 88.115 101.585 88.365 ;
        RECT 101.805 88.115 102.480 88.365 ;
        RECT 100.905 87.945 101.075 88.035 ;
        RECT 103.130 88.015 103.480 88.665 ;
        RECT 100.905 87.755 102.295 87.945 ;
        RECT 103.650 87.845 103.880 88.835 ;
        RECT 100.365 87.295 100.925 87.585 ;
        RECT 101.095 87.125 101.345 87.585 ;
        RECT 101.965 87.395 102.295 87.755 ;
        RECT 103.215 87.675 103.880 87.845 ;
        RECT 103.215 87.385 103.385 87.675 ;
        RECT 103.555 87.125 103.885 87.505 ;
        RECT 104.055 87.385 104.280 89.505 ;
        RECT 104.495 89.175 104.825 89.675 ;
        RECT 104.995 89.005 105.165 89.505 ;
        RECT 105.400 89.290 106.230 89.460 ;
        RECT 106.470 89.295 106.850 89.675 ;
        RECT 104.470 88.835 105.165 89.005 ;
        RECT 104.470 87.865 104.640 88.835 ;
        RECT 104.810 88.045 105.220 88.665 ;
        RECT 105.390 88.615 105.890 88.995 ;
        RECT 104.470 87.675 105.165 87.865 ;
        RECT 105.390 87.745 105.610 88.615 ;
        RECT 106.060 88.445 106.230 89.290 ;
        RECT 107.030 89.125 107.200 89.415 ;
        RECT 107.370 89.295 107.700 89.675 ;
        RECT 108.170 89.205 108.800 89.455 ;
        RECT 108.980 89.295 109.400 89.675 ;
        RECT 108.630 89.125 108.800 89.205 ;
        RECT 109.600 89.125 109.840 89.415 ;
        RECT 106.400 88.875 107.770 89.125 ;
        RECT 106.400 88.615 106.650 88.875 ;
        RECT 107.160 88.445 107.410 88.605 ;
        RECT 106.060 88.275 107.410 88.445 ;
        RECT 106.060 88.235 106.480 88.275 ;
        RECT 105.790 87.685 106.140 88.055 ;
        RECT 104.495 87.125 104.825 87.505 ;
        RECT 104.995 87.345 105.165 87.675 ;
        RECT 106.310 87.505 106.480 88.235 ;
        RECT 107.580 88.105 107.770 88.875 ;
        RECT 106.650 87.775 107.060 88.105 ;
        RECT 107.350 87.765 107.770 88.105 ;
        RECT 107.940 88.695 108.460 89.005 ;
        RECT 108.630 88.955 109.840 89.125 ;
        RECT 110.070 88.985 110.400 89.675 ;
        RECT 107.940 87.935 108.110 88.695 ;
        RECT 108.280 88.105 108.460 88.515 ;
        RECT 108.630 88.445 108.800 88.955 ;
        RECT 110.570 88.805 110.740 89.415 ;
        RECT 111.010 88.955 111.340 89.465 ;
        RECT 110.570 88.785 110.890 88.805 ;
        RECT 108.970 88.615 110.890 88.785 ;
        RECT 108.630 88.275 110.530 88.445 ;
        RECT 108.860 87.935 109.190 88.055 ;
        RECT 107.940 87.765 109.190 87.935 ;
        RECT 105.465 87.305 106.480 87.505 ;
        RECT 106.650 87.125 107.060 87.565 ;
        RECT 107.350 87.335 107.600 87.765 ;
        RECT 107.800 87.125 108.120 87.585 ;
        RECT 109.360 87.515 109.530 88.275 ;
        RECT 110.200 88.215 110.530 88.275 ;
        RECT 109.720 88.045 110.050 88.105 ;
        RECT 109.720 87.775 110.380 88.045 ;
        RECT 110.700 87.720 110.890 88.615 ;
        RECT 108.680 87.345 109.530 87.515 ;
        RECT 109.730 87.125 110.390 87.605 ;
        RECT 110.570 87.390 110.890 87.720 ;
        RECT 111.090 88.365 111.340 88.955 ;
        RECT 111.520 88.875 111.805 89.675 ;
        RECT 111.985 88.695 112.240 89.365 ;
        RECT 111.090 88.035 111.890 88.365 ;
        RECT 111.090 87.385 111.340 88.035 ;
        RECT 112.060 87.835 112.240 88.695 ;
        RECT 112.845 88.535 113.055 89.675 ;
        RECT 113.225 88.525 113.555 89.505 ;
        RECT 113.725 88.535 113.955 89.675 ;
        RECT 114.165 88.600 114.435 89.505 ;
        RECT 114.605 88.915 114.935 89.675 ;
        RECT 115.115 88.745 115.285 89.505 ;
        RECT 111.985 87.635 112.240 87.835 ;
        RECT 111.520 87.125 111.805 87.585 ;
        RECT 111.985 87.465 112.325 87.635 ;
        RECT 111.985 87.305 112.240 87.465 ;
        RECT 112.845 87.125 113.055 87.945 ;
        RECT 113.225 87.925 113.475 88.525 ;
        RECT 113.645 88.115 113.975 88.365 ;
        RECT 113.225 87.295 113.555 87.925 ;
        RECT 113.725 87.125 113.955 87.945 ;
        RECT 114.165 87.800 114.335 88.600 ;
        RECT 114.620 88.575 115.285 88.745 ;
        RECT 114.620 88.430 114.790 88.575 ;
        RECT 115.585 88.535 115.815 89.675 ;
        RECT 115.985 88.525 116.315 89.505 ;
        RECT 116.485 88.535 116.695 89.675 ;
        RECT 117.385 88.585 118.595 89.675 ;
        RECT 114.505 88.100 114.790 88.430 ;
        RECT 114.620 87.845 114.790 88.100 ;
        RECT 115.025 88.025 115.355 88.395 ;
        RECT 115.565 88.115 115.895 88.365 ;
        RECT 114.165 87.295 114.425 87.800 ;
        RECT 114.620 87.675 115.285 87.845 ;
        RECT 114.605 87.125 114.935 87.505 ;
        RECT 115.115 87.295 115.285 87.675 ;
        RECT 115.585 87.125 115.815 87.945 ;
        RECT 116.065 87.925 116.315 88.525 ;
        RECT 117.385 88.045 117.905 88.585 ;
        RECT 115.985 87.295 116.315 87.925 ;
        RECT 116.485 87.125 116.695 87.945 ;
        RECT 118.075 87.875 118.595 88.415 ;
        RECT 117.385 87.125 118.595 87.875 ;
        RECT 5.520 86.955 118.680 87.125 ;
        RECT 5.605 86.205 6.815 86.955 ;
        RECT 5.605 85.665 6.125 86.205 ;
        RECT 6.985 86.185 8.655 86.955 ;
        RECT 8.825 86.280 9.085 86.785 ;
        RECT 9.265 86.575 9.595 86.955 ;
        RECT 9.775 86.405 9.945 86.785 ;
        RECT 6.295 85.495 6.815 86.035 ;
        RECT 6.985 85.665 7.735 86.185 ;
        RECT 7.905 85.495 8.655 86.015 ;
        RECT 5.605 84.405 6.815 85.495 ;
        RECT 6.985 84.405 8.655 85.495 ;
        RECT 8.825 85.480 8.995 86.280 ;
        RECT 9.280 86.235 9.945 86.405 ;
        RECT 10.295 86.405 10.465 86.695 ;
        RECT 10.635 86.575 10.965 86.955 ;
        RECT 10.295 86.235 10.960 86.405 ;
        RECT 9.280 85.980 9.450 86.235 ;
        RECT 9.165 85.650 9.450 85.980 ;
        RECT 9.685 85.685 10.015 86.055 ;
        RECT 9.280 85.505 9.450 85.650 ;
        RECT 8.825 84.575 9.095 85.480 ;
        RECT 9.280 85.335 9.945 85.505 ;
        RECT 10.210 85.415 10.560 86.065 ;
        RECT 9.265 84.405 9.595 85.165 ;
        RECT 9.775 84.575 9.945 85.335 ;
        RECT 10.730 85.245 10.960 86.235 ;
        RECT 10.295 85.075 10.960 85.245 ;
        RECT 10.295 84.575 10.465 85.075 ;
        RECT 10.635 84.405 10.965 84.905 ;
        RECT 11.135 84.575 11.360 86.695 ;
        RECT 11.575 86.575 11.905 86.955 ;
        RECT 12.075 86.405 12.245 86.735 ;
        RECT 12.545 86.575 13.560 86.775 ;
        RECT 11.550 86.215 12.245 86.405 ;
        RECT 11.550 85.245 11.720 86.215 ;
        RECT 11.890 85.415 12.300 86.035 ;
        RECT 12.470 85.465 12.690 86.335 ;
        RECT 12.870 86.025 13.220 86.395 ;
        RECT 13.390 85.845 13.560 86.575 ;
        RECT 13.730 86.515 14.140 86.955 ;
        RECT 14.430 86.315 14.680 86.745 ;
        RECT 14.880 86.495 15.200 86.955 ;
        RECT 15.760 86.565 16.610 86.735 ;
        RECT 13.730 85.975 14.140 86.305 ;
        RECT 14.430 85.975 14.850 86.315 ;
        RECT 13.140 85.805 13.560 85.845 ;
        RECT 13.140 85.635 14.490 85.805 ;
        RECT 11.550 85.075 12.245 85.245 ;
        RECT 12.470 85.085 12.970 85.465 ;
        RECT 11.575 84.405 11.905 84.905 ;
        RECT 12.075 84.575 12.245 85.075 ;
        RECT 13.140 84.790 13.310 85.635 ;
        RECT 14.240 85.475 14.490 85.635 ;
        RECT 13.480 85.205 13.730 85.465 ;
        RECT 14.660 85.205 14.850 85.975 ;
        RECT 13.480 84.955 14.850 85.205 ;
        RECT 15.020 86.145 16.270 86.315 ;
        RECT 15.020 85.385 15.190 86.145 ;
        RECT 15.940 86.025 16.270 86.145 ;
        RECT 15.360 85.565 15.540 85.975 ;
        RECT 16.440 85.805 16.610 86.565 ;
        RECT 16.810 86.475 17.470 86.955 ;
        RECT 17.650 86.360 17.970 86.690 ;
        RECT 16.800 86.035 17.460 86.305 ;
        RECT 16.800 85.975 17.130 86.035 ;
        RECT 17.280 85.805 17.610 85.865 ;
        RECT 15.710 85.635 17.610 85.805 ;
        RECT 15.020 85.075 15.540 85.385 ;
        RECT 15.710 85.125 15.880 85.635 ;
        RECT 17.780 85.465 17.970 86.360 ;
        RECT 16.050 85.295 17.970 85.465 ;
        RECT 17.650 85.275 17.970 85.295 ;
        RECT 18.170 86.045 18.420 86.695 ;
        RECT 18.600 86.495 18.885 86.955 ;
        RECT 19.065 86.275 19.320 86.775 ;
        RECT 19.065 86.245 19.405 86.275 ;
        RECT 19.140 86.105 19.405 86.245 ;
        RECT 19.870 86.215 20.125 86.785 ;
        RECT 20.295 86.555 20.625 86.955 ;
        RECT 21.050 86.420 21.580 86.785 ;
        RECT 21.050 86.385 21.225 86.420 ;
        RECT 20.295 86.215 21.225 86.385 ;
        RECT 18.170 85.715 18.970 86.045 ;
        RECT 15.710 84.955 16.920 85.125 ;
        RECT 12.480 84.620 13.310 84.790 ;
        RECT 13.550 84.405 13.930 84.785 ;
        RECT 14.110 84.665 14.280 84.955 ;
        RECT 15.710 84.875 15.880 84.955 ;
        RECT 14.450 84.405 14.780 84.785 ;
        RECT 15.250 84.625 15.880 84.875 ;
        RECT 16.060 84.405 16.480 84.785 ;
        RECT 16.680 84.665 16.920 84.955 ;
        RECT 17.150 84.405 17.480 85.095 ;
        RECT 17.650 84.665 17.820 85.275 ;
        RECT 18.170 85.125 18.420 85.715 ;
        RECT 19.140 85.385 19.320 86.105 ;
        RECT 18.090 84.615 18.420 85.125 ;
        RECT 18.600 84.405 18.885 85.205 ;
        RECT 19.065 84.715 19.320 85.385 ;
        RECT 19.870 85.545 20.040 86.215 ;
        RECT 20.295 86.045 20.465 86.215 ;
        RECT 20.210 85.715 20.465 86.045 ;
        RECT 20.690 85.715 20.885 86.045 ;
        RECT 19.870 84.575 20.205 85.545 ;
        RECT 20.375 84.405 20.545 85.545 ;
        RECT 20.715 84.745 20.885 85.715 ;
        RECT 21.055 85.085 21.225 86.215 ;
        RECT 21.395 85.425 21.565 86.225 ;
        RECT 21.770 85.935 22.045 86.785 ;
        RECT 21.765 85.765 22.045 85.935 ;
        RECT 21.770 85.625 22.045 85.765 ;
        RECT 22.215 85.425 22.405 86.785 ;
        RECT 22.585 86.420 23.095 86.955 ;
        RECT 23.315 86.145 23.560 86.750 ;
        RECT 25.015 86.405 25.185 86.785 ;
        RECT 25.365 86.575 25.695 86.955 ;
        RECT 25.015 86.235 25.680 86.405 ;
        RECT 25.875 86.280 26.135 86.785 ;
        RECT 22.605 85.975 23.835 86.145 ;
        RECT 21.395 85.255 22.405 85.425 ;
        RECT 22.575 85.410 23.325 85.600 ;
        RECT 21.055 84.915 22.180 85.085 ;
        RECT 22.575 84.745 22.745 85.410 ;
        RECT 23.495 85.165 23.835 85.975 ;
        RECT 24.945 85.685 25.275 86.055 ;
        RECT 25.510 85.980 25.680 86.235 ;
        RECT 25.510 85.650 25.795 85.980 ;
        RECT 25.510 85.505 25.680 85.650 ;
        RECT 20.715 84.575 22.745 84.745 ;
        RECT 22.915 84.405 23.085 85.165 ;
        RECT 23.320 84.755 23.835 85.165 ;
        RECT 25.015 85.335 25.680 85.505 ;
        RECT 25.965 85.480 26.135 86.280 ;
        RECT 25.015 84.575 25.185 85.335 ;
        RECT 25.365 84.405 25.695 85.165 ;
        RECT 25.865 84.575 26.135 85.480 ;
        RECT 26.310 86.215 26.565 86.785 ;
        RECT 26.735 86.555 27.065 86.955 ;
        RECT 27.490 86.420 28.020 86.785 ;
        RECT 27.490 86.385 27.665 86.420 ;
        RECT 26.735 86.215 27.665 86.385 ;
        RECT 26.310 85.545 26.480 86.215 ;
        RECT 26.735 86.045 26.905 86.215 ;
        RECT 26.650 85.715 26.905 86.045 ;
        RECT 27.130 85.715 27.325 86.045 ;
        RECT 26.310 84.575 26.645 85.545 ;
        RECT 26.815 84.405 26.985 85.545 ;
        RECT 27.155 84.745 27.325 85.715 ;
        RECT 27.495 85.085 27.665 86.215 ;
        RECT 27.835 85.425 28.005 86.225 ;
        RECT 28.210 85.935 28.485 86.785 ;
        RECT 28.205 85.765 28.485 85.935 ;
        RECT 28.210 85.625 28.485 85.765 ;
        RECT 28.655 85.425 28.845 86.785 ;
        RECT 29.025 86.420 29.535 86.955 ;
        RECT 29.755 86.145 30.000 86.750 ;
        RECT 31.365 86.230 31.655 86.955 ;
        RECT 31.825 86.155 32.165 86.785 ;
        RECT 32.335 86.155 32.585 86.955 ;
        RECT 32.775 86.305 33.105 86.785 ;
        RECT 33.275 86.495 33.500 86.955 ;
        RECT 33.670 86.305 34.000 86.785 ;
        RECT 29.045 85.975 30.275 86.145 ;
        RECT 27.835 85.255 28.845 85.425 ;
        RECT 29.015 85.410 29.765 85.600 ;
        RECT 27.495 84.915 28.620 85.085 ;
        RECT 29.015 84.745 29.185 85.410 ;
        RECT 29.935 85.165 30.275 85.975 ;
        RECT 27.155 84.575 29.185 84.745 ;
        RECT 29.355 84.405 29.525 85.165 ;
        RECT 29.760 84.755 30.275 85.165 ;
        RECT 31.365 84.405 31.655 85.570 ;
        RECT 31.825 85.545 32.000 86.155 ;
        RECT 32.775 86.135 34.000 86.305 ;
        RECT 34.630 86.175 35.130 86.785 ;
        RECT 32.170 85.795 32.865 85.965 ;
        RECT 32.695 85.545 32.865 85.795 ;
        RECT 33.040 85.765 33.460 85.965 ;
        RECT 33.630 85.765 33.960 85.965 ;
        RECT 34.130 85.765 34.460 85.965 ;
        RECT 34.630 85.545 34.800 86.175 ;
        RECT 36.240 86.145 36.485 86.750 ;
        RECT 36.705 86.420 37.215 86.955 ;
        RECT 35.965 85.975 37.195 86.145 ;
        RECT 34.985 85.715 35.335 85.965 ;
        RECT 31.825 84.575 32.165 85.545 ;
        RECT 32.335 84.405 32.505 85.545 ;
        RECT 32.695 85.375 35.130 85.545 ;
        RECT 32.775 84.405 33.025 85.205 ;
        RECT 33.670 84.575 34.000 85.375 ;
        RECT 34.300 84.405 34.630 85.205 ;
        RECT 34.800 84.575 35.130 85.375 ;
        RECT 35.965 85.165 36.305 85.975 ;
        RECT 36.475 85.410 37.225 85.600 ;
        RECT 35.965 84.755 36.480 85.165 ;
        RECT 36.715 84.405 36.885 85.165 ;
        RECT 37.055 84.745 37.225 85.410 ;
        RECT 37.395 85.425 37.585 86.785 ;
        RECT 37.755 86.615 38.030 86.785 ;
        RECT 37.755 86.445 38.035 86.615 ;
        RECT 37.755 85.625 38.030 86.445 ;
        RECT 38.220 86.420 38.750 86.785 ;
        RECT 39.175 86.555 39.505 86.955 ;
        RECT 38.575 86.385 38.750 86.420 ;
        RECT 38.235 85.425 38.405 86.225 ;
        RECT 37.395 85.255 38.405 85.425 ;
        RECT 38.575 86.215 39.505 86.385 ;
        RECT 39.675 86.215 39.930 86.785 ;
        RECT 40.195 86.405 40.365 86.695 ;
        RECT 40.535 86.575 40.865 86.955 ;
        RECT 40.195 86.235 40.860 86.405 ;
        RECT 38.575 85.085 38.745 86.215 ;
        RECT 39.335 86.045 39.505 86.215 ;
        RECT 37.620 84.915 38.745 85.085 ;
        RECT 38.915 85.715 39.110 86.045 ;
        RECT 39.335 85.715 39.590 86.045 ;
        RECT 38.915 84.745 39.085 85.715 ;
        RECT 39.760 85.545 39.930 86.215 ;
        RECT 37.055 84.575 39.085 84.745 ;
        RECT 39.255 84.405 39.425 85.545 ;
        RECT 39.595 84.575 39.930 85.545 ;
        RECT 40.110 85.415 40.460 86.065 ;
        RECT 40.630 85.245 40.860 86.235 ;
        RECT 40.195 85.075 40.860 85.245 ;
        RECT 40.195 84.575 40.365 85.075 ;
        RECT 40.535 84.405 40.865 84.905 ;
        RECT 41.035 84.575 41.260 86.695 ;
        RECT 41.475 86.575 41.805 86.955 ;
        RECT 41.975 86.405 42.145 86.735 ;
        RECT 42.445 86.575 43.460 86.775 ;
        RECT 41.450 86.215 42.145 86.405 ;
        RECT 41.450 85.245 41.620 86.215 ;
        RECT 41.790 85.415 42.200 86.035 ;
        RECT 42.370 85.465 42.590 86.335 ;
        RECT 42.770 86.025 43.120 86.395 ;
        RECT 43.290 85.845 43.460 86.575 ;
        RECT 43.630 86.515 44.040 86.955 ;
        RECT 44.330 86.315 44.580 86.745 ;
        RECT 44.780 86.495 45.100 86.955 ;
        RECT 45.660 86.565 46.510 86.735 ;
        RECT 43.630 85.975 44.040 86.305 ;
        RECT 44.330 85.975 44.750 86.315 ;
        RECT 43.040 85.805 43.460 85.845 ;
        RECT 43.040 85.635 44.390 85.805 ;
        RECT 41.450 85.075 42.145 85.245 ;
        RECT 42.370 85.085 42.870 85.465 ;
        RECT 41.475 84.405 41.805 84.905 ;
        RECT 41.975 84.575 42.145 85.075 ;
        RECT 43.040 84.790 43.210 85.635 ;
        RECT 44.140 85.475 44.390 85.635 ;
        RECT 43.380 85.205 43.630 85.465 ;
        RECT 44.560 85.205 44.750 85.975 ;
        RECT 43.380 84.955 44.750 85.205 ;
        RECT 44.920 86.145 46.170 86.315 ;
        RECT 44.920 85.385 45.090 86.145 ;
        RECT 45.840 86.025 46.170 86.145 ;
        RECT 45.260 85.565 45.440 85.975 ;
        RECT 46.340 85.805 46.510 86.565 ;
        RECT 46.710 86.475 47.370 86.955 ;
        RECT 47.550 86.360 47.870 86.690 ;
        RECT 46.700 86.035 47.360 86.305 ;
        RECT 46.700 85.975 47.030 86.035 ;
        RECT 47.180 85.805 47.510 85.865 ;
        RECT 45.610 85.635 47.510 85.805 ;
        RECT 44.920 85.075 45.440 85.385 ;
        RECT 45.610 85.125 45.780 85.635 ;
        RECT 47.680 85.465 47.870 86.360 ;
        RECT 45.950 85.295 47.870 85.465 ;
        RECT 47.550 85.275 47.870 85.295 ;
        RECT 48.070 86.045 48.320 86.695 ;
        RECT 48.500 86.495 48.785 86.955 ;
        RECT 48.965 86.245 49.220 86.775 ;
        RECT 48.070 85.715 48.870 86.045 ;
        RECT 45.610 84.955 46.820 85.125 ;
        RECT 42.380 84.620 43.210 84.790 ;
        RECT 43.450 84.405 43.830 84.785 ;
        RECT 44.010 84.665 44.180 84.955 ;
        RECT 45.610 84.875 45.780 84.955 ;
        RECT 44.350 84.405 44.680 84.785 ;
        RECT 45.150 84.625 45.780 84.875 ;
        RECT 45.960 84.405 46.380 84.785 ;
        RECT 46.580 84.665 46.820 84.955 ;
        RECT 47.050 84.405 47.380 85.095 ;
        RECT 47.550 84.665 47.720 85.275 ;
        RECT 48.070 85.125 48.320 85.715 ;
        RECT 49.040 85.385 49.220 86.245 ;
        RECT 49.970 86.175 50.470 86.785 ;
        RECT 49.765 85.715 50.115 85.965 ;
        RECT 50.300 85.545 50.470 86.175 ;
        RECT 51.100 86.305 51.430 86.785 ;
        RECT 51.600 86.495 51.825 86.955 ;
        RECT 51.995 86.305 52.325 86.785 ;
        RECT 51.100 86.135 52.325 86.305 ;
        RECT 52.515 86.155 52.765 86.955 ;
        RECT 52.935 86.155 53.275 86.785 ;
        RECT 53.455 86.455 53.785 86.955 ;
        RECT 53.985 86.385 54.155 86.735 ;
        RECT 54.355 86.555 54.685 86.955 ;
        RECT 54.855 86.385 55.025 86.735 ;
        RECT 55.195 86.555 55.575 86.955 ;
        RECT 50.640 85.765 50.970 85.965 ;
        RECT 51.140 85.765 51.470 85.965 ;
        RECT 51.640 85.765 52.060 85.965 ;
        RECT 52.235 85.795 52.930 85.965 ;
        RECT 52.235 85.545 52.405 85.795 ;
        RECT 53.100 85.545 53.275 86.155 ;
        RECT 53.450 85.715 53.800 86.285 ;
        RECT 53.985 86.215 55.595 86.385 ;
        RECT 55.765 86.280 56.035 86.625 ;
        RECT 55.425 86.045 55.595 86.215 ;
        RECT 47.990 84.615 48.320 85.125 ;
        RECT 48.500 84.405 48.785 85.205 ;
        RECT 48.965 84.915 49.220 85.385 ;
        RECT 49.970 85.375 52.405 85.545 ;
        RECT 48.965 84.745 49.305 84.915 ;
        RECT 48.965 84.715 49.220 84.745 ;
        RECT 49.970 84.575 50.300 85.375 ;
        RECT 50.470 84.405 50.800 85.205 ;
        RECT 51.100 84.575 51.430 85.375 ;
        RECT 52.075 84.405 52.325 85.205 ;
        RECT 52.595 84.405 52.765 85.545 ;
        RECT 52.935 84.575 53.275 85.545 ;
        RECT 53.450 85.255 53.770 85.545 ;
        RECT 53.970 85.425 54.680 86.045 ;
        RECT 54.850 85.715 55.255 86.045 ;
        RECT 55.425 85.715 55.695 86.045 ;
        RECT 55.425 85.545 55.595 85.715 ;
        RECT 55.865 85.545 56.035 86.280 ;
        RECT 57.125 86.230 57.415 86.955 ;
        RECT 57.585 86.185 61.095 86.955 ;
        RECT 61.725 86.455 61.985 86.785 ;
        RECT 62.155 86.595 62.485 86.955 ;
        RECT 62.740 86.575 64.040 86.785 ;
        RECT 57.585 85.665 59.235 86.185 ;
        RECT 54.870 85.375 55.595 85.545 ;
        RECT 54.870 85.255 55.040 85.375 ;
        RECT 53.450 85.085 55.040 85.255 ;
        RECT 53.450 84.625 55.105 84.915 ;
        RECT 55.275 84.405 55.555 85.205 ;
        RECT 55.765 84.575 56.035 85.545 ;
        RECT 57.125 84.405 57.415 85.570 ;
        RECT 59.405 85.495 61.095 86.015 ;
        RECT 57.585 84.405 61.095 85.495 ;
        RECT 61.725 85.255 61.895 86.455 ;
        RECT 62.740 86.425 62.910 86.575 ;
        RECT 62.155 86.300 62.910 86.425 ;
        RECT 62.065 86.255 62.910 86.300 ;
        RECT 62.065 86.135 62.335 86.255 ;
        RECT 62.065 85.560 62.235 86.135 ;
        RECT 62.465 85.695 62.875 86.000 ;
        RECT 63.165 85.965 63.375 86.365 ;
        RECT 63.045 85.755 63.375 85.965 ;
        RECT 63.620 85.965 63.840 86.365 ;
        RECT 64.315 86.190 64.770 86.955 ;
        RECT 64.945 86.215 65.330 86.785 ;
        RECT 65.500 86.495 65.825 86.955 ;
        RECT 66.345 86.325 66.625 86.785 ;
        RECT 63.620 85.755 64.095 85.965 ;
        RECT 64.285 85.765 64.775 85.965 ;
        RECT 62.065 85.525 62.265 85.560 ;
        RECT 63.595 85.525 64.770 85.585 ;
        RECT 62.065 85.415 64.770 85.525 ;
        RECT 62.125 85.355 63.925 85.415 ;
        RECT 63.595 85.325 63.925 85.355 ;
        RECT 61.725 84.575 61.985 85.255 ;
        RECT 62.155 84.405 62.405 85.185 ;
        RECT 62.655 85.155 63.490 85.165 ;
        RECT 64.080 85.155 64.265 85.245 ;
        RECT 62.655 84.955 64.265 85.155 ;
        RECT 62.655 84.575 62.905 84.955 ;
        RECT 64.035 84.915 64.265 84.955 ;
        RECT 64.515 84.795 64.770 85.415 ;
        RECT 63.075 84.405 63.430 84.785 ;
        RECT 64.435 84.575 64.770 84.795 ;
        RECT 64.945 85.545 65.225 86.215 ;
        RECT 65.500 86.155 66.625 86.325 ;
        RECT 65.500 86.045 65.950 86.155 ;
        RECT 65.395 85.715 65.950 86.045 ;
        RECT 66.815 85.985 67.215 86.785 ;
        RECT 67.615 86.495 67.885 86.955 ;
        RECT 68.055 86.325 68.340 86.785 ;
        RECT 64.945 84.575 65.330 85.545 ;
        RECT 65.500 85.255 65.950 85.715 ;
        RECT 66.120 85.425 67.215 85.985 ;
        RECT 65.500 85.035 66.625 85.255 ;
        RECT 65.500 84.405 65.825 84.865 ;
        RECT 66.345 84.575 66.625 85.035 ;
        RECT 66.815 84.575 67.215 85.425 ;
        RECT 67.385 86.155 68.340 86.325 ;
        RECT 68.830 86.175 69.330 86.785 ;
        RECT 67.385 85.255 67.595 86.155 ;
        RECT 67.765 85.425 68.455 85.985 ;
        RECT 68.625 85.715 68.975 85.965 ;
        RECT 69.160 85.545 69.330 86.175 ;
        RECT 69.960 86.305 70.290 86.785 ;
        RECT 70.460 86.495 70.685 86.955 ;
        RECT 70.855 86.305 71.185 86.785 ;
        RECT 69.960 86.135 71.185 86.305 ;
        RECT 71.375 86.155 71.625 86.955 ;
        RECT 71.795 86.155 72.135 86.785 ;
        RECT 69.500 85.765 69.830 85.965 ;
        RECT 70.000 85.765 70.330 85.965 ;
        RECT 70.500 85.765 70.920 85.965 ;
        RECT 71.095 85.795 71.790 85.965 ;
        RECT 71.095 85.545 71.265 85.795 ;
        RECT 71.960 85.545 72.135 86.155 ;
        RECT 72.305 86.185 73.975 86.955 ;
        RECT 74.145 86.280 74.405 86.785 ;
        RECT 74.585 86.575 74.915 86.955 ;
        RECT 75.095 86.405 75.265 86.785 ;
        RECT 72.305 85.665 73.055 86.185 ;
        RECT 68.830 85.375 71.265 85.545 ;
        RECT 67.385 85.035 68.340 85.255 ;
        RECT 67.615 84.405 67.885 84.865 ;
        RECT 68.055 84.575 68.340 85.035 ;
        RECT 68.830 84.575 69.160 85.375 ;
        RECT 69.330 84.405 69.660 85.205 ;
        RECT 69.960 84.575 70.290 85.375 ;
        RECT 70.935 84.405 71.185 85.205 ;
        RECT 71.455 84.405 71.625 85.545 ;
        RECT 71.795 84.575 72.135 85.545 ;
        RECT 73.225 85.495 73.975 86.015 ;
        RECT 72.305 84.405 73.975 85.495 ;
        RECT 74.145 85.480 74.315 86.280 ;
        RECT 74.600 86.235 75.265 86.405 ;
        RECT 74.600 85.980 74.770 86.235 ;
        RECT 75.990 86.215 76.245 86.785 ;
        RECT 76.415 86.555 76.745 86.955 ;
        RECT 77.170 86.420 77.700 86.785 ;
        RECT 77.170 86.385 77.345 86.420 ;
        RECT 76.415 86.215 77.345 86.385 ;
        RECT 74.485 85.650 74.770 85.980 ;
        RECT 75.005 85.685 75.335 86.055 ;
        RECT 74.600 85.505 74.770 85.650 ;
        RECT 75.990 85.545 76.160 86.215 ;
        RECT 76.415 86.045 76.585 86.215 ;
        RECT 76.330 85.715 76.585 86.045 ;
        RECT 76.810 85.715 77.005 86.045 ;
        RECT 74.145 84.575 74.415 85.480 ;
        RECT 74.600 85.335 75.265 85.505 ;
        RECT 74.585 84.405 74.915 85.165 ;
        RECT 75.095 84.575 75.265 85.335 ;
        RECT 75.990 84.575 76.325 85.545 ;
        RECT 76.495 84.405 76.665 85.545 ;
        RECT 76.835 84.745 77.005 85.715 ;
        RECT 77.175 85.085 77.345 86.215 ;
        RECT 77.515 85.425 77.685 86.225 ;
        RECT 77.890 85.935 78.165 86.785 ;
        RECT 77.885 85.765 78.165 85.935 ;
        RECT 77.890 85.625 78.165 85.765 ;
        RECT 78.335 85.425 78.525 86.785 ;
        RECT 78.705 86.420 79.215 86.955 ;
        RECT 79.435 86.145 79.680 86.750 ;
        RECT 80.125 86.185 82.715 86.955 ;
        RECT 82.885 86.230 83.175 86.955 ;
        RECT 78.725 85.975 79.955 86.145 ;
        RECT 77.515 85.255 78.525 85.425 ;
        RECT 78.695 85.410 79.445 85.600 ;
        RECT 77.175 84.915 78.300 85.085 ;
        RECT 78.695 84.745 78.865 85.410 ;
        RECT 79.615 85.165 79.955 85.975 ;
        RECT 80.125 85.665 81.335 86.185 ;
        RECT 83.550 86.175 84.050 86.785 ;
        RECT 81.505 85.495 82.715 86.015 ;
        RECT 83.345 85.715 83.695 85.965 ;
        RECT 76.835 84.575 78.865 84.745 ;
        RECT 79.035 84.405 79.205 85.165 ;
        RECT 79.440 84.755 79.955 85.165 ;
        RECT 80.125 84.405 82.715 85.495 ;
        RECT 82.885 84.405 83.175 85.570 ;
        RECT 83.880 85.545 84.050 86.175 ;
        RECT 84.680 86.305 85.010 86.785 ;
        RECT 85.180 86.495 85.405 86.955 ;
        RECT 85.575 86.305 85.905 86.785 ;
        RECT 84.680 86.135 85.905 86.305 ;
        RECT 86.095 86.155 86.345 86.955 ;
        RECT 86.515 86.155 86.855 86.785 ;
        RECT 87.035 86.455 87.365 86.955 ;
        RECT 87.565 86.385 87.735 86.735 ;
        RECT 87.935 86.555 88.265 86.955 ;
        RECT 88.435 86.385 88.605 86.735 ;
        RECT 88.775 86.555 89.155 86.955 ;
        RECT 86.625 86.105 86.855 86.155 ;
        RECT 84.220 85.765 84.550 85.965 ;
        RECT 84.720 85.765 85.050 85.965 ;
        RECT 85.220 85.765 85.640 85.965 ;
        RECT 85.815 85.795 86.510 85.965 ;
        RECT 85.815 85.545 85.985 85.795 ;
        RECT 86.680 85.545 86.855 86.105 ;
        RECT 87.030 85.715 87.380 86.285 ;
        RECT 87.565 86.215 89.175 86.385 ;
        RECT 89.345 86.280 89.615 86.625 ;
        RECT 89.005 86.045 89.175 86.215 ;
        RECT 87.550 85.595 88.260 86.045 ;
        RECT 88.430 85.715 88.835 86.045 ;
        RECT 89.005 85.715 89.275 86.045 ;
        RECT 83.550 85.375 85.985 85.545 ;
        RECT 83.550 84.575 83.880 85.375 ;
        RECT 84.050 84.405 84.380 85.205 ;
        RECT 84.680 84.575 85.010 85.375 ;
        RECT 85.655 84.405 85.905 85.205 ;
        RECT 86.175 84.405 86.345 85.545 ;
        RECT 86.515 84.575 86.855 85.545 ;
        RECT 87.030 85.255 87.350 85.545 ;
        RECT 87.545 85.425 88.260 85.595 ;
        RECT 89.005 85.545 89.175 85.715 ;
        RECT 89.445 85.545 89.615 86.280 ;
        RECT 89.785 86.185 92.375 86.955 ;
        RECT 93.015 86.455 93.345 86.955 ;
        RECT 93.545 86.385 93.715 86.735 ;
        RECT 93.915 86.555 94.245 86.955 ;
        RECT 94.415 86.385 94.585 86.735 ;
        RECT 94.755 86.555 95.135 86.955 ;
        RECT 89.785 85.665 90.995 86.185 ;
        RECT 88.450 85.375 89.175 85.545 ;
        RECT 88.450 85.255 88.620 85.375 ;
        RECT 87.030 85.085 88.620 85.255 ;
        RECT 87.030 84.625 88.685 84.915 ;
        RECT 88.855 84.405 89.135 85.205 ;
        RECT 89.345 84.575 89.615 85.545 ;
        RECT 91.165 85.495 92.375 86.015 ;
        RECT 93.010 85.715 93.360 86.285 ;
        RECT 93.545 86.215 95.155 86.385 ;
        RECT 95.325 86.280 95.595 86.625 ;
        RECT 95.775 86.455 96.105 86.955 ;
        RECT 96.305 86.385 96.475 86.735 ;
        RECT 96.675 86.555 97.005 86.955 ;
        RECT 97.175 86.385 97.345 86.735 ;
        RECT 97.515 86.555 97.895 86.955 ;
        RECT 94.985 86.045 95.155 86.215 ;
        RECT 89.785 84.405 92.375 85.495 ;
        RECT 93.010 85.255 93.330 85.545 ;
        RECT 93.530 85.425 94.240 86.045 ;
        RECT 94.410 85.715 94.815 86.045 ;
        RECT 94.985 85.715 95.255 86.045 ;
        RECT 94.985 85.545 95.155 85.715 ;
        RECT 95.425 85.545 95.595 86.280 ;
        RECT 95.770 85.715 96.120 86.285 ;
        RECT 96.305 86.215 97.915 86.385 ;
        RECT 98.085 86.280 98.355 86.625 ;
        RECT 97.745 86.045 97.915 86.215 ;
        RECT 94.430 85.375 95.155 85.545 ;
        RECT 94.430 85.255 94.600 85.375 ;
        RECT 93.010 85.085 94.600 85.255 ;
        RECT 93.010 84.625 94.665 84.915 ;
        RECT 94.835 84.405 95.115 85.205 ;
        RECT 95.325 84.575 95.595 85.545 ;
        RECT 95.770 85.255 96.090 85.545 ;
        RECT 96.290 85.425 97.000 86.045 ;
        RECT 97.170 85.715 97.575 86.045 ;
        RECT 97.745 85.715 98.015 86.045 ;
        RECT 97.745 85.545 97.915 85.715 ;
        RECT 98.185 85.545 98.355 86.280 ;
        RECT 97.190 85.375 97.915 85.545 ;
        RECT 97.190 85.255 97.360 85.375 ;
        RECT 95.770 85.085 97.360 85.255 ;
        RECT 95.770 84.625 97.425 84.915 ;
        RECT 97.595 84.405 97.875 85.205 ;
        RECT 98.085 84.575 98.355 85.545 ;
        RECT 98.525 86.495 99.085 86.785 ;
        RECT 99.255 86.495 99.505 86.955 ;
        RECT 98.525 85.125 98.775 86.495 ;
        RECT 100.125 86.325 100.455 86.685 ;
        RECT 99.065 86.135 100.455 86.325 ;
        RECT 101.100 86.145 101.345 86.750 ;
        RECT 101.565 86.420 102.075 86.955 ;
        RECT 99.065 86.045 99.235 86.135 ;
        RECT 98.945 85.715 99.235 86.045 ;
        RECT 100.825 85.975 102.055 86.145 ;
        RECT 99.405 85.715 99.745 85.965 ;
        RECT 99.965 85.715 100.640 85.965 ;
        RECT 99.065 85.465 99.235 85.715 ;
        RECT 99.065 85.295 100.005 85.465 ;
        RECT 100.375 85.355 100.640 85.715 ;
        RECT 98.525 84.575 98.985 85.125 ;
        RECT 99.175 84.405 99.505 85.125 ;
        RECT 99.705 84.745 100.005 85.295 ;
        RECT 100.825 85.165 101.165 85.975 ;
        RECT 101.335 85.410 102.085 85.600 ;
        RECT 100.175 84.405 100.455 85.075 ;
        RECT 100.825 84.755 101.340 85.165 ;
        RECT 101.575 84.405 101.745 85.165 ;
        RECT 101.915 84.745 102.085 85.410 ;
        RECT 102.255 85.425 102.445 86.785 ;
        RECT 102.615 86.275 102.890 86.785 ;
        RECT 103.080 86.420 103.610 86.785 ;
        RECT 104.035 86.555 104.365 86.955 ;
        RECT 103.435 86.385 103.610 86.420 ;
        RECT 102.615 86.105 102.895 86.275 ;
        RECT 102.615 85.625 102.890 86.105 ;
        RECT 103.095 85.425 103.265 86.225 ;
        RECT 102.255 85.255 103.265 85.425 ;
        RECT 103.435 86.215 104.365 86.385 ;
        RECT 104.535 86.215 104.790 86.785 ;
        RECT 103.435 85.085 103.605 86.215 ;
        RECT 104.195 86.045 104.365 86.215 ;
        RECT 102.480 84.915 103.605 85.085 ;
        RECT 103.775 85.715 103.970 86.045 ;
        RECT 104.195 85.715 104.450 86.045 ;
        RECT 103.775 84.745 103.945 85.715 ;
        RECT 104.620 85.545 104.790 86.215 ;
        RECT 104.965 86.185 108.475 86.955 ;
        RECT 108.645 86.230 108.935 86.955 ;
        RECT 104.965 85.665 106.615 86.185 ;
        RECT 109.380 86.145 109.625 86.750 ;
        RECT 109.845 86.420 110.355 86.955 ;
        RECT 101.915 84.575 103.945 84.745 ;
        RECT 104.115 84.405 104.285 85.545 ;
        RECT 104.455 84.575 104.790 85.545 ;
        RECT 106.785 85.495 108.475 86.015 ;
        RECT 109.105 85.975 110.335 86.145 ;
        RECT 104.965 84.405 108.475 85.495 ;
        RECT 108.645 84.405 108.935 85.570 ;
        RECT 109.105 85.165 109.445 85.975 ;
        RECT 109.615 85.410 110.365 85.600 ;
        RECT 109.105 84.755 109.620 85.165 ;
        RECT 109.855 84.405 110.025 85.165 ;
        RECT 110.195 84.745 110.365 85.410 ;
        RECT 110.535 85.425 110.725 86.785 ;
        RECT 110.895 85.935 111.170 86.785 ;
        RECT 111.360 86.420 111.890 86.785 ;
        RECT 112.315 86.555 112.645 86.955 ;
        RECT 111.715 86.385 111.890 86.420 ;
        RECT 110.895 85.765 111.175 85.935 ;
        RECT 110.895 85.625 111.170 85.765 ;
        RECT 111.375 85.425 111.545 86.225 ;
        RECT 110.535 85.255 111.545 85.425 ;
        RECT 111.715 86.215 112.645 86.385 ;
        RECT 112.815 86.215 113.070 86.785 ;
        RECT 111.715 85.085 111.885 86.215 ;
        RECT 112.475 86.045 112.645 86.215 ;
        RECT 110.760 84.915 111.885 85.085 ;
        RECT 112.055 85.715 112.250 86.045 ;
        RECT 112.475 85.715 112.730 86.045 ;
        RECT 112.055 84.745 112.225 85.715 ;
        RECT 112.900 85.545 113.070 86.215 ;
        RECT 113.245 86.185 116.755 86.955 ;
        RECT 117.385 86.205 118.595 86.955 ;
        RECT 113.245 85.665 114.895 86.185 ;
        RECT 110.195 84.575 112.225 84.745 ;
        RECT 112.395 84.405 112.565 85.545 ;
        RECT 112.735 84.575 113.070 85.545 ;
        RECT 115.065 85.495 116.755 86.015 ;
        RECT 113.245 84.405 116.755 85.495 ;
        RECT 117.385 85.495 117.905 86.035 ;
        RECT 118.075 85.665 118.595 86.205 ;
        RECT 117.385 84.405 118.595 85.495 ;
        RECT 5.520 84.235 118.680 84.405 ;
        RECT 5.605 83.145 6.815 84.235 ;
        RECT 7.075 83.565 7.245 84.065 ;
        RECT 7.415 83.735 7.745 84.235 ;
        RECT 7.075 83.395 7.740 83.565 ;
        RECT 5.605 82.435 6.125 82.975 ;
        RECT 6.295 82.605 6.815 83.145 ;
        RECT 6.990 82.575 7.340 83.225 ;
        RECT 5.605 81.685 6.815 82.435 ;
        RECT 7.510 82.405 7.740 83.395 ;
        RECT 7.075 82.235 7.740 82.405 ;
        RECT 7.075 81.945 7.245 82.235 ;
        RECT 7.415 81.685 7.745 82.065 ;
        RECT 7.915 81.945 8.140 84.065 ;
        RECT 8.355 83.735 8.685 84.235 ;
        RECT 8.855 83.565 9.025 84.065 ;
        RECT 9.260 83.850 10.090 84.020 ;
        RECT 10.330 83.855 10.710 84.235 ;
        RECT 8.330 83.395 9.025 83.565 ;
        RECT 8.330 82.425 8.500 83.395 ;
        RECT 8.670 82.605 9.080 83.225 ;
        RECT 9.250 83.175 9.750 83.555 ;
        RECT 8.330 82.235 9.025 82.425 ;
        RECT 9.250 82.305 9.470 83.175 ;
        RECT 9.920 83.005 10.090 83.850 ;
        RECT 10.890 83.685 11.060 83.975 ;
        RECT 11.230 83.855 11.560 84.235 ;
        RECT 12.030 83.765 12.660 84.015 ;
        RECT 12.840 83.855 13.260 84.235 ;
        RECT 12.490 83.685 12.660 83.765 ;
        RECT 13.460 83.685 13.700 83.975 ;
        RECT 10.260 83.435 11.630 83.685 ;
        RECT 10.260 83.175 10.510 83.435 ;
        RECT 11.020 83.005 11.270 83.165 ;
        RECT 9.920 82.835 11.270 83.005 ;
        RECT 9.920 82.795 10.340 82.835 ;
        RECT 9.650 82.245 10.000 82.615 ;
        RECT 8.355 81.685 8.685 82.065 ;
        RECT 8.855 81.905 9.025 82.235 ;
        RECT 10.170 82.065 10.340 82.795 ;
        RECT 11.440 82.665 11.630 83.435 ;
        RECT 10.510 82.335 10.920 82.665 ;
        RECT 11.210 82.325 11.630 82.665 ;
        RECT 11.800 83.255 12.320 83.565 ;
        RECT 12.490 83.515 13.700 83.685 ;
        RECT 13.930 83.545 14.260 84.235 ;
        RECT 11.800 82.495 11.970 83.255 ;
        RECT 12.140 82.665 12.320 83.075 ;
        RECT 12.490 83.005 12.660 83.515 ;
        RECT 14.430 83.365 14.600 83.975 ;
        RECT 14.870 83.515 15.200 84.025 ;
        RECT 14.430 83.345 14.750 83.365 ;
        RECT 12.830 83.175 14.750 83.345 ;
        RECT 12.490 82.835 14.390 83.005 ;
        RECT 12.720 82.495 13.050 82.615 ;
        RECT 11.800 82.325 13.050 82.495 ;
        RECT 9.325 81.865 10.340 82.065 ;
        RECT 10.510 81.685 10.920 82.125 ;
        RECT 11.210 81.895 11.460 82.325 ;
        RECT 11.660 81.685 11.980 82.145 ;
        RECT 13.220 82.075 13.390 82.835 ;
        RECT 14.060 82.775 14.390 82.835 ;
        RECT 13.580 82.605 13.910 82.665 ;
        RECT 13.580 82.335 14.240 82.605 ;
        RECT 14.560 82.280 14.750 83.175 ;
        RECT 12.540 81.905 13.390 82.075 ;
        RECT 13.590 81.685 14.250 82.165 ;
        RECT 14.430 81.950 14.750 82.280 ;
        RECT 14.950 82.925 15.200 83.515 ;
        RECT 15.380 83.435 15.665 84.235 ;
        RECT 15.845 83.255 16.100 83.925 ;
        RECT 14.950 82.595 15.750 82.925 ;
        RECT 14.950 81.945 15.200 82.595 ;
        RECT 15.920 82.535 16.100 83.255 ;
        RECT 16.705 83.095 16.915 84.235 ;
        RECT 17.085 83.085 17.415 84.065 ;
        RECT 17.585 83.095 17.815 84.235 ;
        RECT 15.920 82.395 16.185 82.535 ;
        RECT 15.845 82.365 16.185 82.395 ;
        RECT 15.380 81.685 15.665 82.145 ;
        RECT 15.845 81.865 16.100 82.365 ;
        RECT 16.705 81.685 16.915 82.505 ;
        RECT 17.085 82.485 17.335 83.085 ;
        RECT 18.485 83.070 18.775 84.235 ;
        RECT 19.865 83.095 20.205 84.065 ;
        RECT 20.375 83.095 20.545 84.235 ;
        RECT 20.815 83.435 21.065 84.235 ;
        RECT 21.710 83.265 22.040 84.065 ;
        RECT 22.340 83.435 22.670 84.235 ;
        RECT 22.840 83.265 23.170 84.065 ;
        RECT 20.735 83.095 23.170 83.265 ;
        RECT 23.545 83.145 25.215 84.235 ;
        RECT 25.935 83.565 26.105 84.065 ;
        RECT 26.275 83.735 26.605 84.235 ;
        RECT 25.935 83.395 26.600 83.565 ;
        RECT 17.505 82.675 17.835 82.925 ;
        RECT 19.865 82.535 20.040 83.095 ;
        RECT 20.735 82.845 20.905 83.095 ;
        RECT 20.210 82.675 20.905 82.845 ;
        RECT 21.080 82.675 21.500 82.875 ;
        RECT 21.670 82.675 22.000 82.875 ;
        RECT 22.170 82.675 22.500 82.875 ;
        RECT 17.085 81.855 17.415 82.485 ;
        RECT 17.585 81.685 17.815 82.505 ;
        RECT 19.865 82.485 20.095 82.535 ;
        RECT 18.485 81.685 18.775 82.410 ;
        RECT 19.865 81.855 20.205 82.485 ;
        RECT 20.375 81.685 20.625 82.485 ;
        RECT 20.815 82.335 22.040 82.505 ;
        RECT 20.815 81.855 21.145 82.335 ;
        RECT 21.315 81.685 21.540 82.145 ;
        RECT 21.710 81.855 22.040 82.335 ;
        RECT 22.670 82.465 22.840 83.095 ;
        RECT 23.025 82.675 23.375 82.925 ;
        RECT 22.670 81.855 23.170 82.465 ;
        RECT 23.545 82.455 24.295 82.975 ;
        RECT 24.465 82.625 25.215 83.145 ;
        RECT 25.850 82.575 26.200 83.225 ;
        RECT 23.545 81.685 25.215 82.455 ;
        RECT 26.370 82.405 26.600 83.395 ;
        RECT 25.935 82.235 26.600 82.405 ;
        RECT 25.935 81.945 26.105 82.235 ;
        RECT 26.275 81.685 26.605 82.065 ;
        RECT 26.775 81.945 27.000 84.065 ;
        RECT 27.215 83.735 27.545 84.235 ;
        RECT 27.715 83.565 27.885 84.065 ;
        RECT 28.120 83.850 28.950 84.020 ;
        RECT 29.190 83.855 29.570 84.235 ;
        RECT 27.190 83.395 27.885 83.565 ;
        RECT 27.190 82.425 27.360 83.395 ;
        RECT 27.530 82.605 27.940 83.225 ;
        RECT 28.110 83.175 28.610 83.555 ;
        RECT 27.190 82.235 27.885 82.425 ;
        RECT 28.110 82.305 28.330 83.175 ;
        RECT 28.780 83.005 28.950 83.850 ;
        RECT 29.750 83.685 29.920 83.975 ;
        RECT 30.090 83.855 30.420 84.235 ;
        RECT 30.890 83.765 31.520 84.015 ;
        RECT 31.700 83.855 32.120 84.235 ;
        RECT 31.350 83.685 31.520 83.765 ;
        RECT 32.320 83.685 32.560 83.975 ;
        RECT 29.120 83.435 30.490 83.685 ;
        RECT 29.120 83.175 29.370 83.435 ;
        RECT 29.880 83.005 30.130 83.165 ;
        RECT 28.780 82.835 30.130 83.005 ;
        RECT 28.780 82.795 29.200 82.835 ;
        RECT 28.510 82.245 28.860 82.615 ;
        RECT 27.215 81.685 27.545 82.065 ;
        RECT 27.715 81.905 27.885 82.235 ;
        RECT 29.030 82.065 29.200 82.795 ;
        RECT 30.300 82.665 30.490 83.435 ;
        RECT 29.370 82.335 29.780 82.665 ;
        RECT 30.070 82.325 30.490 82.665 ;
        RECT 30.660 83.255 31.180 83.565 ;
        RECT 31.350 83.515 32.560 83.685 ;
        RECT 32.790 83.545 33.120 84.235 ;
        RECT 30.660 82.495 30.830 83.255 ;
        RECT 31.000 82.665 31.180 83.075 ;
        RECT 31.350 83.005 31.520 83.515 ;
        RECT 33.290 83.365 33.460 83.975 ;
        RECT 33.730 83.515 34.060 84.025 ;
        RECT 33.290 83.345 33.610 83.365 ;
        RECT 31.690 83.175 33.610 83.345 ;
        RECT 31.350 82.835 33.250 83.005 ;
        RECT 31.580 82.495 31.910 82.615 ;
        RECT 30.660 82.325 31.910 82.495 ;
        RECT 28.185 81.865 29.200 82.065 ;
        RECT 29.370 81.685 29.780 82.125 ;
        RECT 30.070 81.895 30.320 82.325 ;
        RECT 30.520 81.685 30.840 82.145 ;
        RECT 32.080 82.075 32.250 82.835 ;
        RECT 32.920 82.775 33.250 82.835 ;
        RECT 32.440 82.605 32.770 82.665 ;
        RECT 32.440 82.335 33.100 82.605 ;
        RECT 33.420 82.280 33.610 83.175 ;
        RECT 31.400 81.905 32.250 82.075 ;
        RECT 32.450 81.685 33.110 82.165 ;
        RECT 33.290 81.950 33.610 82.280 ;
        RECT 33.810 82.925 34.060 83.515 ;
        RECT 34.240 83.435 34.525 84.235 ;
        RECT 34.705 83.255 34.960 83.925 ;
        RECT 35.505 83.800 40.850 84.235 ;
        RECT 34.780 83.215 34.960 83.255 ;
        RECT 34.780 83.045 35.045 83.215 ;
        RECT 33.810 82.595 34.610 82.925 ;
        RECT 33.810 81.945 34.060 82.595 ;
        RECT 34.780 82.395 34.960 83.045 ;
        RECT 34.240 81.685 34.525 82.145 ;
        RECT 34.705 81.865 34.960 82.395 ;
        RECT 37.090 82.230 37.430 83.060 ;
        RECT 38.910 82.550 39.260 83.800 ;
        RECT 41.025 83.145 42.695 84.235 ;
        RECT 41.025 82.455 41.775 82.975 ;
        RECT 41.945 82.625 42.695 83.145 ;
        RECT 42.865 83.160 43.135 84.065 ;
        RECT 43.305 83.475 43.635 84.235 ;
        RECT 43.815 83.305 43.985 84.065 ;
        RECT 35.505 81.685 40.850 82.230 ;
        RECT 41.025 81.685 42.695 82.455 ;
        RECT 42.865 82.360 43.035 83.160 ;
        RECT 43.320 83.135 43.985 83.305 ;
        RECT 43.320 82.990 43.490 83.135 ;
        RECT 44.245 83.070 44.535 84.235 ;
        RECT 44.710 83.095 45.045 84.065 ;
        RECT 45.215 83.095 45.385 84.235 ;
        RECT 45.555 83.895 47.585 84.065 ;
        RECT 43.205 82.660 43.490 82.990 ;
        RECT 43.320 82.405 43.490 82.660 ;
        RECT 43.725 82.585 44.055 82.955 ;
        RECT 44.710 82.425 44.880 83.095 ;
        RECT 45.555 82.925 45.725 83.895 ;
        RECT 45.050 82.595 45.305 82.925 ;
        RECT 45.530 82.595 45.725 82.925 ;
        RECT 45.895 83.555 47.020 83.725 ;
        RECT 45.135 82.425 45.305 82.595 ;
        RECT 45.895 82.425 46.065 83.555 ;
        RECT 42.865 81.855 43.125 82.360 ;
        RECT 43.320 82.235 43.985 82.405 ;
        RECT 43.305 81.685 43.635 82.065 ;
        RECT 43.815 81.855 43.985 82.235 ;
        RECT 44.245 81.685 44.535 82.410 ;
        RECT 44.710 81.855 44.965 82.425 ;
        RECT 45.135 82.255 46.065 82.425 ;
        RECT 46.235 83.215 47.245 83.385 ;
        RECT 46.235 82.415 46.405 83.215 ;
        RECT 46.610 82.875 46.885 83.015 ;
        RECT 46.605 82.705 46.885 82.875 ;
        RECT 45.890 82.220 46.065 82.255 ;
        RECT 45.135 81.685 45.465 82.085 ;
        RECT 45.890 81.855 46.420 82.220 ;
        RECT 46.610 81.855 46.885 82.705 ;
        RECT 47.055 81.855 47.245 83.215 ;
        RECT 47.415 83.230 47.585 83.895 ;
        RECT 47.755 83.475 47.925 84.235 ;
        RECT 48.160 83.475 48.675 83.885 ;
        RECT 47.415 83.040 48.165 83.230 ;
        RECT 48.335 82.665 48.675 83.475 ;
        RECT 48.845 83.145 50.055 84.235 ;
        RECT 47.445 82.495 48.675 82.665 ;
        RECT 47.425 81.685 47.935 82.220 ;
        RECT 48.155 81.890 48.400 82.495 ;
        RECT 48.845 82.435 49.365 82.975 ;
        RECT 49.535 82.605 50.055 83.145 ;
        RECT 50.430 83.265 50.760 84.065 ;
        RECT 50.930 83.435 51.260 84.235 ;
        RECT 51.560 83.265 51.890 84.065 ;
        RECT 52.535 83.435 52.785 84.235 ;
        RECT 50.430 83.095 52.865 83.265 ;
        RECT 53.055 83.095 53.225 84.235 ;
        RECT 53.395 83.095 53.735 84.065 ;
        RECT 53.905 83.145 55.575 84.235 ;
        RECT 56.295 83.565 56.465 84.065 ;
        RECT 56.635 83.735 56.965 84.235 ;
        RECT 56.295 83.395 56.960 83.565 ;
        RECT 50.225 82.675 50.575 82.925 ;
        RECT 50.760 82.465 50.930 83.095 ;
        RECT 51.100 82.675 51.430 82.875 ;
        RECT 51.600 82.675 51.930 82.875 ;
        RECT 52.100 82.675 52.520 82.875 ;
        RECT 52.695 82.845 52.865 83.095 ;
        RECT 52.695 82.675 53.390 82.845 ;
        RECT 48.845 81.685 50.055 82.435 ;
        RECT 50.430 81.855 50.930 82.465 ;
        RECT 51.560 82.335 52.785 82.505 ;
        RECT 53.560 82.485 53.735 83.095 ;
        RECT 51.560 81.855 51.890 82.335 ;
        RECT 52.060 81.685 52.285 82.145 ;
        RECT 52.455 81.855 52.785 82.335 ;
        RECT 52.975 81.685 53.225 82.485 ;
        RECT 53.395 81.855 53.735 82.485 ;
        RECT 53.905 82.455 54.655 82.975 ;
        RECT 54.825 82.625 55.575 83.145 ;
        RECT 56.210 82.575 56.560 83.225 ;
        RECT 53.905 81.685 55.575 82.455 ;
        RECT 56.730 82.405 56.960 83.395 ;
        RECT 56.295 82.235 56.960 82.405 ;
        RECT 56.295 81.945 56.465 82.235 ;
        RECT 56.635 81.685 56.965 82.065 ;
        RECT 57.135 81.945 57.360 84.065 ;
        RECT 57.575 83.735 57.905 84.235 ;
        RECT 58.075 83.565 58.245 84.065 ;
        RECT 58.480 83.850 59.310 84.020 ;
        RECT 59.550 83.855 59.930 84.235 ;
        RECT 57.550 83.395 58.245 83.565 ;
        RECT 57.550 82.425 57.720 83.395 ;
        RECT 57.890 82.605 58.300 83.225 ;
        RECT 58.470 83.175 58.970 83.555 ;
        RECT 57.550 82.235 58.245 82.425 ;
        RECT 58.470 82.305 58.690 83.175 ;
        RECT 59.140 83.005 59.310 83.850 ;
        RECT 60.110 83.685 60.280 83.975 ;
        RECT 60.450 83.855 60.780 84.235 ;
        RECT 61.250 83.765 61.880 84.015 ;
        RECT 62.060 83.855 62.480 84.235 ;
        RECT 61.710 83.685 61.880 83.765 ;
        RECT 62.680 83.685 62.920 83.975 ;
        RECT 59.480 83.435 60.850 83.685 ;
        RECT 59.480 83.175 59.730 83.435 ;
        RECT 60.240 83.005 60.490 83.165 ;
        RECT 59.140 82.835 60.490 83.005 ;
        RECT 59.140 82.795 59.560 82.835 ;
        RECT 58.870 82.245 59.220 82.615 ;
        RECT 57.575 81.685 57.905 82.065 ;
        RECT 58.075 81.905 58.245 82.235 ;
        RECT 59.390 82.065 59.560 82.795 ;
        RECT 60.660 82.665 60.850 83.435 ;
        RECT 59.730 82.335 60.140 82.665 ;
        RECT 60.430 82.325 60.850 82.665 ;
        RECT 61.020 83.255 61.540 83.565 ;
        RECT 61.710 83.515 62.920 83.685 ;
        RECT 63.150 83.545 63.480 84.235 ;
        RECT 61.020 82.495 61.190 83.255 ;
        RECT 61.360 82.665 61.540 83.075 ;
        RECT 61.710 83.005 61.880 83.515 ;
        RECT 63.650 83.365 63.820 83.975 ;
        RECT 64.090 83.515 64.420 84.025 ;
        RECT 63.650 83.345 63.970 83.365 ;
        RECT 62.050 83.175 63.970 83.345 ;
        RECT 61.710 82.835 63.610 83.005 ;
        RECT 61.940 82.495 62.270 82.615 ;
        RECT 61.020 82.325 62.270 82.495 ;
        RECT 58.545 81.865 59.560 82.065 ;
        RECT 59.730 81.685 60.140 82.125 ;
        RECT 60.430 81.895 60.680 82.325 ;
        RECT 60.880 81.685 61.200 82.145 ;
        RECT 62.440 82.075 62.610 82.835 ;
        RECT 63.280 82.775 63.610 82.835 ;
        RECT 62.800 82.605 63.130 82.665 ;
        RECT 62.800 82.335 63.460 82.605 ;
        RECT 63.780 82.280 63.970 83.175 ;
        RECT 61.760 81.905 62.610 82.075 ;
        RECT 62.810 81.685 63.470 82.165 ;
        RECT 63.650 81.950 63.970 82.280 ;
        RECT 64.170 82.925 64.420 83.515 ;
        RECT 64.600 83.435 64.885 84.235 ;
        RECT 65.065 83.255 65.320 83.925 ;
        RECT 64.170 82.595 64.970 82.925 ;
        RECT 64.170 81.945 64.420 82.595 ;
        RECT 65.140 82.395 65.320 83.255 ;
        RECT 66.070 83.265 66.400 84.065 ;
        RECT 66.570 83.435 66.900 84.235 ;
        RECT 67.200 83.265 67.530 84.065 ;
        RECT 68.175 83.435 68.425 84.235 ;
        RECT 66.070 83.095 68.505 83.265 ;
        RECT 68.695 83.095 68.865 84.235 ;
        RECT 69.035 83.095 69.375 84.065 ;
        RECT 65.865 82.675 66.215 82.925 ;
        RECT 66.400 82.465 66.570 83.095 ;
        RECT 66.740 82.675 67.070 82.875 ;
        RECT 67.240 82.675 67.570 82.875 ;
        RECT 67.740 82.675 68.160 82.875 ;
        RECT 68.335 82.845 68.505 83.095 ;
        RECT 68.335 82.675 69.030 82.845 ;
        RECT 65.065 82.195 65.320 82.395 ;
        RECT 64.600 81.685 64.885 82.145 ;
        RECT 65.065 82.025 65.405 82.195 ;
        RECT 65.065 81.865 65.320 82.025 ;
        RECT 66.070 81.855 66.570 82.465 ;
        RECT 67.200 82.335 68.425 82.505 ;
        RECT 69.200 82.485 69.375 83.095 ;
        RECT 70.005 83.070 70.295 84.235 ;
        RECT 70.670 83.265 71.000 84.065 ;
        RECT 71.170 83.435 71.500 84.235 ;
        RECT 71.800 83.265 72.130 84.065 ;
        RECT 72.775 83.435 73.025 84.235 ;
        RECT 70.670 83.095 73.105 83.265 ;
        RECT 73.295 83.095 73.465 84.235 ;
        RECT 73.635 83.095 73.975 84.065 ;
        RECT 74.145 83.145 75.815 84.235 ;
        RECT 70.465 82.675 70.815 82.925 ;
        RECT 67.200 81.855 67.530 82.335 ;
        RECT 67.700 81.685 67.925 82.145 ;
        RECT 68.095 81.855 68.425 82.335 ;
        RECT 68.615 81.685 68.865 82.485 ;
        RECT 69.035 81.855 69.375 82.485 ;
        RECT 71.000 82.465 71.170 83.095 ;
        RECT 71.340 82.675 71.670 82.875 ;
        RECT 71.840 82.675 72.170 82.875 ;
        RECT 72.340 82.675 72.760 82.875 ;
        RECT 72.935 82.845 73.105 83.095 ;
        RECT 72.935 82.675 73.630 82.845 ;
        RECT 70.005 81.685 70.295 82.410 ;
        RECT 70.670 81.855 71.170 82.465 ;
        RECT 71.800 82.335 73.025 82.505 ;
        RECT 73.800 82.485 73.975 83.095 ;
        RECT 71.800 81.855 72.130 82.335 ;
        RECT 72.300 81.685 72.525 82.145 ;
        RECT 72.695 81.855 73.025 82.335 ;
        RECT 73.215 81.685 73.465 82.485 ;
        RECT 73.635 81.855 73.975 82.485 ;
        RECT 74.145 82.455 74.895 82.975 ;
        RECT 75.065 82.625 75.815 83.145 ;
        RECT 76.505 83.095 76.715 84.235 ;
        RECT 76.885 83.085 77.215 84.065 ;
        RECT 77.385 83.095 77.615 84.235 ;
        RECT 77.825 83.800 83.170 84.235 ;
        RECT 83.345 83.800 88.690 84.235 ;
        RECT 74.145 81.685 75.815 82.455 ;
        RECT 76.505 81.685 76.715 82.505 ;
        RECT 76.885 82.485 77.135 83.085 ;
        RECT 77.305 82.675 77.635 82.925 ;
        RECT 76.885 81.855 77.215 82.485 ;
        RECT 77.385 81.685 77.615 82.505 ;
        RECT 79.410 82.230 79.750 83.060 ;
        RECT 81.230 82.550 81.580 83.800 ;
        RECT 84.930 82.230 85.270 83.060 ;
        RECT 86.750 82.550 87.100 83.800 ;
        RECT 88.865 83.145 91.455 84.235 ;
        RECT 92.090 83.725 93.745 84.015 ;
        RECT 88.865 82.455 90.075 82.975 ;
        RECT 90.245 82.625 91.455 83.145 ;
        RECT 92.090 83.385 93.680 83.555 ;
        RECT 93.915 83.435 94.195 84.235 ;
        RECT 92.090 83.095 92.410 83.385 ;
        RECT 93.510 83.265 93.680 83.385 ;
        RECT 77.825 81.685 83.170 82.230 ;
        RECT 83.345 81.685 88.690 82.230 ;
        RECT 88.865 81.685 91.455 82.455 ;
        RECT 92.090 82.355 92.440 82.925 ;
        RECT 92.610 82.595 93.320 83.215 ;
        RECT 93.510 83.095 94.235 83.265 ;
        RECT 94.405 83.095 94.675 84.065 ;
        RECT 94.065 82.925 94.235 83.095 ;
        RECT 93.490 82.595 93.895 82.925 ;
        RECT 94.065 82.595 94.335 82.925 ;
        RECT 94.065 82.425 94.235 82.595 ;
        RECT 92.625 82.255 94.235 82.425 ;
        RECT 94.505 82.360 94.675 83.095 ;
        RECT 95.765 83.070 96.055 84.235 ;
        RECT 97.145 83.515 97.605 84.065 ;
        RECT 97.795 83.515 98.125 84.235 ;
        RECT 92.095 81.685 92.425 82.185 ;
        RECT 92.625 81.905 92.795 82.255 ;
        RECT 92.995 81.685 93.325 82.085 ;
        RECT 93.495 81.905 93.665 82.255 ;
        RECT 93.835 81.685 94.215 82.085 ;
        RECT 94.405 82.015 94.675 82.360 ;
        RECT 95.765 81.685 96.055 82.410 ;
        RECT 97.145 82.145 97.395 83.515 ;
        RECT 98.325 83.345 98.625 83.895 ;
        RECT 98.795 83.565 99.075 84.235 ;
        RECT 99.445 83.800 104.790 84.235 ;
        RECT 97.685 83.175 98.625 83.345 ;
        RECT 97.685 82.925 97.855 83.175 ;
        RECT 98.995 82.925 99.260 83.285 ;
        RECT 97.565 82.595 97.855 82.925 ;
        RECT 98.025 82.675 98.365 82.925 ;
        RECT 98.585 82.675 99.260 82.925 ;
        RECT 97.685 82.505 97.855 82.595 ;
        RECT 97.685 82.315 99.075 82.505 ;
        RECT 97.145 81.855 97.705 82.145 ;
        RECT 97.875 81.685 98.125 82.145 ;
        RECT 98.745 81.955 99.075 82.315 ;
        RECT 101.030 82.230 101.370 83.060 ;
        RECT 102.850 82.550 103.200 83.800 ;
        RECT 104.965 83.145 107.555 84.235 ;
        RECT 107.815 83.565 107.985 84.065 ;
        RECT 108.155 83.735 108.485 84.235 ;
        RECT 107.815 83.395 108.480 83.565 ;
        RECT 104.965 82.455 106.175 82.975 ;
        RECT 106.345 82.625 107.555 83.145 ;
        RECT 107.730 82.575 108.080 83.225 ;
        RECT 99.445 81.685 104.790 82.230 ;
        RECT 104.965 81.685 107.555 82.455 ;
        RECT 108.250 82.405 108.480 83.395 ;
        RECT 107.815 82.235 108.480 82.405 ;
        RECT 107.815 81.945 107.985 82.235 ;
        RECT 108.155 81.685 108.485 82.065 ;
        RECT 108.655 81.945 108.880 84.065 ;
        RECT 109.095 83.735 109.425 84.235 ;
        RECT 109.595 83.565 109.765 84.065 ;
        RECT 110.000 83.850 110.830 84.020 ;
        RECT 111.070 83.855 111.450 84.235 ;
        RECT 109.070 83.395 109.765 83.565 ;
        RECT 109.070 82.425 109.240 83.395 ;
        RECT 109.410 82.605 109.820 83.225 ;
        RECT 109.990 83.175 110.490 83.555 ;
        RECT 109.070 82.235 109.765 82.425 ;
        RECT 109.990 82.305 110.210 83.175 ;
        RECT 110.660 83.005 110.830 83.850 ;
        RECT 111.630 83.685 111.800 83.975 ;
        RECT 111.970 83.855 112.300 84.235 ;
        RECT 112.770 83.765 113.400 84.015 ;
        RECT 113.580 83.855 114.000 84.235 ;
        RECT 113.230 83.685 113.400 83.765 ;
        RECT 114.200 83.685 114.440 83.975 ;
        RECT 111.000 83.435 112.370 83.685 ;
        RECT 111.000 83.175 111.250 83.435 ;
        RECT 111.760 83.005 112.010 83.165 ;
        RECT 110.660 82.835 112.010 83.005 ;
        RECT 110.660 82.795 111.080 82.835 ;
        RECT 110.390 82.245 110.740 82.615 ;
        RECT 109.095 81.685 109.425 82.065 ;
        RECT 109.595 81.905 109.765 82.235 ;
        RECT 110.910 82.065 111.080 82.795 ;
        RECT 112.180 82.665 112.370 83.435 ;
        RECT 111.250 82.335 111.660 82.665 ;
        RECT 111.950 82.325 112.370 82.665 ;
        RECT 112.540 83.255 113.060 83.565 ;
        RECT 113.230 83.515 114.440 83.685 ;
        RECT 114.670 83.545 115.000 84.235 ;
        RECT 112.540 82.495 112.710 83.255 ;
        RECT 112.880 82.665 113.060 83.075 ;
        RECT 113.230 83.005 113.400 83.515 ;
        RECT 115.170 83.365 115.340 83.975 ;
        RECT 115.610 83.515 115.940 84.025 ;
        RECT 115.170 83.345 115.490 83.365 ;
        RECT 113.570 83.175 115.490 83.345 ;
        RECT 113.230 82.835 115.130 83.005 ;
        RECT 113.460 82.495 113.790 82.615 ;
        RECT 112.540 82.325 113.790 82.495 ;
        RECT 110.065 81.865 111.080 82.065 ;
        RECT 111.250 81.685 111.660 82.125 ;
        RECT 111.950 81.895 112.200 82.325 ;
        RECT 112.400 81.685 112.720 82.145 ;
        RECT 113.960 82.075 114.130 82.835 ;
        RECT 114.800 82.775 115.130 82.835 ;
        RECT 114.320 82.605 114.650 82.665 ;
        RECT 114.320 82.335 114.980 82.605 ;
        RECT 115.300 82.280 115.490 83.175 ;
        RECT 113.280 81.905 114.130 82.075 ;
        RECT 114.330 81.685 114.990 82.165 ;
        RECT 115.170 81.950 115.490 82.280 ;
        RECT 115.690 82.925 115.940 83.515 ;
        RECT 116.120 83.435 116.405 84.235 ;
        RECT 116.585 83.895 116.840 83.925 ;
        RECT 116.585 83.725 116.925 83.895 ;
        RECT 116.585 83.255 116.840 83.725 ;
        RECT 115.690 82.595 116.490 82.925 ;
        RECT 115.690 81.945 115.940 82.595 ;
        RECT 116.660 82.395 116.840 83.255 ;
        RECT 117.385 83.145 118.595 84.235 ;
        RECT 117.385 82.605 117.905 83.145 ;
        RECT 118.075 82.435 118.595 82.975 ;
        RECT 116.120 81.685 116.405 82.145 ;
        RECT 116.585 81.865 116.840 82.395 ;
        RECT 117.385 81.685 118.595 82.435 ;
        RECT 5.520 81.515 118.680 81.685 ;
        RECT 5.605 80.765 6.815 81.515 ;
        RECT 5.605 80.225 6.125 80.765 ;
        RECT 6.985 80.745 10.495 81.515 ;
        RECT 10.665 80.765 11.875 81.515 ;
        RECT 6.295 80.055 6.815 80.595 ;
        RECT 6.985 80.225 8.635 80.745 ;
        RECT 8.805 80.055 10.495 80.575 ;
        RECT 10.665 80.225 11.185 80.765 ;
        RECT 12.105 80.695 12.315 81.515 ;
        RECT 12.485 80.715 12.815 81.345 ;
        RECT 11.355 80.055 11.875 80.595 ;
        RECT 12.485 80.115 12.735 80.715 ;
        RECT 12.985 80.695 13.215 81.515 ;
        RECT 13.430 80.775 13.685 81.345 ;
        RECT 13.855 81.115 14.185 81.515 ;
        RECT 14.610 80.980 15.140 81.345 ;
        RECT 14.610 80.945 14.785 80.980 ;
        RECT 13.855 80.775 14.785 80.945 ;
        RECT 12.905 80.275 13.235 80.525 ;
        RECT 5.605 78.965 6.815 80.055 ;
        RECT 6.985 78.965 10.495 80.055 ;
        RECT 10.665 78.965 11.875 80.055 ;
        RECT 12.105 78.965 12.315 80.105 ;
        RECT 12.485 79.135 12.815 80.115 ;
        RECT 13.430 80.105 13.600 80.775 ;
        RECT 13.855 80.605 14.025 80.775 ;
        RECT 13.770 80.275 14.025 80.605 ;
        RECT 14.250 80.275 14.445 80.605 ;
        RECT 12.985 78.965 13.215 80.105 ;
        RECT 13.430 79.135 13.765 80.105 ;
        RECT 13.935 78.965 14.105 80.105 ;
        RECT 14.275 79.305 14.445 80.275 ;
        RECT 14.615 79.645 14.785 80.775 ;
        RECT 14.955 79.985 15.125 80.785 ;
        RECT 15.330 80.495 15.605 81.345 ;
        RECT 15.325 80.325 15.605 80.495 ;
        RECT 15.330 80.185 15.605 80.325 ;
        RECT 15.775 79.985 15.965 81.345 ;
        RECT 16.145 80.980 16.655 81.515 ;
        RECT 16.875 80.705 17.120 81.310 ;
        RECT 17.565 80.970 22.910 81.515 ;
        RECT 23.085 80.970 28.430 81.515 ;
        RECT 16.165 80.535 17.395 80.705 ;
        RECT 14.955 79.815 15.965 79.985 ;
        RECT 16.135 79.970 16.885 80.160 ;
        RECT 14.615 79.475 15.740 79.645 ;
        RECT 16.135 79.305 16.305 79.970 ;
        RECT 17.055 79.725 17.395 80.535 ;
        RECT 19.150 80.140 19.490 80.970 ;
        RECT 14.275 79.135 16.305 79.305 ;
        RECT 16.475 78.965 16.645 79.725 ;
        RECT 16.880 79.315 17.395 79.725 ;
        RECT 20.970 79.400 21.320 80.650 ;
        RECT 24.670 80.140 25.010 80.970 ;
        RECT 28.605 80.745 31.195 81.515 ;
        RECT 31.365 80.790 31.655 81.515 ;
        RECT 31.825 80.970 37.170 81.515 ;
        RECT 37.345 80.970 42.690 81.515 ;
        RECT 42.865 80.970 48.210 81.515 ;
        RECT 48.385 80.970 53.730 81.515 ;
        RECT 26.490 79.400 26.840 80.650 ;
        RECT 28.605 80.225 29.815 80.745 ;
        RECT 29.985 80.055 31.195 80.575 ;
        RECT 33.410 80.140 33.750 80.970 ;
        RECT 17.565 78.965 22.910 79.400 ;
        RECT 23.085 78.965 28.430 79.400 ;
        RECT 28.605 78.965 31.195 80.055 ;
        RECT 31.365 78.965 31.655 80.130 ;
        RECT 35.230 79.400 35.580 80.650 ;
        RECT 38.930 80.140 39.270 80.970 ;
        RECT 40.750 79.400 41.100 80.650 ;
        RECT 44.450 80.140 44.790 80.970 ;
        RECT 46.270 79.400 46.620 80.650 ;
        RECT 49.970 80.140 50.310 80.970 ;
        RECT 53.905 80.745 56.495 81.515 ;
        RECT 57.125 80.790 57.415 81.515 ;
        RECT 57.585 80.745 60.175 81.515 ;
        RECT 51.790 79.400 52.140 80.650 ;
        RECT 53.905 80.225 55.115 80.745 ;
        RECT 55.285 80.055 56.495 80.575 ;
        RECT 57.585 80.225 58.795 80.745 ;
        RECT 60.385 80.695 60.615 81.515 ;
        RECT 60.785 80.715 61.115 81.345 ;
        RECT 31.825 78.965 37.170 79.400 ;
        RECT 37.345 78.965 42.690 79.400 ;
        RECT 42.865 78.965 48.210 79.400 ;
        RECT 48.385 78.965 53.730 79.400 ;
        RECT 53.905 78.965 56.495 80.055 ;
        RECT 57.125 78.965 57.415 80.130 ;
        RECT 58.965 80.055 60.175 80.575 ;
        RECT 60.365 80.275 60.695 80.525 ;
        RECT 60.865 80.115 61.115 80.715 ;
        RECT 61.285 80.695 61.495 81.515 ;
        RECT 61.725 80.765 62.935 81.515 ;
        RECT 63.195 80.965 63.365 81.345 ;
        RECT 63.545 81.135 63.875 81.515 ;
        RECT 63.195 80.795 63.860 80.965 ;
        RECT 64.055 80.840 64.315 81.345 ;
        RECT 61.725 80.225 62.245 80.765 ;
        RECT 57.585 78.965 60.175 80.055 ;
        RECT 60.385 78.965 60.615 80.105 ;
        RECT 60.785 79.135 61.115 80.115 ;
        RECT 61.285 78.965 61.495 80.105 ;
        RECT 62.415 80.055 62.935 80.595 ;
        RECT 63.125 80.245 63.455 80.615 ;
        RECT 63.690 80.540 63.860 80.795 ;
        RECT 63.690 80.210 63.975 80.540 ;
        RECT 63.690 80.065 63.860 80.210 ;
        RECT 61.725 78.965 62.935 80.055 ;
        RECT 63.195 79.895 63.860 80.065 ;
        RECT 64.145 80.040 64.315 80.840 ;
        RECT 64.490 80.965 64.745 81.255 ;
        RECT 64.915 81.135 65.245 81.515 ;
        RECT 64.490 80.795 65.240 80.965 ;
        RECT 63.195 79.135 63.365 79.895 ;
        RECT 63.545 78.965 63.875 79.725 ;
        RECT 64.045 79.135 64.315 80.040 ;
        RECT 64.490 79.975 64.840 80.625 ;
        RECT 65.010 79.805 65.240 80.795 ;
        RECT 64.490 79.635 65.240 79.805 ;
        RECT 64.490 79.135 64.745 79.635 ;
        RECT 64.915 78.965 65.245 79.465 ;
        RECT 65.415 79.135 65.585 81.255 ;
        RECT 65.945 81.155 66.275 81.515 ;
        RECT 66.445 81.125 66.940 81.295 ;
        RECT 67.145 81.125 68.000 81.295 ;
        RECT 65.815 79.935 66.275 80.985 ;
        RECT 65.755 79.150 66.080 79.935 ;
        RECT 66.445 79.765 66.615 81.125 ;
        RECT 66.785 80.215 67.135 80.835 ;
        RECT 67.305 80.615 67.660 80.835 ;
        RECT 67.305 80.025 67.475 80.615 ;
        RECT 67.830 80.415 68.000 81.125 ;
        RECT 68.875 81.055 69.205 81.515 ;
        RECT 69.415 81.155 69.765 81.325 ;
        RECT 68.205 80.585 68.995 80.835 ;
        RECT 69.415 80.765 69.675 81.155 ;
        RECT 69.985 81.065 70.935 81.345 ;
        RECT 71.105 81.075 71.295 81.515 ;
        RECT 71.465 81.135 72.535 81.305 ;
        RECT 69.165 80.415 69.335 80.595 ;
        RECT 66.445 79.595 66.840 79.765 ;
        RECT 67.010 79.635 67.475 80.025 ;
        RECT 67.645 80.245 69.335 80.415 ;
        RECT 66.670 79.465 66.840 79.595 ;
        RECT 67.645 79.465 67.815 80.245 ;
        RECT 69.505 80.075 69.675 80.765 ;
        RECT 68.175 79.905 69.675 80.075 ;
        RECT 69.865 80.105 70.075 80.895 ;
        RECT 70.245 80.275 70.595 80.895 ;
        RECT 70.765 80.285 70.935 81.065 ;
        RECT 71.465 80.905 71.635 81.135 ;
        RECT 71.105 80.735 71.635 80.905 ;
        RECT 71.105 80.455 71.325 80.735 ;
        RECT 71.805 80.565 72.045 80.965 ;
        RECT 70.765 80.115 71.170 80.285 ;
        RECT 71.505 80.195 72.045 80.565 ;
        RECT 72.215 80.780 72.535 81.135 ;
        RECT 72.780 81.055 73.085 81.515 ;
        RECT 73.255 80.805 73.510 81.335 ;
        RECT 72.215 80.605 72.540 80.780 ;
        RECT 72.215 80.305 73.130 80.605 ;
        RECT 72.390 80.275 73.130 80.305 ;
        RECT 69.865 79.945 70.540 80.105 ;
        RECT 71.000 80.025 71.170 80.115 ;
        RECT 69.865 79.935 70.830 79.945 ;
        RECT 69.505 79.765 69.675 79.905 ;
        RECT 66.250 78.965 66.500 79.425 ;
        RECT 66.670 79.135 66.920 79.465 ;
        RECT 67.135 79.135 67.815 79.465 ;
        RECT 67.985 79.565 69.060 79.735 ;
        RECT 69.505 79.595 70.065 79.765 ;
        RECT 70.370 79.645 70.830 79.935 ;
        RECT 71.000 79.855 72.220 80.025 ;
        RECT 67.985 79.225 68.155 79.565 ;
        RECT 68.390 78.965 68.720 79.395 ;
        RECT 68.890 79.225 69.060 79.565 ;
        RECT 69.355 78.965 69.725 79.425 ;
        RECT 69.895 79.135 70.065 79.595 ;
        RECT 71.000 79.475 71.170 79.855 ;
        RECT 72.390 79.685 72.560 80.275 ;
        RECT 73.300 80.155 73.510 80.805 ;
        RECT 70.300 79.135 71.170 79.475 ;
        RECT 71.760 79.515 72.560 79.685 ;
        RECT 71.340 78.965 71.590 79.425 ;
        RECT 71.760 79.225 71.930 79.515 ;
        RECT 72.110 78.965 72.440 79.345 ;
        RECT 72.780 78.965 73.085 80.105 ;
        RECT 73.255 79.275 73.510 80.155 ;
        RECT 73.685 80.775 74.070 81.345 ;
        RECT 74.240 81.055 74.565 81.515 ;
        RECT 75.085 80.885 75.365 81.345 ;
        RECT 73.685 80.105 73.965 80.775 ;
        RECT 74.240 80.715 75.365 80.885 ;
        RECT 74.240 80.605 74.690 80.715 ;
        RECT 74.135 80.275 74.690 80.605 ;
        RECT 75.555 80.545 75.955 81.345 ;
        RECT 76.355 81.055 76.625 81.515 ;
        RECT 76.795 80.885 77.080 81.345 ;
        RECT 73.685 79.135 74.070 80.105 ;
        RECT 74.240 79.815 74.690 80.275 ;
        RECT 74.860 79.985 75.955 80.545 ;
        RECT 74.240 79.595 75.365 79.815 ;
        RECT 74.240 78.965 74.565 79.425 ;
        RECT 75.085 79.135 75.365 79.595 ;
        RECT 75.555 79.135 75.955 79.985 ;
        RECT 76.125 80.715 77.080 80.885 ;
        RECT 77.570 80.735 78.070 81.345 ;
        RECT 76.125 79.815 76.335 80.715 ;
        RECT 76.505 79.985 77.195 80.545 ;
        RECT 77.365 80.275 77.715 80.525 ;
        RECT 77.900 80.105 78.070 80.735 ;
        RECT 78.700 80.865 79.030 81.345 ;
        RECT 79.200 81.055 79.425 81.515 ;
        RECT 79.595 80.865 79.925 81.345 ;
        RECT 78.700 80.695 79.925 80.865 ;
        RECT 80.115 80.715 80.365 81.515 ;
        RECT 80.535 80.715 80.875 81.345 ;
        RECT 80.645 80.665 80.875 80.715 ;
        RECT 78.240 80.325 78.570 80.525 ;
        RECT 78.740 80.325 79.070 80.525 ;
        RECT 79.240 80.325 79.660 80.525 ;
        RECT 79.835 80.355 80.530 80.525 ;
        RECT 79.835 80.105 80.005 80.355 ;
        RECT 80.700 80.105 80.875 80.665 ;
        RECT 81.045 80.745 82.715 81.515 ;
        RECT 82.885 80.790 83.175 81.515 ;
        RECT 83.355 81.015 83.685 81.515 ;
        RECT 83.885 80.945 84.055 81.295 ;
        RECT 84.255 81.115 84.585 81.515 ;
        RECT 84.755 80.945 84.925 81.295 ;
        RECT 85.095 81.115 85.475 81.515 ;
        RECT 81.045 80.225 81.795 80.745 ;
        RECT 77.570 79.935 80.005 80.105 ;
        RECT 76.125 79.595 77.080 79.815 ;
        RECT 76.355 78.965 76.625 79.425 ;
        RECT 76.795 79.135 77.080 79.595 ;
        RECT 77.570 79.135 77.900 79.935 ;
        RECT 78.070 78.965 78.400 79.765 ;
        RECT 78.700 79.135 79.030 79.935 ;
        RECT 79.675 78.965 79.925 79.765 ;
        RECT 80.195 78.965 80.365 80.105 ;
        RECT 80.535 79.135 80.875 80.105 ;
        RECT 81.965 80.055 82.715 80.575 ;
        RECT 83.350 80.275 83.700 80.845 ;
        RECT 83.885 80.775 85.495 80.945 ;
        RECT 85.665 80.840 85.935 81.185 ;
        RECT 86.105 80.970 91.450 81.515 ;
        RECT 85.325 80.605 85.495 80.775 ;
        RECT 81.045 78.965 82.715 80.055 ;
        RECT 82.885 78.965 83.175 80.130 ;
        RECT 83.350 79.815 83.670 80.105 ;
        RECT 83.870 79.985 84.580 80.605 ;
        RECT 84.750 80.275 85.155 80.605 ;
        RECT 85.325 80.275 85.595 80.605 ;
        RECT 85.325 80.105 85.495 80.275 ;
        RECT 85.765 80.105 85.935 80.840 ;
        RECT 87.690 80.140 88.030 80.970 ;
        RECT 91.625 80.745 95.135 81.515 ;
        RECT 96.235 81.015 96.565 81.515 ;
        RECT 96.765 80.945 96.935 81.295 ;
        RECT 97.135 81.115 97.465 81.515 ;
        RECT 97.635 80.945 97.805 81.295 ;
        RECT 97.975 81.115 98.355 81.515 ;
        RECT 84.770 79.935 85.495 80.105 ;
        RECT 84.770 79.815 84.940 79.935 ;
        RECT 83.350 79.645 84.940 79.815 ;
        RECT 83.350 79.185 85.005 79.475 ;
        RECT 85.175 78.965 85.455 79.765 ;
        RECT 85.665 79.135 85.935 80.105 ;
        RECT 89.510 79.400 89.860 80.650 ;
        RECT 91.625 80.225 93.275 80.745 ;
        RECT 93.445 80.055 95.135 80.575 ;
        RECT 96.230 80.275 96.580 80.845 ;
        RECT 96.765 80.775 98.375 80.945 ;
        RECT 98.545 80.840 98.815 81.185 ;
        RECT 98.985 80.970 104.330 81.515 ;
        RECT 98.205 80.605 98.375 80.775 ;
        RECT 86.105 78.965 91.450 79.400 ;
        RECT 91.625 78.965 95.135 80.055 ;
        RECT 96.230 79.815 96.550 80.105 ;
        RECT 96.750 79.985 97.460 80.605 ;
        RECT 97.630 80.275 98.035 80.605 ;
        RECT 98.205 80.275 98.475 80.605 ;
        RECT 98.205 80.105 98.375 80.275 ;
        RECT 98.645 80.105 98.815 80.840 ;
        RECT 100.570 80.140 100.910 80.970 ;
        RECT 104.505 80.745 108.015 81.515 ;
        RECT 108.645 80.790 108.935 81.515 ;
        RECT 109.105 80.970 114.450 81.515 ;
        RECT 97.650 79.935 98.375 80.105 ;
        RECT 97.650 79.815 97.820 79.935 ;
        RECT 96.230 79.645 97.820 79.815 ;
        RECT 96.230 79.185 97.885 79.475 ;
        RECT 98.055 78.965 98.335 79.765 ;
        RECT 98.545 79.135 98.815 80.105 ;
        RECT 102.390 79.400 102.740 80.650 ;
        RECT 104.505 80.225 106.155 80.745 ;
        RECT 106.325 80.055 108.015 80.575 ;
        RECT 110.690 80.140 111.030 80.970 ;
        RECT 114.625 80.745 117.215 81.515 ;
        RECT 117.385 80.765 118.595 81.515 ;
        RECT 98.985 78.965 104.330 79.400 ;
        RECT 104.505 78.965 108.015 80.055 ;
        RECT 108.645 78.965 108.935 80.130 ;
        RECT 112.510 79.400 112.860 80.650 ;
        RECT 114.625 80.225 115.835 80.745 ;
        RECT 116.005 80.055 117.215 80.575 ;
        RECT 109.105 78.965 114.450 79.400 ;
        RECT 114.625 78.965 117.215 80.055 ;
        RECT 117.385 80.055 117.905 80.595 ;
        RECT 118.075 80.225 118.595 80.765 ;
        RECT 117.385 78.965 118.595 80.055 ;
        RECT 5.520 78.795 118.680 78.965 ;
        RECT 5.605 77.705 6.815 78.795 ;
        RECT 6.985 77.705 10.495 78.795 ;
        RECT 5.605 76.995 6.125 77.535 ;
        RECT 6.295 77.165 6.815 77.705 ;
        RECT 6.985 77.015 8.635 77.535 ;
        RECT 8.805 77.185 10.495 77.705 ;
        RECT 10.665 77.720 10.935 78.625 ;
        RECT 11.105 78.035 11.435 78.795 ;
        RECT 11.615 77.865 11.785 78.625 ;
        RECT 5.605 76.245 6.815 76.995 ;
        RECT 6.985 76.245 10.495 77.015 ;
        RECT 10.665 76.920 10.835 77.720 ;
        RECT 11.120 77.695 11.785 77.865 ;
        RECT 11.120 77.550 11.290 77.695 ;
        RECT 12.565 77.655 12.775 78.795 ;
        RECT 11.005 77.220 11.290 77.550 ;
        RECT 12.945 77.645 13.275 78.625 ;
        RECT 13.445 77.655 13.675 78.795 ;
        RECT 13.890 77.655 14.225 78.625 ;
        RECT 14.395 77.655 14.565 78.795 ;
        RECT 14.735 78.455 16.765 78.625 ;
        RECT 11.120 76.965 11.290 77.220 ;
        RECT 11.525 77.145 11.855 77.515 ;
        RECT 10.665 76.415 10.925 76.920 ;
        RECT 11.120 76.795 11.785 76.965 ;
        RECT 11.105 76.245 11.435 76.625 ;
        RECT 11.615 76.415 11.785 76.795 ;
        RECT 12.565 76.245 12.775 77.065 ;
        RECT 12.945 77.045 13.195 77.645 ;
        RECT 13.365 77.235 13.695 77.485 ;
        RECT 12.945 76.415 13.275 77.045 ;
        RECT 13.445 76.245 13.675 77.065 ;
        RECT 13.890 76.985 14.060 77.655 ;
        RECT 14.735 77.485 14.905 78.455 ;
        RECT 14.230 77.155 14.485 77.485 ;
        RECT 14.710 77.155 14.905 77.485 ;
        RECT 15.075 78.115 16.200 78.285 ;
        RECT 14.315 76.985 14.485 77.155 ;
        RECT 15.075 76.985 15.245 78.115 ;
        RECT 13.890 76.415 14.145 76.985 ;
        RECT 14.315 76.815 15.245 76.985 ;
        RECT 15.415 77.775 16.425 77.945 ;
        RECT 15.415 76.975 15.585 77.775 ;
        RECT 15.070 76.780 15.245 76.815 ;
        RECT 14.315 76.245 14.645 76.645 ;
        RECT 15.070 76.415 15.600 76.780 ;
        RECT 15.790 76.755 16.065 77.575 ;
        RECT 15.785 76.585 16.065 76.755 ;
        RECT 15.790 76.415 16.065 76.585 ;
        RECT 16.235 76.415 16.425 77.775 ;
        RECT 16.595 77.790 16.765 78.455 ;
        RECT 16.935 78.035 17.105 78.795 ;
        RECT 17.340 78.035 17.855 78.445 ;
        RECT 16.595 77.600 17.345 77.790 ;
        RECT 17.515 77.225 17.855 78.035 ;
        RECT 18.485 77.630 18.775 78.795 ;
        RECT 20.070 77.825 20.400 78.625 ;
        RECT 20.570 77.995 20.900 78.795 ;
        RECT 21.200 77.825 21.530 78.625 ;
        RECT 22.175 77.995 22.425 78.795 ;
        RECT 20.070 77.655 22.505 77.825 ;
        RECT 22.695 77.655 22.865 78.795 ;
        RECT 23.035 77.655 23.375 78.625 ;
        RECT 19.865 77.235 20.215 77.485 ;
        RECT 16.625 77.055 17.855 77.225 ;
        RECT 16.605 76.245 17.115 76.780 ;
        RECT 17.335 76.450 17.580 77.055 ;
        RECT 20.400 77.025 20.570 77.655 ;
        RECT 20.740 77.235 21.070 77.435 ;
        RECT 21.240 77.235 21.570 77.435 ;
        RECT 21.740 77.235 22.160 77.435 ;
        RECT 22.335 77.405 22.505 77.655 ;
        RECT 22.335 77.235 23.030 77.405 ;
        RECT 23.200 77.095 23.375 77.655 ;
        RECT 18.485 76.245 18.775 76.970 ;
        RECT 20.070 76.415 20.570 77.025 ;
        RECT 21.200 76.895 22.425 77.065 ;
        RECT 23.145 77.045 23.375 77.095 ;
        RECT 21.200 76.415 21.530 76.895 ;
        RECT 21.700 76.245 21.925 76.705 ;
        RECT 22.095 76.415 22.425 76.895 ;
        RECT 22.615 76.245 22.865 77.045 ;
        RECT 23.035 76.415 23.375 77.045 ;
        RECT 23.545 77.655 23.815 78.625 ;
        RECT 24.025 77.995 24.305 78.795 ;
        RECT 24.475 78.285 26.130 78.575 ;
        RECT 26.305 78.360 31.650 78.795 ;
        RECT 24.540 77.945 26.130 78.115 ;
        RECT 24.540 77.825 24.710 77.945 ;
        RECT 23.985 77.655 24.710 77.825 ;
        RECT 23.545 76.920 23.715 77.655 ;
        RECT 23.985 77.485 24.155 77.655 ;
        RECT 23.885 77.155 24.155 77.485 ;
        RECT 24.325 77.155 24.730 77.485 ;
        RECT 24.900 77.155 25.610 77.775 ;
        RECT 25.810 77.655 26.130 77.945 ;
        RECT 23.985 76.985 24.155 77.155 ;
        RECT 23.545 76.575 23.815 76.920 ;
        RECT 23.985 76.815 25.595 76.985 ;
        RECT 25.780 76.915 26.130 77.485 ;
        RECT 24.005 76.245 24.385 76.645 ;
        RECT 24.555 76.465 24.725 76.815 ;
        RECT 24.895 76.245 25.225 76.645 ;
        RECT 25.425 76.465 25.595 76.815 ;
        RECT 27.890 76.790 28.230 77.620 ;
        RECT 29.710 77.110 30.060 78.360 ;
        RECT 31.825 77.705 35.335 78.795 ;
        RECT 31.825 77.015 33.475 77.535 ;
        RECT 33.645 77.185 35.335 77.705 ;
        RECT 35.965 77.655 36.350 78.625 ;
        RECT 36.520 78.335 36.845 78.795 ;
        RECT 37.365 78.165 37.645 78.625 ;
        RECT 36.520 77.945 37.645 78.165 ;
        RECT 25.795 76.245 26.125 76.745 ;
        RECT 26.305 76.245 31.650 76.790 ;
        RECT 31.825 76.245 35.335 77.015 ;
        RECT 35.965 76.985 36.245 77.655 ;
        RECT 36.520 77.485 36.970 77.945 ;
        RECT 37.835 77.775 38.235 78.625 ;
        RECT 38.635 78.335 38.905 78.795 ;
        RECT 39.075 78.165 39.360 78.625 ;
        RECT 36.415 77.155 36.970 77.485 ;
        RECT 37.140 77.215 38.235 77.775 ;
        RECT 36.520 77.045 36.970 77.155 ;
        RECT 35.965 76.415 36.350 76.985 ;
        RECT 36.520 76.875 37.645 77.045 ;
        RECT 36.520 76.245 36.845 76.705 ;
        RECT 37.365 76.415 37.645 76.875 ;
        RECT 37.835 76.415 38.235 77.215 ;
        RECT 38.405 77.945 39.360 78.165 ;
        RECT 38.405 77.045 38.615 77.945 ;
        RECT 38.785 77.215 39.475 77.775 ;
        RECT 39.645 77.705 41.315 78.795 ;
        RECT 38.405 76.875 39.360 77.045 ;
        RECT 38.635 76.245 38.905 76.705 ;
        RECT 39.075 76.415 39.360 76.875 ;
        RECT 39.645 77.015 40.395 77.535 ;
        RECT 40.565 77.185 41.315 77.705 ;
        RECT 41.945 77.720 42.215 78.625 ;
        RECT 42.385 78.035 42.715 78.795 ;
        RECT 42.895 77.865 43.065 78.625 ;
        RECT 39.645 76.245 41.315 77.015 ;
        RECT 41.945 76.920 42.115 77.720 ;
        RECT 42.400 77.695 43.065 77.865 ;
        RECT 42.400 77.550 42.570 77.695 ;
        RECT 44.245 77.630 44.535 78.795 ;
        RECT 44.710 77.655 45.045 78.625 ;
        RECT 45.215 77.655 45.385 78.795 ;
        RECT 45.555 78.455 47.585 78.625 ;
        RECT 42.285 77.220 42.570 77.550 ;
        RECT 42.400 76.965 42.570 77.220 ;
        RECT 42.805 77.145 43.135 77.515 ;
        RECT 44.710 76.985 44.880 77.655 ;
        RECT 45.555 77.485 45.725 78.455 ;
        RECT 45.050 77.155 45.305 77.485 ;
        RECT 45.530 77.155 45.725 77.485 ;
        RECT 45.895 78.115 47.020 78.285 ;
        RECT 45.135 76.985 45.305 77.155 ;
        RECT 45.895 76.985 46.065 78.115 ;
        RECT 41.945 76.415 42.205 76.920 ;
        RECT 42.400 76.795 43.065 76.965 ;
        RECT 42.385 76.245 42.715 76.625 ;
        RECT 42.895 76.415 43.065 76.795 ;
        RECT 44.245 76.245 44.535 76.970 ;
        RECT 44.710 76.415 44.965 76.985 ;
        RECT 45.135 76.815 46.065 76.985 ;
        RECT 46.235 77.775 47.245 77.945 ;
        RECT 46.235 76.975 46.405 77.775 ;
        RECT 46.610 77.435 46.885 77.575 ;
        RECT 46.605 77.265 46.885 77.435 ;
        RECT 45.890 76.780 46.065 76.815 ;
        RECT 45.135 76.245 45.465 76.645 ;
        RECT 45.890 76.415 46.420 76.780 ;
        RECT 46.610 76.415 46.885 77.265 ;
        RECT 47.055 76.415 47.245 77.775 ;
        RECT 47.415 77.790 47.585 78.455 ;
        RECT 47.755 78.035 47.925 78.795 ;
        RECT 48.160 78.035 48.675 78.445 ;
        RECT 47.415 77.600 48.165 77.790 ;
        RECT 48.335 77.225 48.675 78.035 ;
        RECT 48.845 77.705 50.515 78.795 ;
        RECT 47.445 77.055 48.675 77.225 ;
        RECT 47.425 76.245 47.935 76.780 ;
        RECT 48.155 76.450 48.400 77.055 ;
        RECT 48.845 77.015 49.595 77.535 ;
        RECT 49.765 77.185 50.515 77.705 ;
        RECT 51.145 77.655 51.415 78.625 ;
        RECT 51.625 77.995 51.905 78.795 ;
        RECT 52.075 78.285 53.730 78.575 ;
        RECT 53.905 78.360 59.250 78.795 ;
        RECT 59.425 78.360 64.770 78.795 ;
        RECT 52.140 77.945 53.730 78.115 ;
        RECT 52.140 77.825 52.310 77.945 ;
        RECT 51.585 77.655 52.310 77.825 ;
        RECT 48.845 76.245 50.515 77.015 ;
        RECT 51.145 76.920 51.315 77.655 ;
        RECT 51.585 77.485 51.755 77.655 ;
        RECT 51.485 77.155 51.755 77.485 ;
        RECT 51.925 77.155 52.330 77.485 ;
        RECT 52.500 77.155 53.210 77.775 ;
        RECT 53.410 77.655 53.730 77.945 ;
        RECT 51.585 76.985 51.755 77.155 ;
        RECT 51.145 76.575 51.415 76.920 ;
        RECT 51.585 76.815 53.195 76.985 ;
        RECT 53.380 76.915 53.730 77.485 ;
        RECT 51.605 76.245 51.985 76.645 ;
        RECT 52.155 76.465 52.325 76.815 ;
        RECT 52.495 76.245 52.825 76.645 ;
        RECT 53.025 76.465 53.195 76.815 ;
        RECT 55.490 76.790 55.830 77.620 ;
        RECT 57.310 77.110 57.660 78.360 ;
        RECT 61.010 76.790 61.350 77.620 ;
        RECT 62.830 77.110 63.180 78.360 ;
        RECT 65.410 77.655 65.745 78.625 ;
        RECT 65.915 77.655 66.085 78.795 ;
        RECT 66.255 78.455 68.285 78.625 ;
        RECT 65.410 76.985 65.580 77.655 ;
        RECT 66.255 77.485 66.425 78.455 ;
        RECT 65.750 77.155 66.005 77.485 ;
        RECT 66.230 77.155 66.425 77.485 ;
        RECT 66.595 78.115 67.720 78.285 ;
        RECT 65.835 76.985 66.005 77.155 ;
        RECT 66.595 76.985 66.765 78.115 ;
        RECT 53.395 76.245 53.725 76.745 ;
        RECT 53.905 76.245 59.250 76.790 ;
        RECT 59.425 76.245 64.770 76.790 ;
        RECT 65.410 76.415 65.665 76.985 ;
        RECT 65.835 76.815 66.765 76.985 ;
        RECT 66.935 77.775 67.945 77.945 ;
        RECT 66.935 76.975 67.105 77.775 ;
        RECT 67.310 77.435 67.585 77.575 ;
        RECT 67.305 77.265 67.585 77.435 ;
        RECT 66.590 76.780 66.765 76.815 ;
        RECT 65.835 76.245 66.165 76.645 ;
        RECT 66.590 76.415 67.120 76.780 ;
        RECT 67.310 76.415 67.585 77.265 ;
        RECT 67.755 76.415 67.945 77.775 ;
        RECT 68.115 77.790 68.285 78.455 ;
        RECT 68.455 78.035 68.625 78.795 ;
        RECT 68.860 78.035 69.375 78.445 ;
        RECT 68.115 77.600 68.865 77.790 ;
        RECT 69.035 77.225 69.375 78.035 ;
        RECT 70.005 77.630 70.295 78.795 ;
        RECT 70.465 77.705 73.055 78.795 ;
        RECT 68.145 77.055 69.375 77.225 ;
        RECT 68.125 76.245 68.635 76.780 ;
        RECT 68.855 76.450 69.100 77.055 ;
        RECT 70.465 77.015 71.675 77.535 ;
        RECT 71.845 77.185 73.055 77.705 ;
        RECT 73.745 77.655 73.955 78.795 ;
        RECT 74.125 77.645 74.455 78.625 ;
        RECT 74.625 77.655 74.855 78.795 ;
        RECT 75.065 77.705 76.735 78.795 ;
        RECT 70.005 76.245 70.295 76.970 ;
        RECT 70.465 76.245 73.055 77.015 ;
        RECT 73.745 76.245 73.955 77.065 ;
        RECT 74.125 77.045 74.375 77.645 ;
        RECT 74.545 77.235 74.875 77.485 ;
        RECT 74.125 76.415 74.455 77.045 ;
        RECT 74.625 76.245 74.855 77.065 ;
        RECT 75.065 77.015 75.815 77.535 ;
        RECT 75.985 77.185 76.735 77.705 ;
        RECT 77.365 78.035 77.880 78.445 ;
        RECT 78.115 78.035 78.285 78.795 ;
        RECT 78.455 78.455 80.485 78.625 ;
        RECT 77.365 77.225 77.705 78.035 ;
        RECT 78.455 77.790 78.625 78.455 ;
        RECT 79.020 78.115 80.145 78.285 ;
        RECT 77.875 77.600 78.625 77.790 ;
        RECT 78.795 77.775 79.805 77.945 ;
        RECT 77.365 77.055 78.595 77.225 ;
        RECT 75.065 76.245 76.735 77.015 ;
        RECT 77.640 76.450 77.885 77.055 ;
        RECT 78.105 76.245 78.615 76.780 ;
        RECT 78.795 76.415 78.985 77.775 ;
        RECT 79.155 76.755 79.430 77.575 ;
        RECT 79.635 76.975 79.805 77.775 ;
        RECT 79.975 76.985 80.145 78.115 ;
        RECT 80.315 77.485 80.485 78.455 ;
        RECT 80.655 77.655 80.825 78.795 ;
        RECT 80.995 77.655 81.330 78.625 ;
        RECT 81.595 78.125 81.765 78.625 ;
        RECT 81.935 78.295 82.265 78.795 ;
        RECT 81.595 77.955 82.260 78.125 ;
        RECT 80.315 77.155 80.510 77.485 ;
        RECT 80.735 77.155 80.990 77.485 ;
        RECT 80.735 76.985 80.905 77.155 ;
        RECT 81.160 76.985 81.330 77.655 ;
        RECT 81.510 77.135 81.860 77.785 ;
        RECT 79.975 76.815 80.905 76.985 ;
        RECT 79.975 76.780 80.150 76.815 ;
        RECT 79.155 76.585 79.435 76.755 ;
        RECT 79.155 76.415 79.430 76.585 ;
        RECT 79.620 76.415 80.150 76.780 ;
        RECT 80.575 76.245 80.905 76.645 ;
        RECT 81.075 76.415 81.330 76.985 ;
        RECT 82.030 76.965 82.260 77.955 ;
        RECT 81.595 76.795 82.260 76.965 ;
        RECT 81.595 76.505 81.765 76.795 ;
        RECT 81.935 76.245 82.265 76.625 ;
        RECT 82.435 76.505 82.660 78.625 ;
        RECT 82.875 78.295 83.205 78.795 ;
        RECT 83.375 78.125 83.545 78.625 ;
        RECT 83.780 78.410 84.610 78.580 ;
        RECT 84.850 78.415 85.230 78.795 ;
        RECT 82.850 77.955 83.545 78.125 ;
        RECT 82.850 76.985 83.020 77.955 ;
        RECT 83.190 77.165 83.600 77.785 ;
        RECT 83.770 77.735 84.270 78.115 ;
        RECT 82.850 76.795 83.545 76.985 ;
        RECT 83.770 76.865 83.990 77.735 ;
        RECT 84.440 77.565 84.610 78.410 ;
        RECT 85.410 78.245 85.580 78.535 ;
        RECT 85.750 78.415 86.080 78.795 ;
        RECT 86.550 78.325 87.180 78.575 ;
        RECT 87.360 78.415 87.780 78.795 ;
        RECT 87.010 78.245 87.180 78.325 ;
        RECT 87.980 78.245 88.220 78.535 ;
        RECT 84.780 77.995 86.150 78.245 ;
        RECT 84.780 77.735 85.030 77.995 ;
        RECT 85.540 77.565 85.790 77.725 ;
        RECT 84.440 77.395 85.790 77.565 ;
        RECT 84.440 77.355 84.860 77.395 ;
        RECT 84.170 76.805 84.520 77.175 ;
        RECT 82.875 76.245 83.205 76.625 ;
        RECT 83.375 76.465 83.545 76.795 ;
        RECT 84.690 76.625 84.860 77.355 ;
        RECT 85.960 77.225 86.150 77.995 ;
        RECT 85.030 76.895 85.440 77.225 ;
        RECT 85.730 76.885 86.150 77.225 ;
        RECT 86.320 77.815 86.840 78.125 ;
        RECT 87.010 78.075 88.220 78.245 ;
        RECT 88.450 78.105 88.780 78.795 ;
        RECT 86.320 77.055 86.490 77.815 ;
        RECT 86.660 77.225 86.840 77.635 ;
        RECT 87.010 77.565 87.180 78.075 ;
        RECT 88.950 77.925 89.120 78.535 ;
        RECT 89.390 78.075 89.720 78.585 ;
        RECT 88.950 77.905 89.270 77.925 ;
        RECT 87.350 77.735 89.270 77.905 ;
        RECT 87.010 77.395 88.910 77.565 ;
        RECT 87.240 77.055 87.570 77.175 ;
        RECT 86.320 76.885 87.570 77.055 ;
        RECT 83.845 76.425 84.860 76.625 ;
        RECT 85.030 76.245 85.440 76.685 ;
        RECT 85.730 76.455 85.980 76.885 ;
        RECT 86.180 76.245 86.500 76.705 ;
        RECT 87.740 76.635 87.910 77.395 ;
        RECT 88.580 77.335 88.910 77.395 ;
        RECT 88.100 77.165 88.430 77.225 ;
        RECT 88.100 76.895 88.760 77.165 ;
        RECT 89.080 76.840 89.270 77.735 ;
        RECT 87.060 76.465 87.910 76.635 ;
        RECT 88.110 76.245 88.770 76.725 ;
        RECT 88.950 76.510 89.270 76.840 ;
        RECT 89.470 77.485 89.720 78.075 ;
        RECT 89.900 77.995 90.185 78.795 ;
        RECT 90.365 77.815 90.620 78.485 ;
        RECT 90.440 77.775 90.620 77.815 ;
        RECT 90.440 77.605 90.705 77.775 ;
        RECT 91.225 77.655 91.435 78.795 ;
        RECT 91.605 77.645 91.935 78.625 ;
        RECT 92.105 77.655 92.335 78.795 ;
        RECT 92.545 77.705 95.135 78.795 ;
        RECT 89.470 77.155 90.270 77.485 ;
        RECT 89.470 76.505 89.720 77.155 ;
        RECT 90.440 76.955 90.620 77.605 ;
        RECT 89.900 76.245 90.185 76.705 ;
        RECT 90.365 76.425 90.620 76.955 ;
        RECT 91.225 76.245 91.435 77.065 ;
        RECT 91.605 77.045 91.855 77.645 ;
        RECT 92.025 77.235 92.355 77.485 ;
        RECT 91.605 76.415 91.935 77.045 ;
        RECT 92.105 76.245 92.335 77.065 ;
        RECT 92.545 77.015 93.755 77.535 ;
        RECT 93.925 77.185 95.135 77.705 ;
        RECT 95.765 77.630 96.055 78.795 ;
        RECT 96.225 77.705 99.735 78.795 ;
        RECT 99.905 77.705 101.115 78.795 ;
        RECT 101.375 78.125 101.545 78.625 ;
        RECT 101.715 78.295 102.045 78.795 ;
        RECT 101.375 77.955 102.040 78.125 ;
        RECT 96.225 77.015 97.875 77.535 ;
        RECT 98.045 77.185 99.735 77.705 ;
        RECT 92.545 76.245 95.135 77.015 ;
        RECT 95.765 76.245 96.055 76.970 ;
        RECT 96.225 76.245 99.735 77.015 ;
        RECT 99.905 76.995 100.425 77.535 ;
        RECT 100.595 77.165 101.115 77.705 ;
        RECT 101.290 77.135 101.640 77.785 ;
        RECT 99.905 76.245 101.115 76.995 ;
        RECT 101.810 76.965 102.040 77.955 ;
        RECT 101.375 76.795 102.040 76.965 ;
        RECT 101.375 76.505 101.545 76.795 ;
        RECT 101.715 76.245 102.045 76.625 ;
        RECT 102.215 76.505 102.440 78.625 ;
        RECT 102.655 78.295 102.985 78.795 ;
        RECT 103.155 78.125 103.325 78.625 ;
        RECT 103.560 78.410 104.390 78.580 ;
        RECT 104.630 78.415 105.010 78.795 ;
        RECT 102.630 77.955 103.325 78.125 ;
        RECT 102.630 76.985 102.800 77.955 ;
        RECT 102.970 77.165 103.380 77.785 ;
        RECT 103.550 77.735 104.050 78.115 ;
        RECT 102.630 76.795 103.325 76.985 ;
        RECT 103.550 76.865 103.770 77.735 ;
        RECT 104.220 77.565 104.390 78.410 ;
        RECT 105.190 78.245 105.360 78.535 ;
        RECT 105.530 78.415 105.860 78.795 ;
        RECT 106.330 78.325 106.960 78.575 ;
        RECT 107.140 78.415 107.560 78.795 ;
        RECT 106.790 78.245 106.960 78.325 ;
        RECT 107.760 78.245 108.000 78.535 ;
        RECT 104.560 77.995 105.930 78.245 ;
        RECT 104.560 77.735 104.810 77.995 ;
        RECT 105.320 77.565 105.570 77.725 ;
        RECT 104.220 77.395 105.570 77.565 ;
        RECT 104.220 77.355 104.640 77.395 ;
        RECT 103.950 76.805 104.300 77.175 ;
        RECT 102.655 76.245 102.985 76.625 ;
        RECT 103.155 76.465 103.325 76.795 ;
        RECT 104.470 76.625 104.640 77.355 ;
        RECT 105.740 77.225 105.930 77.995 ;
        RECT 104.810 76.895 105.220 77.225 ;
        RECT 105.510 76.885 105.930 77.225 ;
        RECT 106.100 77.815 106.620 78.125 ;
        RECT 106.790 78.075 108.000 78.245 ;
        RECT 108.230 78.105 108.560 78.795 ;
        RECT 106.100 77.055 106.270 77.815 ;
        RECT 106.440 77.225 106.620 77.635 ;
        RECT 106.790 77.565 106.960 78.075 ;
        RECT 108.730 77.925 108.900 78.535 ;
        RECT 109.170 78.075 109.500 78.585 ;
        RECT 108.730 77.905 109.050 77.925 ;
        RECT 107.130 77.735 109.050 77.905 ;
        RECT 106.790 77.395 108.690 77.565 ;
        RECT 107.020 77.055 107.350 77.175 ;
        RECT 106.100 76.885 107.350 77.055 ;
        RECT 103.625 76.425 104.640 76.625 ;
        RECT 104.810 76.245 105.220 76.685 ;
        RECT 105.510 76.455 105.760 76.885 ;
        RECT 105.960 76.245 106.280 76.705 ;
        RECT 107.520 76.635 107.690 77.395 ;
        RECT 108.360 77.335 108.690 77.395 ;
        RECT 107.880 77.165 108.210 77.225 ;
        RECT 107.880 76.895 108.540 77.165 ;
        RECT 108.860 76.840 109.050 77.735 ;
        RECT 106.840 76.465 107.690 76.635 ;
        RECT 107.890 76.245 108.550 76.725 ;
        RECT 108.730 76.510 109.050 76.840 ;
        RECT 109.250 77.485 109.500 78.075 ;
        RECT 109.680 77.995 109.965 78.795 ;
        RECT 110.145 77.815 110.400 78.485 ;
        RECT 109.250 77.155 110.050 77.485 ;
        RECT 109.250 76.505 109.500 77.155 ;
        RECT 110.220 76.955 110.400 77.815 ;
        RECT 111.005 77.655 111.215 78.795 ;
        RECT 111.385 77.645 111.715 78.625 ;
        RECT 111.885 77.655 112.115 78.795 ;
        RECT 112.385 77.655 112.595 78.795 ;
        RECT 112.765 77.645 113.095 78.625 ;
        RECT 113.265 77.655 113.495 78.795 ;
        RECT 113.705 77.705 117.215 78.795 ;
        RECT 110.145 76.755 110.400 76.955 ;
        RECT 109.680 76.245 109.965 76.705 ;
        RECT 110.145 76.585 110.485 76.755 ;
        RECT 110.145 76.425 110.400 76.585 ;
        RECT 111.005 76.245 111.215 77.065 ;
        RECT 111.385 77.045 111.635 77.645 ;
        RECT 111.805 77.235 112.135 77.485 ;
        RECT 111.385 76.415 111.715 77.045 ;
        RECT 111.885 76.245 112.115 77.065 ;
        RECT 112.385 76.245 112.595 77.065 ;
        RECT 112.765 77.045 113.015 77.645 ;
        RECT 113.185 77.235 113.515 77.485 ;
        RECT 112.765 76.415 113.095 77.045 ;
        RECT 113.265 76.245 113.495 77.065 ;
        RECT 113.705 77.015 115.355 77.535 ;
        RECT 115.525 77.185 117.215 77.705 ;
        RECT 117.385 77.705 118.595 78.795 ;
        RECT 117.385 77.165 117.905 77.705 ;
        RECT 113.705 76.245 117.215 77.015 ;
        RECT 118.075 76.995 118.595 77.535 ;
        RECT 117.385 76.245 118.595 76.995 ;
        RECT 5.520 76.075 118.680 76.245 ;
        RECT 5.605 75.325 6.815 76.075 ;
        RECT 7.535 75.525 7.705 75.815 ;
        RECT 7.875 75.695 8.205 76.075 ;
        RECT 7.535 75.355 8.200 75.525 ;
        RECT 5.605 74.785 6.125 75.325 ;
        RECT 6.295 74.615 6.815 75.155 ;
        RECT 5.605 73.525 6.815 74.615 ;
        RECT 7.450 74.535 7.800 75.185 ;
        RECT 7.970 74.365 8.200 75.355 ;
        RECT 7.535 74.195 8.200 74.365 ;
        RECT 7.535 73.695 7.705 74.195 ;
        RECT 7.875 73.525 8.205 74.025 ;
        RECT 8.375 73.695 8.600 75.815 ;
        RECT 8.815 75.695 9.145 76.075 ;
        RECT 9.315 75.525 9.485 75.855 ;
        RECT 9.785 75.695 10.800 75.895 ;
        RECT 8.790 75.335 9.485 75.525 ;
        RECT 8.790 74.365 8.960 75.335 ;
        RECT 9.130 74.535 9.540 75.155 ;
        RECT 9.710 74.585 9.930 75.455 ;
        RECT 10.110 75.145 10.460 75.515 ;
        RECT 10.630 74.965 10.800 75.695 ;
        RECT 10.970 75.635 11.380 76.075 ;
        RECT 11.670 75.435 11.920 75.865 ;
        RECT 12.120 75.615 12.440 76.075 ;
        RECT 13.000 75.685 13.850 75.855 ;
        RECT 10.970 75.095 11.380 75.425 ;
        RECT 11.670 75.095 12.090 75.435 ;
        RECT 10.380 74.925 10.800 74.965 ;
        RECT 10.380 74.755 11.730 74.925 ;
        RECT 8.790 74.195 9.485 74.365 ;
        RECT 9.710 74.205 10.210 74.585 ;
        RECT 8.815 73.525 9.145 74.025 ;
        RECT 9.315 73.695 9.485 74.195 ;
        RECT 10.380 73.910 10.550 74.755 ;
        RECT 11.480 74.595 11.730 74.755 ;
        RECT 10.720 74.325 10.970 74.585 ;
        RECT 11.900 74.325 12.090 75.095 ;
        RECT 10.720 74.075 12.090 74.325 ;
        RECT 12.260 75.265 13.510 75.435 ;
        RECT 12.260 74.505 12.430 75.265 ;
        RECT 13.180 75.145 13.510 75.265 ;
        RECT 12.600 74.685 12.780 75.095 ;
        RECT 13.680 74.925 13.850 75.685 ;
        RECT 14.050 75.595 14.710 76.075 ;
        RECT 14.890 75.480 15.210 75.810 ;
        RECT 14.040 75.155 14.700 75.425 ;
        RECT 14.040 75.095 14.370 75.155 ;
        RECT 14.520 74.925 14.850 74.985 ;
        RECT 12.950 74.755 14.850 74.925 ;
        RECT 12.260 74.195 12.780 74.505 ;
        RECT 12.950 74.245 13.120 74.755 ;
        RECT 15.020 74.585 15.210 75.480 ;
        RECT 13.290 74.415 15.210 74.585 ;
        RECT 14.890 74.395 15.210 74.415 ;
        RECT 15.410 75.165 15.660 75.815 ;
        RECT 15.840 75.615 16.125 76.075 ;
        RECT 16.305 75.395 16.560 75.895 ;
        RECT 16.305 75.365 16.645 75.395 ;
        RECT 16.380 75.225 16.645 75.365 ;
        RECT 17.110 75.335 17.365 75.905 ;
        RECT 17.535 75.675 17.865 76.075 ;
        RECT 18.290 75.540 18.820 75.905 ;
        RECT 18.290 75.505 18.465 75.540 ;
        RECT 17.535 75.335 18.465 75.505 ;
        RECT 15.410 74.835 16.210 75.165 ;
        RECT 12.950 74.075 14.160 74.245 ;
        RECT 9.720 73.740 10.550 73.910 ;
        RECT 10.790 73.525 11.170 73.905 ;
        RECT 11.350 73.785 11.520 74.075 ;
        RECT 12.950 73.995 13.120 74.075 ;
        RECT 11.690 73.525 12.020 73.905 ;
        RECT 12.490 73.745 13.120 73.995 ;
        RECT 13.300 73.525 13.720 73.905 ;
        RECT 13.920 73.785 14.160 74.075 ;
        RECT 14.390 73.525 14.720 74.215 ;
        RECT 14.890 73.785 15.060 74.395 ;
        RECT 15.410 74.245 15.660 74.835 ;
        RECT 16.380 74.505 16.560 75.225 ;
        RECT 15.330 73.735 15.660 74.245 ;
        RECT 15.840 73.525 16.125 74.325 ;
        RECT 16.305 73.835 16.560 74.505 ;
        RECT 17.110 74.665 17.280 75.335 ;
        RECT 17.535 75.165 17.705 75.335 ;
        RECT 17.450 74.835 17.705 75.165 ;
        RECT 17.930 74.835 18.125 75.165 ;
        RECT 17.110 73.695 17.445 74.665 ;
        RECT 17.615 73.525 17.785 74.665 ;
        RECT 17.955 73.865 18.125 74.835 ;
        RECT 18.295 74.205 18.465 75.335 ;
        RECT 18.635 74.545 18.805 75.345 ;
        RECT 19.010 75.055 19.285 75.905 ;
        RECT 19.005 74.885 19.285 75.055 ;
        RECT 19.010 74.745 19.285 74.885 ;
        RECT 19.455 74.545 19.645 75.905 ;
        RECT 19.825 75.540 20.335 76.075 ;
        RECT 20.555 75.265 20.800 75.870 ;
        RECT 21.245 75.305 22.915 76.075 ;
        RECT 19.845 75.095 21.075 75.265 ;
        RECT 18.635 74.375 19.645 74.545 ;
        RECT 19.815 74.530 20.565 74.720 ;
        RECT 18.295 74.035 19.420 74.205 ;
        RECT 19.815 73.865 19.985 74.530 ;
        RECT 20.735 74.285 21.075 75.095 ;
        RECT 21.245 74.785 21.995 75.305 ;
        RECT 23.290 75.295 23.790 75.905 ;
        RECT 22.165 74.615 22.915 75.135 ;
        RECT 23.085 74.835 23.435 75.085 ;
        RECT 23.620 74.665 23.790 75.295 ;
        RECT 24.420 75.425 24.750 75.905 ;
        RECT 24.920 75.615 25.145 76.075 ;
        RECT 25.315 75.425 25.645 75.905 ;
        RECT 24.420 75.255 25.645 75.425 ;
        RECT 25.835 75.275 26.085 76.075 ;
        RECT 26.255 75.275 26.595 75.905 ;
        RECT 26.775 75.575 27.105 76.075 ;
        RECT 27.305 75.505 27.475 75.855 ;
        RECT 27.675 75.675 28.005 76.075 ;
        RECT 28.175 75.505 28.345 75.855 ;
        RECT 28.515 75.675 28.895 76.075 ;
        RECT 26.365 75.225 26.595 75.275 ;
        RECT 23.960 74.885 24.290 75.085 ;
        RECT 24.460 74.885 24.790 75.085 ;
        RECT 24.960 74.885 25.380 75.085 ;
        RECT 25.555 74.915 26.250 75.085 ;
        RECT 25.555 74.665 25.725 74.915 ;
        RECT 26.420 74.665 26.595 75.225 ;
        RECT 26.770 74.835 27.120 75.405 ;
        RECT 27.305 75.335 28.915 75.505 ;
        RECT 29.085 75.400 29.355 75.745 ;
        RECT 28.745 75.165 28.915 75.335 ;
        RECT 27.290 74.715 28.000 75.165 ;
        RECT 28.170 74.835 28.575 75.165 ;
        RECT 28.745 74.835 29.015 75.165 ;
        RECT 17.955 73.695 19.985 73.865 ;
        RECT 20.155 73.525 20.325 74.285 ;
        RECT 20.560 73.875 21.075 74.285 ;
        RECT 21.245 73.525 22.915 74.615 ;
        RECT 23.290 74.495 25.725 74.665 ;
        RECT 23.290 73.695 23.620 74.495 ;
        RECT 23.790 73.525 24.120 74.325 ;
        RECT 24.420 73.695 24.750 74.495 ;
        RECT 25.395 73.525 25.645 74.325 ;
        RECT 25.915 73.525 26.085 74.665 ;
        RECT 26.255 73.695 26.595 74.665 ;
        RECT 26.770 74.375 27.090 74.665 ;
        RECT 27.285 74.545 28.000 74.715 ;
        RECT 28.745 74.665 28.915 74.835 ;
        RECT 29.185 74.665 29.355 75.400 ;
        RECT 28.190 74.495 28.915 74.665 ;
        RECT 28.190 74.375 28.360 74.495 ;
        RECT 26.770 74.205 28.360 74.375 ;
        RECT 26.770 73.745 28.425 74.035 ;
        RECT 28.595 73.525 28.875 74.325 ;
        RECT 29.085 73.695 29.355 74.665 ;
        RECT 29.985 75.400 30.245 75.905 ;
        RECT 30.425 75.695 30.755 76.075 ;
        RECT 30.935 75.525 31.105 75.905 ;
        RECT 29.985 74.600 30.155 75.400 ;
        RECT 30.440 75.355 31.105 75.525 ;
        RECT 30.440 75.100 30.610 75.355 ;
        RECT 31.365 75.350 31.655 76.075 ;
        RECT 32.750 75.335 33.005 75.905 ;
        RECT 33.175 75.675 33.505 76.075 ;
        RECT 33.930 75.540 34.460 75.905 ;
        RECT 33.930 75.505 34.105 75.540 ;
        RECT 33.175 75.335 34.105 75.505 ;
        RECT 30.325 74.770 30.610 75.100 ;
        RECT 30.845 74.805 31.175 75.175 ;
        RECT 30.440 74.625 30.610 74.770 ;
        RECT 29.985 73.695 30.255 74.600 ;
        RECT 30.440 74.455 31.105 74.625 ;
        RECT 30.425 73.525 30.755 74.285 ;
        RECT 30.935 73.695 31.105 74.455 ;
        RECT 31.365 73.525 31.655 74.690 ;
        RECT 32.750 74.665 32.920 75.335 ;
        RECT 33.175 75.165 33.345 75.335 ;
        RECT 33.090 74.835 33.345 75.165 ;
        RECT 33.570 74.835 33.765 75.165 ;
        RECT 32.750 73.695 33.085 74.665 ;
        RECT 33.255 73.525 33.425 74.665 ;
        RECT 33.595 73.865 33.765 74.835 ;
        RECT 33.935 74.205 34.105 75.335 ;
        RECT 34.275 74.545 34.445 75.345 ;
        RECT 34.650 75.055 34.925 75.905 ;
        RECT 34.645 74.885 34.925 75.055 ;
        RECT 34.650 74.745 34.925 74.885 ;
        RECT 35.095 74.545 35.285 75.905 ;
        RECT 35.465 75.540 35.975 76.075 ;
        RECT 36.195 75.265 36.440 75.870 ;
        RECT 35.485 75.095 36.715 75.265 ;
        RECT 36.945 75.255 37.155 76.075 ;
        RECT 37.325 75.275 37.655 75.905 ;
        RECT 34.275 74.375 35.285 74.545 ;
        RECT 35.455 74.530 36.205 74.720 ;
        RECT 33.935 74.035 35.060 74.205 ;
        RECT 35.455 73.865 35.625 74.530 ;
        RECT 36.375 74.285 36.715 75.095 ;
        RECT 37.325 74.675 37.575 75.275 ;
        RECT 37.825 75.255 38.055 76.075 ;
        RECT 38.815 75.525 38.985 75.815 ;
        RECT 39.155 75.695 39.485 76.075 ;
        RECT 38.815 75.355 39.480 75.525 ;
        RECT 37.745 74.835 38.075 75.085 ;
        RECT 33.595 73.695 35.625 73.865 ;
        RECT 35.795 73.525 35.965 74.285 ;
        RECT 36.200 73.875 36.715 74.285 ;
        RECT 36.945 73.525 37.155 74.665 ;
        RECT 37.325 73.695 37.655 74.675 ;
        RECT 37.825 73.525 38.055 74.665 ;
        RECT 38.730 74.535 39.080 75.185 ;
        RECT 39.250 74.365 39.480 75.355 ;
        RECT 38.815 74.195 39.480 74.365 ;
        RECT 38.815 73.695 38.985 74.195 ;
        RECT 39.155 73.525 39.485 74.025 ;
        RECT 39.655 73.695 39.880 75.815 ;
        RECT 40.095 75.695 40.425 76.075 ;
        RECT 40.595 75.525 40.765 75.855 ;
        RECT 41.065 75.695 42.080 75.895 ;
        RECT 40.070 75.335 40.765 75.525 ;
        RECT 40.070 74.365 40.240 75.335 ;
        RECT 40.410 74.535 40.820 75.155 ;
        RECT 40.990 74.585 41.210 75.455 ;
        RECT 41.390 75.145 41.740 75.515 ;
        RECT 41.910 74.965 42.080 75.695 ;
        RECT 42.250 75.635 42.660 76.075 ;
        RECT 42.950 75.435 43.200 75.865 ;
        RECT 43.400 75.615 43.720 76.075 ;
        RECT 44.280 75.685 45.130 75.855 ;
        RECT 42.250 75.095 42.660 75.425 ;
        RECT 42.950 75.095 43.370 75.435 ;
        RECT 41.660 74.925 42.080 74.965 ;
        RECT 41.660 74.755 43.010 74.925 ;
        RECT 40.070 74.195 40.765 74.365 ;
        RECT 40.990 74.205 41.490 74.585 ;
        RECT 40.095 73.525 40.425 74.025 ;
        RECT 40.595 73.695 40.765 74.195 ;
        RECT 41.660 73.910 41.830 74.755 ;
        RECT 42.760 74.595 43.010 74.755 ;
        RECT 42.000 74.325 42.250 74.585 ;
        RECT 43.180 74.325 43.370 75.095 ;
        RECT 42.000 74.075 43.370 74.325 ;
        RECT 43.540 75.265 44.790 75.435 ;
        RECT 43.540 74.505 43.710 75.265 ;
        RECT 44.460 75.145 44.790 75.265 ;
        RECT 43.880 74.685 44.060 75.095 ;
        RECT 44.960 74.925 45.130 75.685 ;
        RECT 45.330 75.595 45.990 76.075 ;
        RECT 46.170 75.480 46.490 75.810 ;
        RECT 45.320 75.155 45.980 75.425 ;
        RECT 45.320 75.095 45.650 75.155 ;
        RECT 45.800 74.925 46.130 74.985 ;
        RECT 44.230 74.755 46.130 74.925 ;
        RECT 43.540 74.195 44.060 74.505 ;
        RECT 44.230 74.245 44.400 74.755 ;
        RECT 46.300 74.585 46.490 75.480 ;
        RECT 44.570 74.415 46.490 74.585 ;
        RECT 46.170 74.395 46.490 74.415 ;
        RECT 46.690 75.165 46.940 75.815 ;
        RECT 47.120 75.615 47.405 76.075 ;
        RECT 47.585 75.735 47.840 75.895 ;
        RECT 47.585 75.565 47.925 75.735 ;
        RECT 47.585 75.365 47.840 75.565 ;
        RECT 46.690 74.835 47.490 75.165 ;
        RECT 44.230 74.075 45.440 74.245 ;
        RECT 41.000 73.740 41.830 73.910 ;
        RECT 42.070 73.525 42.450 73.905 ;
        RECT 42.630 73.785 42.800 74.075 ;
        RECT 44.230 73.995 44.400 74.075 ;
        RECT 42.970 73.525 43.300 73.905 ;
        RECT 43.770 73.745 44.400 73.995 ;
        RECT 44.580 73.525 45.000 73.905 ;
        RECT 45.200 73.785 45.440 74.075 ;
        RECT 45.670 73.525 46.000 74.215 ;
        RECT 46.170 73.785 46.340 74.395 ;
        RECT 46.690 74.245 46.940 74.835 ;
        RECT 47.660 74.505 47.840 75.365 ;
        RECT 48.385 75.325 49.595 76.075 ;
        RECT 48.385 74.785 48.905 75.325 ;
        RECT 49.970 75.295 50.470 75.905 ;
        RECT 49.075 74.615 49.595 75.155 ;
        RECT 49.765 74.835 50.115 75.085 ;
        RECT 50.300 74.665 50.470 75.295 ;
        RECT 51.100 75.425 51.430 75.905 ;
        RECT 51.600 75.615 51.825 76.075 ;
        RECT 51.995 75.425 52.325 75.905 ;
        RECT 51.100 75.255 52.325 75.425 ;
        RECT 52.515 75.275 52.765 76.075 ;
        RECT 52.935 75.275 53.275 75.905 ;
        RECT 50.640 74.885 50.970 75.085 ;
        RECT 51.140 74.885 51.470 75.085 ;
        RECT 51.640 74.885 52.060 75.085 ;
        RECT 52.235 74.915 52.930 75.085 ;
        RECT 52.235 74.665 52.405 74.915 ;
        RECT 53.100 74.665 53.275 75.275 ;
        RECT 46.610 73.735 46.940 74.245 ;
        RECT 47.120 73.525 47.405 74.325 ;
        RECT 47.585 73.835 47.840 74.505 ;
        RECT 48.385 73.525 49.595 74.615 ;
        RECT 49.970 74.495 52.405 74.665 ;
        RECT 49.970 73.695 50.300 74.495 ;
        RECT 50.470 73.525 50.800 74.325 ;
        RECT 51.100 73.695 51.430 74.495 ;
        RECT 52.075 73.525 52.325 74.325 ;
        RECT 52.595 73.525 52.765 74.665 ;
        RECT 52.935 73.695 53.275 74.665 ;
        RECT 53.445 75.275 53.785 75.905 ;
        RECT 53.955 75.275 54.205 76.075 ;
        RECT 54.395 75.425 54.725 75.905 ;
        RECT 54.895 75.615 55.120 76.075 ;
        RECT 55.290 75.425 55.620 75.905 ;
        RECT 53.445 74.665 53.620 75.275 ;
        RECT 54.395 75.255 55.620 75.425 ;
        RECT 56.250 75.295 56.750 75.905 ;
        RECT 57.125 75.350 57.415 76.075 ;
        RECT 57.585 75.325 58.795 76.075 ;
        RECT 53.790 74.915 54.485 75.085 ;
        RECT 54.315 74.665 54.485 74.915 ;
        RECT 54.660 74.885 55.080 75.085 ;
        RECT 55.250 74.885 55.580 75.085 ;
        RECT 55.750 74.885 56.080 75.085 ;
        RECT 56.250 74.665 56.420 75.295 ;
        RECT 56.605 74.835 56.955 75.085 ;
        RECT 57.585 74.785 58.105 75.325 ;
        RECT 58.970 75.235 59.230 76.075 ;
        RECT 59.405 75.330 59.660 75.905 ;
        RECT 59.830 75.695 60.160 76.075 ;
        RECT 60.375 75.525 60.545 75.905 ;
        RECT 59.830 75.355 60.545 75.525 ;
        RECT 60.895 75.525 61.065 75.905 ;
        RECT 61.280 75.695 61.610 76.075 ;
        RECT 60.895 75.355 61.610 75.525 ;
        RECT 53.445 73.695 53.785 74.665 ;
        RECT 53.955 73.525 54.125 74.665 ;
        RECT 54.315 74.495 56.750 74.665 ;
        RECT 54.395 73.525 54.645 74.325 ;
        RECT 55.290 73.695 55.620 74.495 ;
        RECT 55.920 73.525 56.250 74.325 ;
        RECT 56.420 73.695 56.750 74.495 ;
        RECT 57.125 73.525 57.415 74.690 ;
        RECT 58.275 74.615 58.795 75.155 ;
        RECT 57.585 73.525 58.795 74.615 ;
        RECT 58.970 73.525 59.230 74.675 ;
        RECT 59.405 74.600 59.575 75.330 ;
        RECT 59.830 75.165 60.000 75.355 ;
        RECT 59.745 74.835 60.000 75.165 ;
        RECT 59.830 74.625 60.000 74.835 ;
        RECT 60.280 74.805 60.635 75.175 ;
        RECT 60.805 74.805 61.160 75.175 ;
        RECT 61.440 75.165 61.610 75.355 ;
        RECT 61.780 75.330 62.035 75.905 ;
        RECT 61.440 74.835 61.695 75.165 ;
        RECT 61.440 74.625 61.610 74.835 ;
        RECT 59.405 73.695 59.660 74.600 ;
        RECT 59.830 74.455 60.545 74.625 ;
        RECT 59.830 73.525 60.160 74.285 ;
        RECT 60.375 73.695 60.545 74.455 ;
        RECT 60.895 74.455 61.610 74.625 ;
        RECT 61.865 74.600 62.035 75.330 ;
        RECT 62.210 75.235 62.470 76.075 ;
        RECT 62.645 75.530 67.990 76.075 ;
        RECT 64.230 74.700 64.570 75.530 ;
        RECT 68.165 75.325 69.375 76.075 ;
        RECT 69.550 75.335 69.805 75.905 ;
        RECT 69.975 75.675 70.305 76.075 ;
        RECT 70.730 75.540 71.260 75.905 ;
        RECT 71.450 75.735 71.725 75.905 ;
        RECT 71.445 75.565 71.725 75.735 ;
        RECT 70.730 75.505 70.905 75.540 ;
        RECT 69.975 75.335 70.905 75.505 ;
        RECT 60.895 73.695 61.065 74.455 ;
        RECT 61.280 73.525 61.610 74.285 ;
        RECT 61.780 73.695 62.035 74.600 ;
        RECT 62.210 73.525 62.470 74.675 ;
        RECT 66.050 73.960 66.400 75.210 ;
        RECT 68.165 74.785 68.685 75.325 ;
        RECT 68.855 74.615 69.375 75.155 ;
        RECT 62.645 73.525 67.990 73.960 ;
        RECT 68.165 73.525 69.375 74.615 ;
        RECT 69.550 74.665 69.720 75.335 ;
        RECT 69.975 75.165 70.145 75.335 ;
        RECT 69.890 74.835 70.145 75.165 ;
        RECT 70.370 74.835 70.565 75.165 ;
        RECT 69.550 73.695 69.885 74.665 ;
        RECT 70.055 73.525 70.225 74.665 ;
        RECT 70.395 73.865 70.565 74.835 ;
        RECT 70.735 74.205 70.905 75.335 ;
        RECT 71.075 74.545 71.245 75.345 ;
        RECT 71.450 74.745 71.725 75.565 ;
        RECT 71.895 74.545 72.085 75.905 ;
        RECT 72.265 75.540 72.775 76.075 ;
        RECT 72.995 75.265 73.240 75.870 ;
        RECT 73.685 75.305 76.275 76.075 ;
        RECT 72.285 75.095 73.515 75.265 ;
        RECT 71.075 74.375 72.085 74.545 ;
        RECT 72.255 74.530 73.005 74.720 ;
        RECT 70.735 74.035 71.860 74.205 ;
        RECT 72.255 73.865 72.425 74.530 ;
        RECT 73.175 74.285 73.515 75.095 ;
        RECT 73.685 74.785 74.895 75.305 ;
        RECT 76.650 75.295 77.150 75.905 ;
        RECT 75.065 74.615 76.275 75.135 ;
        RECT 76.445 74.835 76.795 75.085 ;
        RECT 76.980 74.665 77.150 75.295 ;
        RECT 77.780 75.425 78.110 75.905 ;
        RECT 78.280 75.615 78.505 76.075 ;
        RECT 78.675 75.425 79.005 75.905 ;
        RECT 77.780 75.255 79.005 75.425 ;
        RECT 79.195 75.275 79.445 76.075 ;
        RECT 79.615 75.275 79.955 75.905 ;
        RECT 81.135 75.525 81.305 75.905 ;
        RECT 81.485 75.695 81.815 76.075 ;
        RECT 81.135 75.355 81.800 75.525 ;
        RECT 81.995 75.400 82.255 75.905 ;
        RECT 77.320 74.885 77.650 75.085 ;
        RECT 77.820 74.885 78.150 75.085 ;
        RECT 78.320 74.885 78.740 75.085 ;
        RECT 78.915 74.915 79.610 75.085 ;
        RECT 78.915 74.665 79.085 74.915 ;
        RECT 79.780 74.665 79.955 75.275 ;
        RECT 81.065 74.805 81.395 75.175 ;
        RECT 81.630 75.100 81.800 75.355 ;
        RECT 70.395 73.695 72.425 73.865 ;
        RECT 72.595 73.525 72.765 74.285 ;
        RECT 73.000 73.875 73.515 74.285 ;
        RECT 73.685 73.525 76.275 74.615 ;
        RECT 76.650 74.495 79.085 74.665 ;
        RECT 76.650 73.695 76.980 74.495 ;
        RECT 77.150 73.525 77.480 74.325 ;
        RECT 77.780 73.695 78.110 74.495 ;
        RECT 78.755 73.525 79.005 74.325 ;
        RECT 79.275 73.525 79.445 74.665 ;
        RECT 79.615 73.695 79.955 74.665 ;
        RECT 81.630 74.770 81.915 75.100 ;
        RECT 81.630 74.625 81.800 74.770 ;
        RECT 81.135 74.455 81.800 74.625 ;
        RECT 82.085 74.600 82.255 75.400 ;
        RECT 82.885 75.350 83.175 76.075 ;
        RECT 83.345 75.400 83.615 75.745 ;
        RECT 83.805 75.675 84.185 76.075 ;
        RECT 84.355 75.505 84.525 75.855 ;
        RECT 84.695 75.675 85.025 76.075 ;
        RECT 85.225 75.505 85.395 75.855 ;
        RECT 85.595 75.575 85.925 76.075 ;
        RECT 81.135 73.695 81.305 74.455 ;
        RECT 81.485 73.525 81.815 74.285 ;
        RECT 81.985 73.695 82.255 74.600 ;
        RECT 82.885 73.525 83.175 74.690 ;
        RECT 83.345 74.665 83.515 75.400 ;
        RECT 83.785 75.335 85.395 75.505 ;
        RECT 83.785 75.165 83.955 75.335 ;
        RECT 83.685 74.835 83.955 75.165 ;
        RECT 84.125 74.835 84.530 75.165 ;
        RECT 83.785 74.665 83.955 74.835 ;
        RECT 83.345 73.695 83.615 74.665 ;
        RECT 83.785 74.495 84.510 74.665 ;
        RECT 84.700 74.545 85.410 75.165 ;
        RECT 85.580 74.835 85.930 75.405 ;
        RECT 86.105 75.305 89.615 76.075 ;
        RECT 86.105 74.785 87.755 75.305 ;
        RECT 90.450 75.295 90.950 75.905 ;
        RECT 84.340 74.375 84.510 74.495 ;
        RECT 85.610 74.375 85.930 74.665 ;
        RECT 87.925 74.615 89.615 75.135 ;
        RECT 90.245 74.835 90.595 75.085 ;
        RECT 90.780 74.665 90.950 75.295 ;
        RECT 91.580 75.425 91.910 75.905 ;
        RECT 92.080 75.615 92.305 76.075 ;
        RECT 92.475 75.425 92.805 75.905 ;
        RECT 91.580 75.255 92.805 75.425 ;
        RECT 92.995 75.275 93.245 76.075 ;
        RECT 93.415 75.275 93.755 75.905 ;
        RECT 93.525 75.225 93.755 75.275 ;
        RECT 91.120 74.885 91.450 75.085 ;
        RECT 91.620 74.885 91.950 75.085 ;
        RECT 92.120 74.885 92.540 75.085 ;
        RECT 92.715 74.915 93.410 75.085 ;
        RECT 92.715 74.665 92.885 74.915 ;
        RECT 93.580 74.665 93.755 75.225 ;
        RECT 83.825 73.525 84.105 74.325 ;
        RECT 84.340 74.205 85.930 74.375 ;
        RECT 84.275 73.745 85.930 74.035 ;
        RECT 86.105 73.525 89.615 74.615 ;
        RECT 90.450 74.495 92.885 74.665 ;
        RECT 90.450 73.695 90.780 74.495 ;
        RECT 90.950 73.525 91.280 74.325 ;
        RECT 91.580 73.695 91.910 74.495 ;
        RECT 92.555 73.525 92.805 74.325 ;
        RECT 93.075 73.525 93.245 74.665 ;
        RECT 93.415 73.695 93.755 74.665 ;
        RECT 93.925 75.275 94.265 75.905 ;
        RECT 94.435 75.275 94.685 76.075 ;
        RECT 94.875 75.425 95.205 75.905 ;
        RECT 95.375 75.615 95.600 76.075 ;
        RECT 95.770 75.425 96.100 75.905 ;
        RECT 93.925 74.665 94.100 75.275 ;
        RECT 94.875 75.255 96.100 75.425 ;
        RECT 96.730 75.295 97.230 75.905 ;
        RECT 97.605 75.305 99.275 76.075 ;
        RECT 94.270 74.915 94.965 75.085 ;
        RECT 94.795 74.665 94.965 74.915 ;
        RECT 95.140 74.885 95.560 75.085 ;
        RECT 95.730 74.885 96.060 75.085 ;
        RECT 96.230 74.885 96.560 75.085 ;
        RECT 96.730 74.665 96.900 75.295 ;
        RECT 97.085 74.835 97.435 75.085 ;
        RECT 97.605 74.785 98.355 75.305 ;
        RECT 100.180 75.265 100.425 75.870 ;
        RECT 100.645 75.540 101.155 76.075 ;
        RECT 93.925 73.695 94.265 74.665 ;
        RECT 94.435 73.525 94.605 74.665 ;
        RECT 94.795 74.495 97.230 74.665 ;
        RECT 98.525 74.615 99.275 75.135 ;
        RECT 94.875 73.525 95.125 74.325 ;
        RECT 95.770 73.695 96.100 74.495 ;
        RECT 96.400 73.525 96.730 74.325 ;
        RECT 96.900 73.695 97.230 74.495 ;
        RECT 97.605 73.525 99.275 74.615 ;
        RECT 99.905 75.095 101.135 75.265 ;
        RECT 99.905 74.285 100.245 75.095 ;
        RECT 100.415 74.530 101.165 74.720 ;
        RECT 99.905 73.875 100.420 74.285 ;
        RECT 100.655 73.525 100.825 74.285 ;
        RECT 100.995 73.865 101.165 74.530 ;
        RECT 101.335 74.545 101.525 75.905 ;
        RECT 101.695 75.055 101.970 75.905 ;
        RECT 102.160 75.540 102.690 75.905 ;
        RECT 103.115 75.675 103.445 76.075 ;
        RECT 102.515 75.505 102.690 75.540 ;
        RECT 101.695 74.885 101.975 75.055 ;
        RECT 101.695 74.745 101.970 74.885 ;
        RECT 102.175 74.545 102.345 75.345 ;
        RECT 101.335 74.375 102.345 74.545 ;
        RECT 102.515 75.335 103.445 75.505 ;
        RECT 103.615 75.335 103.870 75.905 ;
        RECT 102.515 74.205 102.685 75.335 ;
        RECT 103.275 75.165 103.445 75.335 ;
        RECT 101.560 74.035 102.685 74.205 ;
        RECT 102.855 74.835 103.050 75.165 ;
        RECT 103.275 74.835 103.530 75.165 ;
        RECT 102.855 73.865 103.025 74.835 ;
        RECT 103.700 74.665 103.870 75.335 ;
        RECT 100.995 73.695 103.025 73.865 ;
        RECT 103.195 73.525 103.365 74.665 ;
        RECT 103.535 73.695 103.870 74.665 ;
        RECT 104.045 75.400 104.305 75.905 ;
        RECT 104.485 75.695 104.815 76.075 ;
        RECT 104.995 75.525 105.165 75.905 ;
        RECT 104.045 74.600 104.215 75.400 ;
        RECT 104.500 75.355 105.165 75.525 ;
        RECT 104.500 75.100 104.670 75.355 ;
        RECT 105.425 75.305 107.095 76.075 ;
        RECT 107.355 75.525 107.525 75.905 ;
        RECT 107.705 75.695 108.035 76.075 ;
        RECT 107.355 75.355 108.020 75.525 ;
        RECT 108.215 75.400 108.475 75.905 ;
        RECT 104.385 74.770 104.670 75.100 ;
        RECT 104.905 74.805 105.235 75.175 ;
        RECT 105.425 74.785 106.175 75.305 ;
        RECT 104.500 74.625 104.670 74.770 ;
        RECT 104.045 73.695 104.315 74.600 ;
        RECT 104.500 74.455 105.165 74.625 ;
        RECT 106.345 74.615 107.095 75.135 ;
        RECT 107.285 74.805 107.615 75.175 ;
        RECT 107.850 75.100 108.020 75.355 ;
        RECT 107.850 74.770 108.135 75.100 ;
        RECT 107.850 74.625 108.020 74.770 ;
        RECT 104.485 73.525 104.815 74.285 ;
        RECT 104.995 73.695 105.165 74.455 ;
        RECT 105.425 73.525 107.095 74.615 ;
        RECT 107.355 74.455 108.020 74.625 ;
        RECT 108.305 74.600 108.475 75.400 ;
        RECT 108.645 75.350 108.935 76.075 ;
        RECT 109.110 75.335 109.365 75.905 ;
        RECT 109.535 75.675 109.865 76.075 ;
        RECT 110.290 75.540 110.820 75.905 ;
        RECT 110.290 75.505 110.465 75.540 ;
        RECT 109.535 75.335 110.465 75.505 ;
        RECT 111.010 75.395 111.285 75.905 ;
        RECT 107.355 73.695 107.525 74.455 ;
        RECT 107.705 73.525 108.035 74.285 ;
        RECT 108.205 73.695 108.475 74.600 ;
        RECT 108.645 73.525 108.935 74.690 ;
        RECT 109.110 74.665 109.280 75.335 ;
        RECT 109.535 75.165 109.705 75.335 ;
        RECT 109.450 74.835 109.705 75.165 ;
        RECT 109.930 74.835 110.125 75.165 ;
        RECT 109.110 73.695 109.445 74.665 ;
        RECT 109.615 73.525 109.785 74.665 ;
        RECT 109.955 73.865 110.125 74.835 ;
        RECT 110.295 74.205 110.465 75.335 ;
        RECT 110.635 74.545 110.805 75.345 ;
        RECT 111.005 75.225 111.285 75.395 ;
        RECT 111.010 74.745 111.285 75.225 ;
        RECT 111.455 74.545 111.645 75.905 ;
        RECT 111.825 75.540 112.335 76.075 ;
        RECT 112.555 75.265 112.800 75.870 ;
        RECT 113.245 75.305 116.755 76.075 ;
        RECT 117.385 75.325 118.595 76.075 ;
        RECT 111.845 75.095 113.075 75.265 ;
        RECT 110.635 74.375 111.645 74.545 ;
        RECT 111.815 74.530 112.565 74.720 ;
        RECT 110.295 74.035 111.420 74.205 ;
        RECT 111.815 73.865 111.985 74.530 ;
        RECT 112.735 74.285 113.075 75.095 ;
        RECT 113.245 74.785 114.895 75.305 ;
        RECT 115.065 74.615 116.755 75.135 ;
        RECT 109.955 73.695 111.985 73.865 ;
        RECT 112.155 73.525 112.325 74.285 ;
        RECT 112.560 73.875 113.075 74.285 ;
        RECT 113.245 73.525 116.755 74.615 ;
        RECT 117.385 74.615 117.905 75.155 ;
        RECT 118.075 74.785 118.595 75.325 ;
        RECT 117.385 73.525 118.595 74.615 ;
        RECT 5.520 73.355 118.680 73.525 ;
        RECT 5.605 72.265 6.815 73.355 ;
        RECT 6.985 72.265 8.195 73.355 ;
        RECT 8.370 72.685 8.625 73.185 ;
        RECT 8.795 72.855 9.125 73.355 ;
        RECT 8.370 72.515 9.120 72.685 ;
        RECT 5.605 71.555 6.125 72.095 ;
        RECT 6.295 71.725 6.815 72.265 ;
        RECT 6.985 71.555 7.505 72.095 ;
        RECT 7.675 71.725 8.195 72.265 ;
        RECT 8.370 71.695 8.720 72.345 ;
        RECT 5.605 70.805 6.815 71.555 ;
        RECT 6.985 70.805 8.195 71.555 ;
        RECT 8.890 71.525 9.120 72.515 ;
        RECT 8.370 71.355 9.120 71.525 ;
        RECT 8.370 71.065 8.625 71.355 ;
        RECT 8.795 70.805 9.125 71.185 ;
        RECT 9.295 71.065 9.465 73.185 ;
        RECT 9.635 72.385 9.960 73.170 ;
        RECT 10.130 72.895 10.380 73.355 ;
        RECT 10.550 72.855 10.800 73.185 ;
        RECT 11.015 72.855 11.695 73.185 ;
        RECT 10.550 72.725 10.720 72.855 ;
        RECT 10.325 72.555 10.720 72.725 ;
        RECT 9.695 71.335 10.155 72.385 ;
        RECT 10.325 71.195 10.495 72.555 ;
        RECT 10.890 72.295 11.355 72.685 ;
        RECT 10.665 71.485 11.015 72.105 ;
        RECT 11.185 71.705 11.355 72.295 ;
        RECT 11.525 72.075 11.695 72.855 ;
        RECT 11.865 72.755 12.035 73.095 ;
        RECT 12.270 72.925 12.600 73.355 ;
        RECT 12.770 72.755 12.940 73.095 ;
        RECT 13.235 72.895 13.605 73.355 ;
        RECT 11.865 72.585 12.940 72.755 ;
        RECT 13.775 72.725 13.945 73.185 ;
        RECT 14.180 72.845 15.050 73.185 ;
        RECT 15.220 72.895 15.470 73.355 ;
        RECT 13.385 72.555 13.945 72.725 ;
        RECT 13.385 72.415 13.555 72.555 ;
        RECT 12.055 72.245 13.555 72.415 ;
        RECT 14.250 72.385 14.710 72.675 ;
        RECT 11.525 71.905 13.215 72.075 ;
        RECT 11.185 71.485 11.540 71.705 ;
        RECT 11.710 71.195 11.880 71.905 ;
        RECT 12.085 71.485 12.875 71.735 ;
        RECT 13.045 71.725 13.215 71.905 ;
        RECT 13.385 71.555 13.555 72.245 ;
        RECT 9.825 70.805 10.155 71.165 ;
        RECT 10.325 71.025 10.820 71.195 ;
        RECT 11.025 71.025 11.880 71.195 ;
        RECT 12.755 70.805 13.085 71.265 ;
        RECT 13.295 71.165 13.555 71.555 ;
        RECT 13.745 72.375 14.710 72.385 ;
        RECT 14.880 72.465 15.050 72.845 ;
        RECT 15.640 72.805 15.810 73.095 ;
        RECT 15.990 72.975 16.320 73.355 ;
        RECT 15.640 72.635 16.440 72.805 ;
        RECT 13.745 72.215 14.420 72.375 ;
        RECT 14.880 72.295 16.100 72.465 ;
        RECT 13.745 71.425 13.955 72.215 ;
        RECT 14.880 72.205 15.050 72.295 ;
        RECT 14.125 71.425 14.475 72.045 ;
        RECT 14.645 72.035 15.050 72.205 ;
        RECT 14.645 71.255 14.815 72.035 ;
        RECT 14.985 71.585 15.205 71.865 ;
        RECT 15.385 71.755 15.925 72.125 ;
        RECT 16.270 72.045 16.440 72.635 ;
        RECT 16.660 72.215 16.965 73.355 ;
        RECT 17.135 72.165 17.390 73.045 ;
        RECT 18.485 72.190 18.775 73.355 ;
        RECT 18.945 72.215 19.330 73.185 ;
        RECT 19.500 72.895 19.825 73.355 ;
        RECT 20.345 72.725 20.625 73.185 ;
        RECT 19.500 72.505 20.625 72.725 ;
        RECT 16.270 72.015 17.010 72.045 ;
        RECT 14.985 71.415 15.515 71.585 ;
        RECT 13.295 70.995 13.645 71.165 ;
        RECT 13.865 70.975 14.815 71.255 ;
        RECT 14.985 70.805 15.175 71.245 ;
        RECT 15.345 71.185 15.515 71.415 ;
        RECT 15.685 71.355 15.925 71.755 ;
        RECT 16.095 71.715 17.010 72.015 ;
        RECT 16.095 71.540 16.420 71.715 ;
        RECT 16.095 71.185 16.415 71.540 ;
        RECT 17.180 71.515 17.390 72.165 ;
        RECT 18.945 71.545 19.225 72.215 ;
        RECT 19.500 72.045 19.950 72.505 ;
        RECT 20.815 72.335 21.215 73.185 ;
        RECT 21.615 72.895 21.885 73.355 ;
        RECT 22.055 72.725 22.340 73.185 ;
        RECT 19.395 71.715 19.950 72.045 ;
        RECT 20.120 71.775 21.215 72.335 ;
        RECT 19.500 71.605 19.950 71.715 ;
        RECT 15.345 71.015 16.415 71.185 ;
        RECT 16.660 70.805 16.965 71.265 ;
        RECT 17.135 70.985 17.390 71.515 ;
        RECT 18.485 70.805 18.775 71.530 ;
        RECT 18.945 70.975 19.330 71.545 ;
        RECT 19.500 71.435 20.625 71.605 ;
        RECT 19.500 70.805 19.825 71.265 ;
        RECT 20.345 70.975 20.625 71.435 ;
        RECT 20.815 70.975 21.215 71.775 ;
        RECT 21.385 72.505 22.340 72.725 ;
        RECT 21.385 71.605 21.595 72.505 ;
        RECT 22.830 72.385 23.160 73.185 ;
        RECT 23.330 72.555 23.660 73.355 ;
        RECT 23.960 72.385 24.290 73.185 ;
        RECT 24.935 72.555 25.185 73.355 ;
        RECT 21.765 71.775 22.455 72.335 ;
        RECT 22.830 72.215 25.265 72.385 ;
        RECT 25.455 72.215 25.625 73.355 ;
        RECT 25.795 72.215 26.135 73.185 ;
        RECT 26.305 72.265 27.515 73.355 ;
        RECT 27.690 72.685 27.945 73.185 ;
        RECT 28.115 72.855 28.445 73.355 ;
        RECT 27.690 72.515 28.440 72.685 ;
        RECT 22.625 71.795 22.975 72.045 ;
        RECT 21.385 71.435 22.340 71.605 ;
        RECT 23.160 71.585 23.330 72.215 ;
        RECT 23.500 71.795 23.830 71.995 ;
        RECT 24.000 71.795 24.330 71.995 ;
        RECT 24.500 71.795 24.920 71.995 ;
        RECT 25.095 71.965 25.265 72.215 ;
        RECT 25.095 71.795 25.790 71.965 ;
        RECT 21.615 70.805 21.885 71.265 ;
        RECT 22.055 70.975 22.340 71.435 ;
        RECT 22.830 70.975 23.330 71.585 ;
        RECT 23.960 71.455 25.185 71.625 ;
        RECT 25.960 71.605 26.135 72.215 ;
        RECT 23.960 70.975 24.290 71.455 ;
        RECT 24.460 70.805 24.685 71.265 ;
        RECT 24.855 70.975 25.185 71.455 ;
        RECT 25.375 70.805 25.625 71.605 ;
        RECT 25.795 70.975 26.135 71.605 ;
        RECT 26.305 71.555 26.825 72.095 ;
        RECT 26.995 71.725 27.515 72.265 ;
        RECT 27.690 71.695 28.040 72.345 ;
        RECT 26.305 70.805 27.515 71.555 ;
        RECT 28.210 71.525 28.440 72.515 ;
        RECT 27.690 71.355 28.440 71.525 ;
        RECT 27.690 71.065 27.945 71.355 ;
        RECT 28.115 70.805 28.445 71.185 ;
        RECT 28.615 71.065 28.785 73.185 ;
        RECT 28.955 72.385 29.280 73.170 ;
        RECT 29.450 72.895 29.700 73.355 ;
        RECT 29.870 72.855 30.120 73.185 ;
        RECT 30.335 72.855 31.015 73.185 ;
        RECT 29.870 72.725 30.040 72.855 ;
        RECT 29.645 72.555 30.040 72.725 ;
        RECT 29.015 71.335 29.475 72.385 ;
        RECT 29.645 71.195 29.815 72.555 ;
        RECT 30.210 72.295 30.675 72.685 ;
        RECT 29.985 71.485 30.335 72.105 ;
        RECT 30.505 71.705 30.675 72.295 ;
        RECT 30.845 72.075 31.015 72.855 ;
        RECT 31.185 72.755 31.355 73.095 ;
        RECT 31.590 72.925 31.920 73.355 ;
        RECT 32.090 72.755 32.260 73.095 ;
        RECT 32.555 72.895 32.925 73.355 ;
        RECT 31.185 72.585 32.260 72.755 ;
        RECT 33.095 72.725 33.265 73.185 ;
        RECT 33.500 72.845 34.370 73.185 ;
        RECT 34.540 72.895 34.790 73.355 ;
        RECT 32.705 72.555 33.265 72.725 ;
        RECT 32.705 72.415 32.875 72.555 ;
        RECT 31.375 72.245 32.875 72.415 ;
        RECT 33.570 72.385 34.030 72.675 ;
        RECT 30.845 71.905 32.535 72.075 ;
        RECT 30.505 71.485 30.860 71.705 ;
        RECT 31.030 71.195 31.200 71.905 ;
        RECT 31.405 71.485 32.195 71.735 ;
        RECT 32.365 71.725 32.535 71.905 ;
        RECT 32.705 71.555 32.875 72.245 ;
        RECT 29.145 70.805 29.475 71.165 ;
        RECT 29.645 71.025 30.140 71.195 ;
        RECT 30.345 71.025 31.200 71.195 ;
        RECT 32.075 70.805 32.405 71.265 ;
        RECT 32.615 71.165 32.875 71.555 ;
        RECT 33.065 72.375 34.030 72.385 ;
        RECT 34.200 72.465 34.370 72.845 ;
        RECT 34.960 72.805 35.130 73.095 ;
        RECT 35.310 72.975 35.640 73.355 ;
        RECT 34.960 72.635 35.760 72.805 ;
        RECT 33.065 72.215 33.740 72.375 ;
        RECT 34.200 72.295 35.420 72.465 ;
        RECT 33.065 71.425 33.275 72.215 ;
        RECT 34.200 72.205 34.370 72.295 ;
        RECT 33.445 71.425 33.795 72.045 ;
        RECT 33.965 72.035 34.370 72.205 ;
        RECT 33.965 71.255 34.135 72.035 ;
        RECT 34.305 71.585 34.525 71.865 ;
        RECT 34.705 71.755 35.245 72.125 ;
        RECT 35.590 72.045 35.760 72.635 ;
        RECT 35.980 72.215 36.285 73.355 ;
        RECT 36.455 72.165 36.710 73.045 ;
        RECT 36.885 72.265 38.555 73.355 ;
        RECT 35.590 72.015 36.330 72.045 ;
        RECT 34.305 71.415 34.835 71.585 ;
        RECT 32.615 70.995 32.965 71.165 ;
        RECT 33.185 70.975 34.135 71.255 ;
        RECT 34.305 70.805 34.495 71.245 ;
        RECT 34.665 71.185 34.835 71.415 ;
        RECT 35.005 71.355 35.245 71.755 ;
        RECT 35.415 71.715 36.330 72.015 ;
        RECT 35.415 71.540 35.740 71.715 ;
        RECT 35.415 71.185 35.735 71.540 ;
        RECT 36.500 71.515 36.710 72.165 ;
        RECT 34.665 71.015 35.735 71.185 ;
        RECT 35.980 70.805 36.285 71.265 ;
        RECT 36.455 70.985 36.710 71.515 ;
        RECT 36.885 71.575 37.635 72.095 ;
        RECT 37.805 71.745 38.555 72.265 ;
        RECT 38.765 72.215 38.995 73.355 ;
        RECT 39.165 72.205 39.495 73.185 ;
        RECT 39.665 72.215 39.875 73.355 ;
        RECT 40.105 72.280 40.375 73.185 ;
        RECT 40.545 72.595 40.875 73.355 ;
        RECT 41.055 72.425 41.225 73.185 ;
        RECT 38.745 71.795 39.075 72.045 ;
        RECT 36.885 70.805 38.555 71.575 ;
        RECT 38.765 70.805 38.995 71.625 ;
        RECT 39.245 71.605 39.495 72.205 ;
        RECT 39.165 70.975 39.495 71.605 ;
        RECT 39.665 70.805 39.875 71.625 ;
        RECT 40.105 71.480 40.275 72.280 ;
        RECT 40.560 72.255 41.225 72.425 ;
        RECT 40.560 72.110 40.730 72.255 ;
        RECT 42.445 72.215 42.675 73.355 ;
        RECT 42.845 72.205 43.175 73.185 ;
        RECT 43.345 72.215 43.555 73.355 ;
        RECT 40.445 71.780 40.730 72.110 ;
        RECT 40.560 71.525 40.730 71.780 ;
        RECT 40.965 71.705 41.295 72.075 ;
        RECT 42.425 71.795 42.755 72.045 ;
        RECT 40.105 70.975 40.365 71.480 ;
        RECT 40.560 71.355 41.225 71.525 ;
        RECT 40.545 70.805 40.875 71.185 ;
        RECT 41.055 70.975 41.225 71.355 ;
        RECT 42.445 70.805 42.675 71.625 ;
        RECT 42.925 71.605 43.175 72.205 ;
        RECT 44.245 72.190 44.535 73.355 ;
        RECT 44.710 72.215 45.045 73.185 ;
        RECT 45.215 72.215 45.385 73.355 ;
        RECT 45.555 73.015 47.585 73.185 ;
        RECT 42.845 70.975 43.175 71.605 ;
        RECT 43.345 70.805 43.555 71.625 ;
        RECT 44.710 71.545 44.880 72.215 ;
        RECT 45.555 72.045 45.725 73.015 ;
        RECT 45.050 71.715 45.305 72.045 ;
        RECT 45.530 71.715 45.725 72.045 ;
        RECT 45.895 72.675 47.020 72.845 ;
        RECT 45.135 71.545 45.305 71.715 ;
        RECT 45.895 71.545 46.065 72.675 ;
        RECT 44.245 70.805 44.535 71.530 ;
        RECT 44.710 70.975 44.965 71.545 ;
        RECT 45.135 71.375 46.065 71.545 ;
        RECT 46.235 72.335 47.245 72.505 ;
        RECT 46.235 71.535 46.405 72.335 ;
        RECT 46.610 71.995 46.885 72.135 ;
        RECT 46.605 71.825 46.885 71.995 ;
        RECT 45.890 71.340 46.065 71.375 ;
        RECT 45.135 70.805 45.465 71.205 ;
        RECT 45.890 70.975 46.420 71.340 ;
        RECT 46.610 70.975 46.885 71.825 ;
        RECT 47.055 70.975 47.245 72.335 ;
        RECT 47.415 72.350 47.585 73.015 ;
        RECT 47.755 72.595 47.925 73.355 ;
        RECT 48.160 72.595 48.675 73.005 ;
        RECT 47.415 72.160 48.165 72.350 ;
        RECT 48.335 71.785 48.675 72.595 ;
        RECT 48.845 72.265 52.355 73.355 ;
        RECT 52.990 72.845 54.645 73.135 ;
        RECT 47.445 71.615 48.675 71.785 ;
        RECT 47.425 70.805 47.935 71.340 ;
        RECT 48.155 71.010 48.400 71.615 ;
        RECT 48.845 71.575 50.495 72.095 ;
        RECT 50.665 71.745 52.355 72.265 ;
        RECT 52.990 72.505 54.580 72.675 ;
        RECT 54.815 72.555 55.095 73.355 ;
        RECT 52.990 72.215 53.310 72.505 ;
        RECT 54.410 72.385 54.580 72.505 ;
        RECT 53.505 72.165 54.220 72.335 ;
        RECT 54.410 72.215 55.135 72.385 ;
        RECT 55.305 72.215 55.575 73.185 ;
        RECT 55.800 72.485 56.085 73.355 ;
        RECT 56.255 72.725 56.515 73.185 ;
        RECT 56.690 72.895 56.945 73.355 ;
        RECT 57.115 72.725 57.375 73.185 ;
        RECT 56.255 72.555 57.375 72.725 ;
        RECT 57.545 72.555 57.855 73.355 ;
        RECT 56.255 72.305 56.515 72.555 ;
        RECT 58.025 72.385 58.335 73.185 ;
        RECT 48.845 70.805 52.355 71.575 ;
        RECT 52.990 71.475 53.340 72.045 ;
        RECT 53.510 71.715 54.220 72.165 ;
        RECT 54.965 72.045 55.135 72.215 ;
        RECT 54.390 71.715 54.795 72.045 ;
        RECT 54.965 71.715 55.235 72.045 ;
        RECT 54.965 71.545 55.135 71.715 ;
        RECT 53.525 71.375 55.135 71.545 ;
        RECT 55.405 71.480 55.575 72.215 ;
        RECT 52.995 70.805 53.325 71.305 ;
        RECT 53.525 71.025 53.695 71.375 ;
        RECT 53.895 70.805 54.225 71.205 ;
        RECT 54.395 71.025 54.565 71.375 ;
        RECT 54.735 70.805 55.115 71.205 ;
        RECT 55.305 71.135 55.575 71.480 ;
        RECT 55.760 72.135 56.515 72.305 ;
        RECT 57.305 72.215 58.335 72.385 ;
        RECT 55.760 71.625 56.165 72.135 ;
        RECT 57.305 71.965 57.475 72.215 ;
        RECT 56.335 71.795 57.475 71.965 ;
        RECT 55.760 71.455 57.410 71.625 ;
        RECT 57.645 71.475 57.995 72.045 ;
        RECT 55.805 70.805 56.085 71.285 ;
        RECT 56.255 71.065 56.515 71.455 ;
        RECT 56.690 70.805 56.945 71.285 ;
        RECT 57.115 71.065 57.410 71.455 ;
        RECT 58.165 71.305 58.335 72.215 ;
        RECT 57.590 70.805 57.865 71.285 ;
        RECT 58.035 70.975 58.335 71.305 ;
        RECT 59.425 72.385 59.735 73.185 ;
        RECT 59.905 72.555 60.215 73.355 ;
        RECT 60.385 72.725 60.645 73.185 ;
        RECT 60.815 72.895 61.070 73.355 ;
        RECT 61.245 72.725 61.505 73.185 ;
        RECT 60.385 72.555 61.505 72.725 ;
        RECT 59.425 72.215 60.455 72.385 ;
        RECT 59.425 71.305 59.595 72.215 ;
        RECT 59.765 71.475 60.115 72.045 ;
        RECT 60.285 71.965 60.455 72.215 ;
        RECT 61.245 72.305 61.505 72.555 ;
        RECT 61.675 72.485 61.960 73.355 ;
        RECT 62.275 72.425 62.445 73.185 ;
        RECT 62.660 72.595 62.990 73.355 ;
        RECT 61.245 72.135 62.000 72.305 ;
        RECT 62.275 72.255 62.990 72.425 ;
        RECT 63.160 72.280 63.415 73.185 ;
        RECT 60.285 71.795 61.425 71.965 ;
        RECT 61.595 71.625 62.000 72.135 ;
        RECT 62.185 71.705 62.540 72.075 ;
        RECT 62.820 72.045 62.990 72.255 ;
        RECT 62.820 71.715 63.075 72.045 ;
        RECT 60.350 71.455 62.000 71.625 ;
        RECT 62.820 71.525 62.990 71.715 ;
        RECT 63.245 71.550 63.415 72.280 ;
        RECT 63.590 72.205 63.850 73.355 ;
        RECT 64.030 72.205 64.290 73.355 ;
        RECT 64.465 72.280 64.720 73.185 ;
        RECT 64.890 72.595 65.220 73.355 ;
        RECT 65.435 72.425 65.605 73.185 ;
        RECT 59.425 70.975 59.725 71.305 ;
        RECT 59.895 70.805 60.170 71.285 ;
        RECT 60.350 71.065 60.645 71.455 ;
        RECT 60.815 70.805 61.070 71.285 ;
        RECT 61.245 71.065 61.505 71.455 ;
        RECT 62.275 71.355 62.990 71.525 ;
        RECT 61.675 70.805 61.955 71.285 ;
        RECT 62.275 70.975 62.445 71.355 ;
        RECT 62.660 70.805 62.990 71.185 ;
        RECT 63.160 70.975 63.415 71.550 ;
        RECT 63.590 70.805 63.850 71.645 ;
        RECT 64.030 70.805 64.290 71.645 ;
        RECT 64.465 71.550 64.635 72.280 ;
        RECT 64.890 72.255 65.605 72.425 ;
        RECT 65.865 72.265 67.535 73.355 ;
        RECT 64.890 72.045 65.060 72.255 ;
        RECT 64.805 71.715 65.060 72.045 ;
        RECT 64.465 70.975 64.720 71.550 ;
        RECT 64.890 71.525 65.060 71.715 ;
        RECT 65.340 71.705 65.695 72.075 ;
        RECT 65.865 71.575 66.615 72.095 ;
        RECT 66.785 71.745 67.535 72.265 ;
        RECT 68.165 72.280 68.435 73.185 ;
        RECT 68.605 72.595 68.935 73.355 ;
        RECT 69.115 72.425 69.285 73.185 ;
        RECT 64.890 71.355 65.605 71.525 ;
        RECT 64.890 70.805 65.220 71.185 ;
        RECT 65.435 70.975 65.605 71.355 ;
        RECT 65.865 70.805 67.535 71.575 ;
        RECT 68.165 71.480 68.335 72.280 ;
        RECT 68.620 72.255 69.285 72.425 ;
        RECT 68.620 72.110 68.790 72.255 ;
        RECT 70.005 72.190 70.295 73.355 ;
        RECT 70.555 72.425 70.725 73.185 ;
        RECT 70.905 72.595 71.235 73.355 ;
        RECT 70.555 72.255 71.220 72.425 ;
        RECT 71.405 72.280 71.675 73.185 ;
        RECT 68.505 71.780 68.790 72.110 ;
        RECT 71.050 72.110 71.220 72.255 ;
        RECT 68.620 71.525 68.790 71.780 ;
        RECT 69.025 71.705 69.355 72.075 ;
        RECT 70.485 71.705 70.815 72.075 ;
        RECT 71.050 71.780 71.335 72.110 ;
        RECT 68.165 70.975 68.425 71.480 ;
        RECT 68.620 71.355 69.285 71.525 ;
        RECT 68.605 70.805 68.935 71.185 ;
        RECT 69.115 70.975 69.285 71.355 ;
        RECT 70.005 70.805 70.295 71.530 ;
        RECT 71.050 71.525 71.220 71.780 ;
        RECT 70.555 71.355 71.220 71.525 ;
        RECT 71.505 71.480 71.675 72.280 ;
        RECT 70.555 70.975 70.725 71.355 ;
        RECT 70.905 70.805 71.235 71.185 ;
        RECT 71.415 70.975 71.675 71.480 ;
        RECT 72.310 72.215 72.645 73.185 ;
        RECT 72.815 72.215 72.985 73.355 ;
        RECT 73.155 73.015 75.185 73.185 ;
        RECT 72.310 71.545 72.480 72.215 ;
        RECT 73.155 72.045 73.325 73.015 ;
        RECT 72.650 71.715 72.905 72.045 ;
        RECT 73.130 71.715 73.325 72.045 ;
        RECT 73.495 72.675 74.620 72.845 ;
        RECT 72.735 71.545 72.905 71.715 ;
        RECT 73.495 71.545 73.665 72.675 ;
        RECT 72.310 70.975 72.565 71.545 ;
        RECT 72.735 71.375 73.665 71.545 ;
        RECT 73.835 72.335 74.845 72.505 ;
        RECT 73.835 71.535 74.005 72.335 ;
        RECT 74.210 71.995 74.485 72.135 ;
        RECT 74.205 71.825 74.485 71.995 ;
        RECT 73.490 71.340 73.665 71.375 ;
        RECT 72.735 70.805 73.065 71.205 ;
        RECT 73.490 70.975 74.020 71.340 ;
        RECT 74.210 70.975 74.485 71.825 ;
        RECT 74.655 70.975 74.845 72.335 ;
        RECT 75.015 72.350 75.185 73.015 ;
        RECT 75.355 72.595 75.525 73.355 ;
        RECT 75.760 72.595 76.275 73.005 ;
        RECT 75.015 72.160 75.765 72.350 ;
        RECT 75.935 71.785 76.275 72.595 ;
        RECT 76.445 72.265 78.115 73.355 ;
        RECT 75.045 71.615 76.275 71.785 ;
        RECT 75.025 70.805 75.535 71.340 ;
        RECT 75.755 71.010 76.000 71.615 ;
        RECT 76.445 71.575 77.195 72.095 ;
        RECT 77.365 71.745 78.115 72.265 ;
        RECT 78.490 72.385 78.820 73.185 ;
        RECT 78.990 72.555 79.320 73.355 ;
        RECT 79.620 72.385 79.950 73.185 ;
        RECT 80.595 72.555 80.845 73.355 ;
        RECT 78.490 72.215 80.925 72.385 ;
        RECT 81.115 72.215 81.285 73.355 ;
        RECT 81.455 72.215 81.795 73.185 ;
        RECT 78.285 71.795 78.635 72.045 ;
        RECT 78.820 71.585 78.990 72.215 ;
        RECT 79.160 71.795 79.490 71.995 ;
        RECT 79.660 71.795 79.990 71.995 ;
        RECT 80.160 71.795 80.580 71.995 ;
        RECT 80.755 71.965 80.925 72.215 ;
        RECT 80.755 71.795 81.450 71.965 ;
        RECT 76.445 70.805 78.115 71.575 ;
        RECT 78.490 70.975 78.990 71.585 ;
        RECT 79.620 71.455 80.845 71.625 ;
        RECT 81.620 71.605 81.795 72.215 ;
        RECT 79.620 70.975 79.950 71.455 ;
        RECT 80.120 70.805 80.345 71.265 ;
        RECT 80.515 70.975 80.845 71.455 ;
        RECT 81.035 70.805 81.285 71.605 ;
        RECT 81.455 70.975 81.795 71.605 ;
        RECT 81.965 72.215 82.235 73.185 ;
        RECT 82.445 72.555 82.725 73.355 ;
        RECT 82.895 72.845 84.550 73.135 ;
        RECT 82.960 72.505 84.550 72.675 ;
        RECT 82.960 72.385 83.130 72.505 ;
        RECT 82.405 72.215 83.130 72.385 ;
        RECT 81.965 71.480 82.135 72.215 ;
        RECT 82.405 72.045 82.575 72.215 ;
        RECT 82.305 71.715 82.575 72.045 ;
        RECT 82.745 71.715 83.150 72.045 ;
        RECT 83.320 71.715 84.030 72.335 ;
        RECT 84.230 72.215 84.550 72.505 ;
        RECT 84.725 72.265 88.235 73.355 ;
        RECT 82.405 71.545 82.575 71.715 ;
        RECT 81.965 71.135 82.235 71.480 ;
        RECT 82.405 71.375 84.015 71.545 ;
        RECT 84.200 71.475 84.550 72.045 ;
        RECT 84.725 71.575 86.375 72.095 ;
        RECT 86.545 71.745 88.235 72.265 ;
        RECT 88.610 72.385 88.940 73.185 ;
        RECT 89.110 72.555 89.440 73.355 ;
        RECT 89.740 72.385 90.070 73.185 ;
        RECT 90.715 72.555 90.965 73.355 ;
        RECT 88.610 72.215 91.045 72.385 ;
        RECT 91.235 72.215 91.405 73.355 ;
        RECT 91.575 72.215 91.915 73.185 ;
        RECT 92.085 72.265 95.595 73.355 ;
        RECT 88.405 71.795 88.755 72.045 ;
        RECT 88.940 71.585 89.110 72.215 ;
        RECT 89.280 71.795 89.610 71.995 ;
        RECT 89.780 71.795 90.110 71.995 ;
        RECT 90.280 71.795 90.700 71.995 ;
        RECT 90.875 71.965 91.045 72.215 ;
        RECT 90.875 71.795 91.570 71.965 ;
        RECT 82.425 70.805 82.805 71.205 ;
        RECT 82.975 71.025 83.145 71.375 ;
        RECT 83.315 70.805 83.645 71.205 ;
        RECT 83.845 71.025 84.015 71.375 ;
        RECT 84.215 70.805 84.545 71.305 ;
        RECT 84.725 70.805 88.235 71.575 ;
        RECT 88.610 70.975 89.110 71.585 ;
        RECT 89.740 71.455 90.965 71.625 ;
        RECT 91.740 71.605 91.915 72.215 ;
        RECT 89.740 70.975 90.070 71.455 ;
        RECT 90.240 70.805 90.465 71.265 ;
        RECT 90.635 70.975 90.965 71.455 ;
        RECT 91.155 70.805 91.405 71.605 ;
        RECT 91.575 70.975 91.915 71.605 ;
        RECT 92.085 71.575 93.735 72.095 ;
        RECT 93.905 71.745 95.595 72.265 ;
        RECT 95.765 72.190 96.055 73.355 ;
        RECT 96.225 72.280 96.495 73.185 ;
        RECT 96.665 72.595 96.995 73.355 ;
        RECT 97.175 72.425 97.345 73.185 ;
        RECT 92.085 70.805 95.595 71.575 ;
        RECT 95.765 70.805 96.055 71.530 ;
        RECT 96.225 71.480 96.395 72.280 ;
        RECT 96.680 72.255 97.345 72.425 ;
        RECT 97.605 72.265 98.815 73.355 ;
        RECT 96.680 72.110 96.850 72.255 ;
        RECT 96.565 71.780 96.850 72.110 ;
        RECT 96.680 71.525 96.850 71.780 ;
        RECT 97.085 71.705 97.415 72.075 ;
        RECT 97.605 71.555 98.125 72.095 ;
        RECT 98.295 71.725 98.815 72.265 ;
        RECT 99.045 72.215 99.255 73.355 ;
        RECT 99.425 72.205 99.755 73.185 ;
        RECT 99.925 72.215 100.155 73.355 ;
        RECT 100.365 72.920 105.710 73.355 ;
        RECT 96.225 70.975 96.485 71.480 ;
        RECT 96.680 71.355 97.345 71.525 ;
        RECT 96.665 70.805 96.995 71.185 ;
        RECT 97.175 70.975 97.345 71.355 ;
        RECT 97.605 70.805 98.815 71.555 ;
        RECT 99.045 70.805 99.255 71.625 ;
        RECT 99.425 71.605 99.675 72.205 ;
        RECT 99.845 71.795 100.175 72.045 ;
        RECT 99.425 70.975 99.755 71.605 ;
        RECT 99.925 70.805 100.155 71.625 ;
        RECT 101.950 71.350 102.290 72.180 ;
        RECT 103.770 71.670 104.120 72.920 ;
        RECT 105.885 72.265 107.095 73.355 ;
        RECT 107.355 72.685 107.525 73.185 ;
        RECT 107.695 72.855 108.025 73.355 ;
        RECT 107.355 72.515 108.020 72.685 ;
        RECT 105.885 71.555 106.405 72.095 ;
        RECT 106.575 71.725 107.095 72.265 ;
        RECT 107.270 71.695 107.620 72.345 ;
        RECT 100.365 70.805 105.710 71.350 ;
        RECT 105.885 70.805 107.095 71.555 ;
        RECT 107.790 71.525 108.020 72.515 ;
        RECT 107.355 71.355 108.020 71.525 ;
        RECT 107.355 71.065 107.525 71.355 ;
        RECT 107.695 70.805 108.025 71.185 ;
        RECT 108.195 71.065 108.420 73.185 ;
        RECT 108.635 72.855 108.965 73.355 ;
        RECT 109.135 72.685 109.305 73.185 ;
        RECT 109.540 72.970 110.370 73.140 ;
        RECT 110.610 72.975 110.990 73.355 ;
        RECT 108.610 72.515 109.305 72.685 ;
        RECT 108.610 71.545 108.780 72.515 ;
        RECT 108.950 71.725 109.360 72.345 ;
        RECT 109.530 72.295 110.030 72.675 ;
        RECT 108.610 71.355 109.305 71.545 ;
        RECT 109.530 71.425 109.750 72.295 ;
        RECT 110.200 72.125 110.370 72.970 ;
        RECT 111.170 72.805 111.340 73.095 ;
        RECT 111.510 72.975 111.840 73.355 ;
        RECT 112.310 72.885 112.940 73.135 ;
        RECT 113.120 72.975 113.540 73.355 ;
        RECT 112.770 72.805 112.940 72.885 ;
        RECT 113.740 72.805 113.980 73.095 ;
        RECT 110.540 72.555 111.910 72.805 ;
        RECT 110.540 72.295 110.790 72.555 ;
        RECT 111.300 72.125 111.550 72.285 ;
        RECT 110.200 71.955 111.550 72.125 ;
        RECT 110.200 71.915 110.620 71.955 ;
        RECT 109.930 71.365 110.280 71.735 ;
        RECT 108.635 70.805 108.965 71.185 ;
        RECT 109.135 71.025 109.305 71.355 ;
        RECT 110.450 71.185 110.620 71.915 ;
        RECT 111.720 71.785 111.910 72.555 ;
        RECT 110.790 71.455 111.200 71.785 ;
        RECT 111.490 71.445 111.910 71.785 ;
        RECT 112.080 72.375 112.600 72.685 ;
        RECT 112.770 72.635 113.980 72.805 ;
        RECT 114.210 72.665 114.540 73.355 ;
        RECT 112.080 71.615 112.250 72.375 ;
        RECT 112.420 71.785 112.600 72.195 ;
        RECT 112.770 72.125 112.940 72.635 ;
        RECT 114.710 72.485 114.880 73.095 ;
        RECT 115.150 72.635 115.480 73.145 ;
        RECT 114.710 72.465 115.030 72.485 ;
        RECT 113.110 72.295 115.030 72.465 ;
        RECT 112.770 71.955 114.670 72.125 ;
        RECT 113.000 71.615 113.330 71.735 ;
        RECT 112.080 71.445 113.330 71.615 ;
        RECT 109.605 70.985 110.620 71.185 ;
        RECT 110.790 70.805 111.200 71.245 ;
        RECT 111.490 71.015 111.740 71.445 ;
        RECT 111.940 70.805 112.260 71.265 ;
        RECT 113.500 71.195 113.670 71.955 ;
        RECT 114.340 71.895 114.670 71.955 ;
        RECT 113.860 71.725 114.190 71.785 ;
        RECT 113.860 71.455 114.520 71.725 ;
        RECT 114.840 71.400 115.030 72.295 ;
        RECT 112.820 71.025 113.670 71.195 ;
        RECT 113.870 70.805 114.530 71.285 ;
        RECT 114.710 71.070 115.030 71.400 ;
        RECT 115.230 72.045 115.480 72.635 ;
        RECT 115.660 72.555 115.945 73.355 ;
        RECT 116.125 72.375 116.380 73.045 ;
        RECT 116.200 72.335 116.380 72.375 ;
        RECT 116.200 72.165 116.465 72.335 ;
        RECT 117.385 72.265 118.595 73.355 ;
        RECT 115.230 71.715 116.030 72.045 ;
        RECT 115.230 71.065 115.480 71.715 ;
        RECT 116.200 71.515 116.380 72.165 ;
        RECT 117.385 71.725 117.905 72.265 ;
        RECT 118.075 71.555 118.595 72.095 ;
        RECT 115.660 70.805 115.945 71.265 ;
        RECT 116.125 70.985 116.380 71.515 ;
        RECT 117.385 70.805 118.595 71.555 ;
        RECT 5.520 70.635 118.680 70.805 ;
        RECT 5.605 69.885 6.815 70.635 ;
        RECT 5.605 69.345 6.125 69.885 ;
        RECT 6.985 69.865 10.495 70.635 ;
        RECT 11.585 69.960 11.845 70.465 ;
        RECT 12.025 70.255 12.355 70.635 ;
        RECT 12.535 70.085 12.705 70.465 ;
        RECT 6.295 69.175 6.815 69.715 ;
        RECT 6.985 69.345 8.635 69.865 ;
        RECT 8.805 69.175 10.495 69.695 ;
        RECT 5.605 68.085 6.815 69.175 ;
        RECT 6.985 68.085 10.495 69.175 ;
        RECT 11.585 69.160 11.755 69.960 ;
        RECT 12.040 69.915 12.705 70.085 ;
        RECT 12.040 69.660 12.210 69.915 ;
        RECT 13.465 69.815 13.695 70.635 ;
        RECT 13.865 69.835 14.195 70.465 ;
        RECT 11.925 69.330 12.210 69.660 ;
        RECT 12.445 69.365 12.775 69.735 ;
        RECT 13.445 69.395 13.775 69.645 ;
        RECT 12.040 69.185 12.210 69.330 ;
        RECT 13.945 69.235 14.195 69.835 ;
        RECT 14.365 69.815 14.575 70.635 ;
        RECT 14.805 70.090 20.150 70.635 ;
        RECT 16.390 69.260 16.730 70.090 ;
        RECT 20.990 69.855 21.490 70.465 ;
        RECT 11.585 68.255 11.855 69.160 ;
        RECT 12.040 69.015 12.705 69.185 ;
        RECT 12.025 68.085 12.355 68.845 ;
        RECT 12.535 68.255 12.705 69.015 ;
        RECT 13.465 68.085 13.695 69.225 ;
        RECT 13.865 68.255 14.195 69.235 ;
        RECT 14.365 68.085 14.575 69.225 ;
        RECT 18.210 68.520 18.560 69.770 ;
        RECT 20.785 69.395 21.135 69.645 ;
        RECT 21.320 69.225 21.490 69.855 ;
        RECT 22.120 69.985 22.450 70.465 ;
        RECT 22.620 70.175 22.845 70.635 ;
        RECT 23.015 69.985 23.345 70.465 ;
        RECT 22.120 69.815 23.345 69.985 ;
        RECT 23.535 69.835 23.785 70.635 ;
        RECT 23.955 69.835 24.295 70.465 ;
        RECT 24.670 69.855 25.170 70.465 ;
        RECT 24.065 69.785 24.295 69.835 ;
        RECT 21.660 69.445 21.990 69.645 ;
        RECT 22.160 69.445 22.490 69.645 ;
        RECT 22.660 69.445 23.080 69.645 ;
        RECT 23.255 69.475 23.950 69.645 ;
        RECT 23.255 69.225 23.425 69.475 ;
        RECT 24.120 69.225 24.295 69.785 ;
        RECT 24.465 69.395 24.815 69.645 ;
        RECT 25.000 69.225 25.170 69.855 ;
        RECT 25.800 69.985 26.130 70.465 ;
        RECT 26.300 70.175 26.525 70.635 ;
        RECT 26.695 69.985 27.025 70.465 ;
        RECT 25.800 69.815 27.025 69.985 ;
        RECT 27.215 69.835 27.465 70.635 ;
        RECT 27.635 69.835 27.975 70.465 ;
        RECT 28.155 70.135 28.485 70.635 ;
        RECT 28.685 70.065 28.855 70.415 ;
        RECT 29.055 70.235 29.385 70.635 ;
        RECT 29.555 70.065 29.725 70.415 ;
        RECT 29.895 70.235 30.275 70.635 ;
        RECT 25.340 69.445 25.670 69.645 ;
        RECT 25.840 69.445 26.170 69.645 ;
        RECT 26.340 69.445 26.760 69.645 ;
        RECT 26.935 69.475 27.630 69.645 ;
        RECT 26.935 69.225 27.105 69.475 ;
        RECT 27.800 69.225 27.975 69.835 ;
        RECT 28.150 69.395 28.500 69.965 ;
        RECT 28.685 69.895 30.295 70.065 ;
        RECT 30.465 69.960 30.735 70.305 ;
        RECT 30.125 69.725 30.295 69.895 ;
        RECT 28.670 69.275 29.380 69.725 ;
        RECT 29.550 69.395 29.955 69.725 ;
        RECT 30.125 69.395 30.395 69.725 ;
        RECT 20.990 69.055 23.425 69.225 ;
        RECT 14.805 68.085 20.150 68.520 ;
        RECT 20.990 68.255 21.320 69.055 ;
        RECT 21.490 68.085 21.820 68.885 ;
        RECT 22.120 68.255 22.450 69.055 ;
        RECT 23.095 68.085 23.345 68.885 ;
        RECT 23.615 68.085 23.785 69.225 ;
        RECT 23.955 68.255 24.295 69.225 ;
        RECT 24.670 69.055 27.105 69.225 ;
        RECT 24.670 68.255 25.000 69.055 ;
        RECT 25.170 68.085 25.500 68.885 ;
        RECT 25.800 68.255 26.130 69.055 ;
        RECT 26.775 68.085 27.025 68.885 ;
        RECT 27.295 68.085 27.465 69.225 ;
        RECT 27.635 68.255 27.975 69.225 ;
        RECT 28.150 68.935 28.470 69.225 ;
        RECT 28.665 69.105 29.380 69.275 ;
        RECT 30.125 69.225 30.295 69.395 ;
        RECT 30.565 69.225 30.735 69.960 ;
        RECT 31.365 69.910 31.655 70.635 ;
        RECT 31.825 70.090 37.170 70.635 ;
        RECT 33.410 69.260 33.750 70.090 ;
        RECT 37.435 70.085 37.605 70.375 ;
        RECT 37.775 70.255 38.105 70.635 ;
        RECT 37.435 69.915 38.100 70.085 ;
        RECT 29.570 69.055 30.295 69.225 ;
        RECT 29.570 68.935 29.740 69.055 ;
        RECT 28.150 68.765 29.740 68.935 ;
        RECT 28.150 68.305 29.805 68.595 ;
        RECT 29.975 68.085 30.255 68.885 ;
        RECT 30.465 68.255 30.735 69.225 ;
        RECT 31.365 68.085 31.655 69.250 ;
        RECT 35.230 68.520 35.580 69.770 ;
        RECT 37.350 69.095 37.700 69.745 ;
        RECT 37.870 68.925 38.100 69.915 ;
        RECT 37.435 68.755 38.100 68.925 ;
        RECT 31.825 68.085 37.170 68.520 ;
        RECT 37.435 68.255 37.605 68.755 ;
        RECT 37.775 68.085 38.105 68.585 ;
        RECT 38.275 68.255 38.500 70.375 ;
        RECT 38.715 70.255 39.045 70.635 ;
        RECT 39.215 70.085 39.385 70.415 ;
        RECT 39.685 70.255 40.700 70.455 ;
        RECT 38.690 69.895 39.385 70.085 ;
        RECT 38.690 68.925 38.860 69.895 ;
        RECT 39.030 69.095 39.440 69.715 ;
        RECT 39.610 69.145 39.830 70.015 ;
        RECT 40.010 69.705 40.360 70.075 ;
        RECT 40.530 69.525 40.700 70.255 ;
        RECT 40.870 70.195 41.280 70.635 ;
        RECT 41.570 69.995 41.820 70.425 ;
        RECT 42.020 70.175 42.340 70.635 ;
        RECT 42.900 70.245 43.750 70.415 ;
        RECT 40.870 69.655 41.280 69.985 ;
        RECT 41.570 69.655 41.990 69.995 ;
        RECT 40.280 69.485 40.700 69.525 ;
        RECT 40.280 69.315 41.630 69.485 ;
        RECT 38.690 68.755 39.385 68.925 ;
        RECT 39.610 68.765 40.110 69.145 ;
        RECT 38.715 68.085 39.045 68.585 ;
        RECT 39.215 68.255 39.385 68.755 ;
        RECT 40.280 68.470 40.450 69.315 ;
        RECT 41.380 69.155 41.630 69.315 ;
        RECT 40.620 68.885 40.870 69.145 ;
        RECT 41.800 68.885 41.990 69.655 ;
        RECT 40.620 68.635 41.990 68.885 ;
        RECT 42.160 69.825 43.410 69.995 ;
        RECT 42.160 69.065 42.330 69.825 ;
        RECT 43.080 69.705 43.410 69.825 ;
        RECT 42.500 69.245 42.680 69.655 ;
        RECT 43.580 69.485 43.750 70.245 ;
        RECT 43.950 70.155 44.610 70.635 ;
        RECT 44.790 70.040 45.110 70.370 ;
        RECT 43.940 69.715 44.600 69.985 ;
        RECT 43.940 69.655 44.270 69.715 ;
        RECT 44.420 69.485 44.750 69.545 ;
        RECT 42.850 69.315 44.750 69.485 ;
        RECT 42.160 68.755 42.680 69.065 ;
        RECT 42.850 68.805 43.020 69.315 ;
        RECT 44.920 69.145 45.110 70.040 ;
        RECT 43.190 68.975 45.110 69.145 ;
        RECT 44.790 68.955 45.110 68.975 ;
        RECT 45.310 69.725 45.560 70.375 ;
        RECT 45.740 70.175 46.025 70.635 ;
        RECT 46.205 70.295 46.460 70.455 ;
        RECT 46.205 70.125 46.545 70.295 ;
        RECT 46.205 69.925 46.460 70.125 ;
        RECT 47.005 70.090 52.350 70.635 ;
        RECT 45.310 69.395 46.110 69.725 ;
        RECT 42.850 68.635 44.060 68.805 ;
        RECT 39.620 68.300 40.450 68.470 ;
        RECT 40.690 68.085 41.070 68.465 ;
        RECT 41.250 68.345 41.420 68.635 ;
        RECT 42.850 68.555 43.020 68.635 ;
        RECT 41.590 68.085 41.920 68.465 ;
        RECT 42.390 68.305 43.020 68.555 ;
        RECT 43.200 68.085 43.620 68.465 ;
        RECT 43.820 68.345 44.060 68.635 ;
        RECT 44.290 68.085 44.620 68.775 ;
        RECT 44.790 68.345 44.960 68.955 ;
        RECT 45.310 68.805 45.560 69.395 ;
        RECT 46.280 69.065 46.460 69.925 ;
        RECT 48.590 69.260 48.930 70.090 ;
        RECT 52.525 69.865 56.035 70.635 ;
        RECT 57.125 69.910 57.415 70.635 ;
        RECT 57.585 69.875 58.295 70.465 ;
        RECT 58.805 70.105 59.135 70.465 ;
        RECT 59.335 70.275 59.665 70.635 ;
        RECT 59.835 70.105 60.165 70.465 ;
        RECT 58.805 69.895 60.165 70.105 ;
        RECT 45.230 68.295 45.560 68.805 ;
        RECT 45.740 68.085 46.025 68.885 ;
        RECT 46.205 68.395 46.460 69.065 ;
        RECT 50.410 68.520 50.760 69.770 ;
        RECT 52.525 69.345 54.175 69.865 ;
        RECT 54.345 69.175 56.035 69.695 ;
        RECT 47.005 68.085 52.350 68.520 ;
        RECT 52.525 68.085 56.035 69.175 ;
        RECT 57.125 68.085 57.415 69.250 ;
        RECT 57.585 68.905 57.790 69.875 ;
        RECT 60.350 69.795 60.610 70.635 ;
        RECT 60.785 69.890 61.040 70.465 ;
        RECT 61.210 70.255 61.540 70.635 ;
        RECT 61.755 70.085 61.925 70.465 ;
        RECT 61.210 69.915 61.925 70.085 ;
        RECT 57.960 69.105 58.290 69.645 ;
        RECT 58.465 69.395 58.960 69.725 ;
        RECT 59.280 69.395 59.655 69.725 ;
        RECT 59.865 69.395 60.175 69.725 ;
        RECT 58.465 69.105 58.790 69.395 ;
        RECT 58.985 68.905 59.315 69.125 ;
        RECT 57.585 68.675 59.315 68.905 ;
        RECT 57.585 68.255 58.285 68.675 ;
        RECT 58.485 68.085 58.815 68.445 ;
        RECT 58.985 68.275 59.315 68.675 ;
        RECT 59.485 68.425 59.655 69.395 ;
        RECT 59.835 68.085 60.165 69.145 ;
        RECT 60.350 68.085 60.610 69.235 ;
        RECT 60.785 69.160 60.955 69.890 ;
        RECT 61.210 69.725 61.380 69.915 ;
        RECT 62.185 69.865 64.775 70.635 ;
        RECT 65.495 70.085 65.665 70.375 ;
        RECT 65.835 70.255 66.165 70.635 ;
        RECT 65.495 69.915 66.160 70.085 ;
        RECT 61.125 69.395 61.380 69.725 ;
        RECT 61.210 69.185 61.380 69.395 ;
        RECT 61.660 69.365 62.015 69.735 ;
        RECT 62.185 69.345 63.395 69.865 ;
        RECT 60.785 68.255 61.040 69.160 ;
        RECT 61.210 69.015 61.925 69.185 ;
        RECT 63.565 69.175 64.775 69.695 ;
        RECT 61.210 68.085 61.540 68.845 ;
        RECT 61.755 68.255 61.925 69.015 ;
        RECT 62.185 68.085 64.775 69.175 ;
        RECT 65.410 69.095 65.760 69.745 ;
        RECT 65.930 68.925 66.160 69.915 ;
        RECT 65.495 68.755 66.160 68.925 ;
        RECT 65.495 68.255 65.665 68.755 ;
        RECT 65.835 68.085 66.165 68.585 ;
        RECT 66.335 68.255 66.560 70.375 ;
        RECT 66.775 70.255 67.105 70.635 ;
        RECT 67.275 70.085 67.445 70.415 ;
        RECT 67.745 70.255 68.760 70.455 ;
        RECT 66.750 69.895 67.445 70.085 ;
        RECT 66.750 68.925 66.920 69.895 ;
        RECT 67.090 69.095 67.500 69.715 ;
        RECT 67.670 69.145 67.890 70.015 ;
        RECT 68.070 69.705 68.420 70.075 ;
        RECT 68.590 69.525 68.760 70.255 ;
        RECT 68.930 70.195 69.340 70.635 ;
        RECT 69.630 69.995 69.880 70.425 ;
        RECT 70.080 70.175 70.400 70.635 ;
        RECT 70.960 70.245 71.810 70.415 ;
        RECT 68.930 69.655 69.340 69.985 ;
        RECT 69.630 69.655 70.050 69.995 ;
        RECT 68.340 69.485 68.760 69.525 ;
        RECT 68.340 69.315 69.690 69.485 ;
        RECT 66.750 68.755 67.445 68.925 ;
        RECT 67.670 68.765 68.170 69.145 ;
        RECT 66.775 68.085 67.105 68.585 ;
        RECT 67.275 68.255 67.445 68.755 ;
        RECT 68.340 68.470 68.510 69.315 ;
        RECT 69.440 69.155 69.690 69.315 ;
        RECT 68.680 68.885 68.930 69.145 ;
        RECT 69.860 68.885 70.050 69.655 ;
        RECT 68.680 68.635 70.050 68.885 ;
        RECT 70.220 69.825 71.470 69.995 ;
        RECT 70.220 69.065 70.390 69.825 ;
        RECT 71.140 69.705 71.470 69.825 ;
        RECT 70.560 69.245 70.740 69.655 ;
        RECT 71.640 69.485 71.810 70.245 ;
        RECT 72.010 70.155 72.670 70.635 ;
        RECT 72.850 70.040 73.170 70.370 ;
        RECT 72.000 69.715 72.660 69.985 ;
        RECT 72.000 69.655 72.330 69.715 ;
        RECT 72.480 69.485 72.810 69.545 ;
        RECT 70.910 69.315 72.810 69.485 ;
        RECT 70.220 68.755 70.740 69.065 ;
        RECT 70.910 68.805 71.080 69.315 ;
        RECT 72.980 69.145 73.170 70.040 ;
        RECT 71.250 68.975 73.170 69.145 ;
        RECT 72.850 68.955 73.170 68.975 ;
        RECT 73.370 69.725 73.620 70.375 ;
        RECT 73.800 70.175 74.085 70.635 ;
        RECT 74.265 70.295 74.520 70.455 ;
        RECT 74.265 70.125 74.605 70.295 ;
        RECT 74.265 69.925 74.520 70.125 ;
        RECT 73.370 69.395 74.170 69.725 ;
        RECT 70.910 68.635 72.120 68.805 ;
        RECT 67.680 68.300 68.510 68.470 ;
        RECT 68.750 68.085 69.130 68.465 ;
        RECT 69.310 68.345 69.480 68.635 ;
        RECT 70.910 68.555 71.080 68.635 ;
        RECT 69.650 68.085 69.980 68.465 ;
        RECT 70.450 68.305 71.080 68.555 ;
        RECT 71.260 68.085 71.680 68.465 ;
        RECT 71.880 68.345 72.120 68.635 ;
        RECT 72.350 68.085 72.680 68.775 ;
        RECT 72.850 68.345 73.020 68.955 ;
        RECT 73.370 68.805 73.620 69.395 ;
        RECT 74.340 69.065 74.520 69.925 ;
        RECT 75.125 69.815 75.335 70.635 ;
        RECT 75.505 69.835 75.835 70.465 ;
        RECT 75.505 69.235 75.755 69.835 ;
        RECT 76.005 69.815 76.235 70.635 ;
        RECT 76.445 70.090 81.790 70.635 ;
        RECT 75.925 69.395 76.255 69.645 ;
        RECT 78.030 69.260 78.370 70.090 ;
        RECT 82.885 69.910 83.175 70.635 ;
        RECT 83.345 70.090 88.690 70.635 ;
        RECT 73.290 68.295 73.620 68.805 ;
        RECT 73.800 68.085 74.085 68.885 ;
        RECT 74.265 68.395 74.520 69.065 ;
        RECT 75.125 68.085 75.335 69.225 ;
        RECT 75.505 68.255 75.835 69.235 ;
        RECT 76.005 68.085 76.235 69.225 ;
        RECT 79.850 68.520 80.200 69.770 ;
        RECT 84.930 69.260 85.270 70.090 ;
        RECT 88.865 69.885 90.075 70.635 ;
        RECT 76.445 68.085 81.790 68.520 ;
        RECT 82.885 68.085 83.175 69.250 ;
        RECT 86.750 68.520 87.100 69.770 ;
        RECT 88.865 69.345 89.385 69.885 ;
        RECT 90.450 69.855 90.950 70.465 ;
        RECT 89.555 69.175 90.075 69.715 ;
        RECT 90.245 69.395 90.595 69.645 ;
        RECT 90.780 69.225 90.950 69.855 ;
        RECT 91.580 69.985 91.910 70.465 ;
        RECT 92.080 70.175 92.305 70.635 ;
        RECT 92.475 69.985 92.805 70.465 ;
        RECT 91.580 69.815 92.805 69.985 ;
        RECT 92.995 69.835 93.245 70.635 ;
        RECT 93.415 69.835 93.755 70.465 ;
        RECT 94.015 70.085 94.185 70.375 ;
        RECT 94.355 70.255 94.685 70.635 ;
        RECT 94.015 69.915 94.680 70.085 ;
        RECT 91.120 69.445 91.450 69.645 ;
        RECT 91.620 69.445 91.950 69.645 ;
        RECT 92.120 69.445 92.540 69.645 ;
        RECT 92.715 69.475 93.410 69.645 ;
        RECT 92.715 69.225 92.885 69.475 ;
        RECT 93.580 69.225 93.755 69.835 ;
        RECT 83.345 68.085 88.690 68.520 ;
        RECT 88.865 68.085 90.075 69.175 ;
        RECT 90.450 69.055 92.885 69.225 ;
        RECT 90.450 68.255 90.780 69.055 ;
        RECT 90.950 68.085 91.280 68.885 ;
        RECT 91.580 68.255 91.910 69.055 ;
        RECT 92.555 68.085 92.805 68.885 ;
        RECT 93.075 68.085 93.245 69.225 ;
        RECT 93.415 68.255 93.755 69.225 ;
        RECT 93.930 69.095 94.280 69.745 ;
        RECT 94.450 68.925 94.680 69.915 ;
        RECT 94.015 68.755 94.680 68.925 ;
        RECT 94.015 68.255 94.185 68.755 ;
        RECT 94.355 68.085 94.685 68.585 ;
        RECT 94.855 68.255 95.080 70.375 ;
        RECT 95.295 70.255 95.625 70.635 ;
        RECT 95.795 70.085 95.965 70.415 ;
        RECT 96.265 70.255 97.280 70.455 ;
        RECT 95.270 69.895 95.965 70.085 ;
        RECT 95.270 68.925 95.440 69.895 ;
        RECT 95.610 69.095 96.020 69.715 ;
        RECT 96.190 69.145 96.410 70.015 ;
        RECT 96.590 69.705 96.940 70.075 ;
        RECT 97.110 69.525 97.280 70.255 ;
        RECT 97.450 70.195 97.860 70.635 ;
        RECT 98.150 69.995 98.400 70.425 ;
        RECT 98.600 70.175 98.920 70.635 ;
        RECT 99.480 70.245 100.330 70.415 ;
        RECT 97.450 69.655 97.860 69.985 ;
        RECT 98.150 69.655 98.570 69.995 ;
        RECT 96.860 69.485 97.280 69.525 ;
        RECT 96.860 69.315 98.210 69.485 ;
        RECT 95.270 68.755 95.965 68.925 ;
        RECT 96.190 68.765 96.690 69.145 ;
        RECT 95.295 68.085 95.625 68.585 ;
        RECT 95.795 68.255 95.965 68.755 ;
        RECT 96.860 68.470 97.030 69.315 ;
        RECT 97.960 69.155 98.210 69.315 ;
        RECT 97.200 68.885 97.450 69.145 ;
        RECT 98.380 68.885 98.570 69.655 ;
        RECT 97.200 68.635 98.570 68.885 ;
        RECT 98.740 69.825 99.990 69.995 ;
        RECT 98.740 69.065 98.910 69.825 ;
        RECT 99.660 69.705 99.990 69.825 ;
        RECT 99.080 69.245 99.260 69.655 ;
        RECT 100.160 69.485 100.330 70.245 ;
        RECT 100.530 70.155 101.190 70.635 ;
        RECT 101.370 70.040 101.690 70.370 ;
        RECT 100.520 69.715 101.180 69.985 ;
        RECT 100.520 69.655 100.850 69.715 ;
        RECT 101.000 69.485 101.330 69.545 ;
        RECT 99.430 69.315 101.330 69.485 ;
        RECT 98.740 68.755 99.260 69.065 ;
        RECT 99.430 68.805 99.600 69.315 ;
        RECT 101.500 69.145 101.690 70.040 ;
        RECT 99.770 68.975 101.690 69.145 ;
        RECT 101.370 68.955 101.690 68.975 ;
        RECT 101.890 69.725 102.140 70.375 ;
        RECT 102.320 70.175 102.605 70.635 ;
        RECT 102.785 70.295 103.040 70.455 ;
        RECT 102.785 70.125 103.125 70.295 ;
        RECT 102.785 69.925 103.040 70.125 ;
        RECT 101.890 69.395 102.690 69.725 ;
        RECT 99.430 68.635 100.640 68.805 ;
        RECT 96.200 68.300 97.030 68.470 ;
        RECT 97.270 68.085 97.650 68.465 ;
        RECT 97.830 68.345 98.000 68.635 ;
        RECT 99.430 68.555 99.600 68.635 ;
        RECT 98.170 68.085 98.500 68.465 ;
        RECT 98.970 68.305 99.600 68.555 ;
        RECT 99.780 68.085 100.200 68.465 ;
        RECT 100.400 68.345 100.640 68.635 ;
        RECT 100.870 68.085 101.200 68.775 ;
        RECT 101.370 68.345 101.540 68.955 ;
        RECT 101.890 68.805 102.140 69.395 ;
        RECT 102.860 69.065 103.040 69.925 ;
        RECT 103.585 69.865 107.095 70.635 ;
        RECT 107.265 69.885 108.475 70.635 ;
        RECT 108.645 69.910 108.935 70.635 ;
        RECT 109.110 69.895 109.365 70.465 ;
        RECT 109.535 70.235 109.865 70.635 ;
        RECT 110.290 70.100 110.820 70.465 ;
        RECT 111.010 70.295 111.285 70.465 ;
        RECT 111.005 70.125 111.285 70.295 ;
        RECT 110.290 70.065 110.465 70.100 ;
        RECT 109.535 69.895 110.465 70.065 ;
        RECT 103.585 69.345 105.235 69.865 ;
        RECT 105.405 69.175 107.095 69.695 ;
        RECT 107.265 69.345 107.785 69.885 ;
        RECT 107.955 69.175 108.475 69.715 ;
        RECT 101.810 68.295 102.140 68.805 ;
        RECT 102.320 68.085 102.605 68.885 ;
        RECT 102.785 68.395 103.040 69.065 ;
        RECT 103.585 68.085 107.095 69.175 ;
        RECT 107.265 68.085 108.475 69.175 ;
        RECT 108.645 68.085 108.935 69.250 ;
        RECT 109.110 69.225 109.280 69.895 ;
        RECT 109.535 69.725 109.705 69.895 ;
        RECT 109.450 69.395 109.705 69.725 ;
        RECT 109.930 69.395 110.125 69.725 ;
        RECT 109.110 68.255 109.445 69.225 ;
        RECT 109.615 68.085 109.785 69.225 ;
        RECT 109.955 68.425 110.125 69.395 ;
        RECT 110.295 68.765 110.465 69.895 ;
        RECT 110.635 69.105 110.805 69.905 ;
        RECT 111.010 69.305 111.285 70.125 ;
        RECT 111.455 69.105 111.645 70.465 ;
        RECT 111.825 70.100 112.335 70.635 ;
        RECT 112.555 69.825 112.800 70.430 ;
        RECT 113.245 69.865 116.755 70.635 ;
        RECT 117.385 69.885 118.595 70.635 ;
        RECT 111.845 69.655 113.075 69.825 ;
        RECT 110.635 68.935 111.645 69.105 ;
        RECT 111.815 69.090 112.565 69.280 ;
        RECT 110.295 68.595 111.420 68.765 ;
        RECT 111.815 68.425 111.985 69.090 ;
        RECT 112.735 68.845 113.075 69.655 ;
        RECT 113.245 69.345 114.895 69.865 ;
        RECT 115.065 69.175 116.755 69.695 ;
        RECT 109.955 68.255 111.985 68.425 ;
        RECT 112.155 68.085 112.325 68.845 ;
        RECT 112.560 68.435 113.075 68.845 ;
        RECT 113.245 68.085 116.755 69.175 ;
        RECT 117.385 69.175 117.905 69.715 ;
        RECT 118.075 69.345 118.595 69.885 ;
        RECT 117.385 68.085 118.595 69.175 ;
        RECT 5.520 67.915 118.680 68.085 ;
        RECT 5.605 66.825 6.815 67.915 ;
        RECT 6.985 67.480 12.330 67.915 ;
        RECT 5.605 66.115 6.125 66.655 ;
        RECT 6.295 66.285 6.815 66.825 ;
        RECT 5.605 65.365 6.815 66.115 ;
        RECT 8.570 65.910 8.910 66.740 ;
        RECT 10.390 66.230 10.740 67.480 ;
        RECT 12.505 66.825 14.175 67.915 ;
        RECT 12.505 66.135 13.255 66.655 ;
        RECT 13.425 66.305 14.175 66.825 ;
        RECT 14.495 66.765 14.825 67.915 ;
        RECT 14.995 66.895 15.165 67.745 ;
        RECT 15.335 67.115 15.665 67.915 ;
        RECT 15.835 66.895 16.005 67.745 ;
        RECT 16.185 67.115 16.425 67.915 ;
        RECT 16.595 66.935 16.925 67.745 ;
        RECT 14.995 66.725 16.005 66.895 ;
        RECT 16.210 66.765 16.925 66.935 ;
        RECT 17.105 66.825 18.315 67.915 ;
        RECT 14.995 66.185 15.490 66.725 ;
        RECT 16.210 66.525 16.380 66.765 ;
        RECT 15.880 66.355 16.380 66.525 ;
        RECT 16.550 66.355 16.930 66.595 ;
        RECT 16.210 66.185 16.380 66.355 ;
        RECT 6.985 65.365 12.330 65.910 ;
        RECT 12.505 65.365 14.175 66.135 ;
        RECT 14.495 65.365 14.825 66.165 ;
        RECT 14.995 66.015 16.005 66.185 ;
        RECT 16.210 66.015 16.845 66.185 ;
        RECT 14.995 65.535 15.165 66.015 ;
        RECT 15.335 65.365 15.665 65.845 ;
        RECT 15.835 65.535 16.005 66.015 ;
        RECT 16.255 65.365 16.495 65.845 ;
        RECT 16.675 65.535 16.845 66.015 ;
        RECT 17.105 66.115 17.625 66.655 ;
        RECT 17.795 66.285 18.315 66.825 ;
        RECT 18.485 66.750 18.775 67.915 ;
        RECT 18.945 66.825 22.455 67.915 ;
        RECT 18.945 66.135 20.595 66.655 ;
        RECT 20.765 66.305 22.455 66.825 ;
        RECT 22.625 66.775 22.965 67.745 ;
        RECT 23.135 66.775 23.305 67.915 ;
        RECT 23.575 67.115 23.825 67.915 ;
        RECT 24.470 66.945 24.800 67.745 ;
        RECT 25.100 67.115 25.430 67.915 ;
        RECT 25.600 66.945 25.930 67.745 ;
        RECT 23.495 66.775 25.930 66.945 ;
        RECT 26.510 66.945 26.840 67.745 ;
        RECT 27.010 67.115 27.340 67.915 ;
        RECT 27.640 66.945 27.970 67.745 ;
        RECT 28.615 67.115 28.865 67.915 ;
        RECT 26.510 66.775 28.945 66.945 ;
        RECT 29.135 66.775 29.305 67.915 ;
        RECT 29.475 66.775 29.815 67.745 ;
        RECT 29.985 66.825 31.655 67.915 ;
        RECT 22.625 66.165 22.800 66.775 ;
        RECT 23.495 66.525 23.665 66.775 ;
        RECT 22.970 66.355 23.665 66.525 ;
        RECT 23.840 66.355 24.260 66.555 ;
        RECT 24.430 66.355 24.760 66.555 ;
        RECT 24.930 66.355 25.260 66.555 ;
        RECT 17.105 65.365 18.315 66.115 ;
        RECT 18.485 65.365 18.775 66.090 ;
        RECT 18.945 65.365 22.455 66.135 ;
        RECT 22.625 65.535 22.965 66.165 ;
        RECT 23.135 65.365 23.385 66.165 ;
        RECT 23.575 66.015 24.800 66.185 ;
        RECT 23.575 65.535 23.905 66.015 ;
        RECT 24.075 65.365 24.300 65.825 ;
        RECT 24.470 65.535 24.800 66.015 ;
        RECT 25.430 66.145 25.600 66.775 ;
        RECT 25.785 66.355 26.135 66.605 ;
        RECT 26.305 66.355 26.655 66.605 ;
        RECT 26.840 66.145 27.010 66.775 ;
        RECT 27.180 66.355 27.510 66.555 ;
        RECT 27.680 66.355 28.010 66.555 ;
        RECT 28.180 66.355 28.600 66.555 ;
        RECT 28.775 66.525 28.945 66.775 ;
        RECT 28.775 66.355 29.470 66.525 ;
        RECT 25.430 65.535 25.930 66.145 ;
        RECT 26.510 65.535 27.010 66.145 ;
        RECT 27.640 66.015 28.865 66.185 ;
        RECT 29.640 66.165 29.815 66.775 ;
        RECT 27.640 65.535 27.970 66.015 ;
        RECT 28.140 65.365 28.365 65.825 ;
        RECT 28.535 65.535 28.865 66.015 ;
        RECT 29.055 65.365 29.305 66.165 ;
        RECT 29.475 65.535 29.815 66.165 ;
        RECT 29.985 66.135 30.735 66.655 ;
        RECT 30.905 66.305 31.655 66.825 ;
        RECT 32.285 66.775 32.625 67.745 ;
        RECT 32.795 66.775 32.965 67.915 ;
        RECT 33.235 67.115 33.485 67.915 ;
        RECT 34.130 66.945 34.460 67.745 ;
        RECT 34.760 67.115 35.090 67.915 ;
        RECT 35.260 66.945 35.590 67.745 ;
        RECT 35.965 67.480 41.310 67.915 ;
        RECT 33.155 66.775 35.590 66.945 ;
        RECT 32.285 66.165 32.460 66.775 ;
        RECT 33.155 66.525 33.325 66.775 ;
        RECT 32.630 66.355 33.325 66.525 ;
        RECT 33.500 66.355 33.920 66.555 ;
        RECT 34.090 66.355 34.420 66.555 ;
        RECT 34.590 66.355 34.920 66.555 ;
        RECT 29.985 65.365 31.655 66.135 ;
        RECT 32.285 65.535 32.625 66.165 ;
        RECT 32.795 65.365 33.045 66.165 ;
        RECT 33.235 66.015 34.460 66.185 ;
        RECT 33.235 65.535 33.565 66.015 ;
        RECT 33.735 65.365 33.960 65.825 ;
        RECT 34.130 65.535 34.460 66.015 ;
        RECT 35.090 66.145 35.260 66.775 ;
        RECT 35.445 66.355 35.795 66.605 ;
        RECT 35.090 65.535 35.590 66.145 ;
        RECT 37.550 65.910 37.890 66.740 ;
        RECT 39.370 66.230 39.720 67.480 ;
        RECT 41.485 66.825 44.075 67.915 ;
        RECT 41.485 66.135 42.695 66.655 ;
        RECT 42.865 66.305 44.075 66.825 ;
        RECT 44.245 66.750 44.535 67.915 ;
        RECT 44.705 66.825 48.215 67.915 ;
        RECT 44.705 66.135 46.355 66.655 ;
        RECT 46.525 66.305 48.215 66.825 ;
        RECT 49.510 66.945 49.840 67.745 ;
        RECT 50.010 67.115 50.340 67.915 ;
        RECT 50.640 66.945 50.970 67.745 ;
        RECT 51.615 67.115 51.865 67.915 ;
        RECT 49.510 66.775 51.945 66.945 ;
        RECT 52.135 66.775 52.305 67.915 ;
        RECT 52.475 66.775 52.815 67.745 ;
        RECT 53.190 66.945 53.520 67.745 ;
        RECT 53.690 67.115 54.020 67.915 ;
        RECT 54.320 66.945 54.650 67.745 ;
        RECT 55.295 67.115 55.545 67.915 ;
        RECT 53.190 66.775 55.625 66.945 ;
        RECT 55.815 66.775 55.985 67.915 ;
        RECT 56.155 66.775 56.495 67.745 ;
        RECT 56.665 66.825 58.335 67.915 ;
        RECT 58.515 67.105 58.810 67.915 ;
        RECT 49.305 66.355 49.655 66.605 ;
        RECT 49.840 66.145 50.010 66.775 ;
        RECT 50.180 66.355 50.510 66.555 ;
        RECT 50.680 66.355 51.010 66.555 ;
        RECT 51.180 66.355 51.600 66.555 ;
        RECT 51.775 66.525 51.945 66.775 ;
        RECT 51.775 66.355 52.470 66.525 ;
        RECT 35.965 65.365 41.310 65.910 ;
        RECT 41.485 65.365 44.075 66.135 ;
        RECT 44.245 65.365 44.535 66.090 ;
        RECT 44.705 65.365 48.215 66.135 ;
        RECT 49.510 65.535 50.010 66.145 ;
        RECT 50.640 66.015 51.865 66.185 ;
        RECT 52.640 66.165 52.815 66.775 ;
        RECT 52.985 66.355 53.335 66.605 ;
        RECT 50.640 65.535 50.970 66.015 ;
        RECT 51.140 65.365 51.365 65.825 ;
        RECT 51.535 65.535 51.865 66.015 ;
        RECT 52.055 65.365 52.305 66.165 ;
        RECT 52.475 65.535 52.815 66.165 ;
        RECT 53.520 66.145 53.690 66.775 ;
        RECT 53.860 66.355 54.190 66.555 ;
        RECT 54.360 66.355 54.690 66.555 ;
        RECT 54.860 66.355 55.280 66.555 ;
        RECT 55.455 66.525 55.625 66.775 ;
        RECT 55.455 66.355 56.150 66.525 ;
        RECT 53.190 65.535 53.690 66.145 ;
        RECT 54.320 66.015 55.545 66.185 ;
        RECT 56.320 66.165 56.495 66.775 ;
        RECT 54.320 65.535 54.650 66.015 ;
        RECT 54.820 65.365 55.045 65.825 ;
        RECT 55.215 65.535 55.545 66.015 ;
        RECT 55.735 65.365 55.985 66.165 ;
        RECT 56.155 65.535 56.495 66.165 ;
        RECT 56.665 66.135 57.415 66.655 ;
        RECT 57.585 66.305 58.335 66.825 ;
        RECT 58.990 66.605 59.235 67.745 ;
        RECT 59.410 67.105 59.670 67.915 ;
        RECT 60.270 67.910 66.545 67.915 ;
        RECT 59.850 66.605 60.100 67.740 ;
        RECT 60.270 67.115 60.530 67.910 ;
        RECT 60.700 67.015 60.960 67.740 ;
        RECT 61.130 67.185 61.390 67.910 ;
        RECT 61.560 67.015 61.820 67.740 ;
        RECT 61.990 67.185 62.250 67.910 ;
        RECT 62.420 67.015 62.680 67.740 ;
        RECT 62.850 67.185 63.110 67.910 ;
        RECT 63.280 67.015 63.540 67.740 ;
        RECT 63.710 67.185 63.955 67.910 ;
        RECT 64.125 67.015 64.385 67.740 ;
        RECT 64.570 67.185 64.815 67.910 ;
        RECT 64.985 67.015 65.245 67.740 ;
        RECT 65.430 67.185 65.675 67.910 ;
        RECT 65.845 67.015 66.105 67.740 ;
        RECT 66.290 67.185 66.545 67.910 ;
        RECT 60.700 67.000 66.105 67.015 ;
        RECT 66.715 67.000 67.005 67.740 ;
        RECT 67.175 67.170 67.445 67.915 ;
        RECT 60.700 66.895 67.445 67.000 ;
        RECT 60.700 66.775 67.475 66.895 ;
        RECT 67.705 66.825 69.375 67.915 ;
        RECT 66.280 66.725 67.475 66.775 ;
        RECT 56.665 65.365 58.335 66.135 ;
        RECT 58.505 66.045 58.820 66.605 ;
        RECT 58.990 66.355 66.110 66.605 ;
        RECT 58.505 65.365 58.810 65.875 ;
        RECT 58.990 65.545 59.240 66.355 ;
        RECT 59.410 65.365 59.670 65.890 ;
        RECT 59.850 65.545 60.100 66.355 ;
        RECT 66.280 66.185 67.445 66.725 ;
        RECT 60.700 66.015 67.445 66.185 ;
        RECT 67.705 66.135 68.455 66.655 ;
        RECT 68.625 66.305 69.375 66.825 ;
        RECT 70.005 66.750 70.295 67.915 ;
        RECT 70.555 67.245 70.725 67.745 ;
        RECT 70.895 67.415 71.225 67.915 ;
        RECT 70.555 67.075 71.220 67.245 ;
        RECT 70.470 66.255 70.820 66.905 ;
        RECT 60.270 65.365 60.530 65.925 ;
        RECT 60.700 65.560 60.960 66.015 ;
        RECT 61.130 65.365 61.390 65.845 ;
        RECT 61.560 65.560 61.820 66.015 ;
        RECT 61.990 65.365 62.250 65.845 ;
        RECT 62.420 65.560 62.680 66.015 ;
        RECT 62.850 65.365 63.095 65.845 ;
        RECT 63.265 65.560 63.540 66.015 ;
        RECT 63.710 65.365 63.955 65.845 ;
        RECT 64.125 65.560 64.385 66.015 ;
        RECT 64.565 65.365 64.815 65.845 ;
        RECT 64.985 65.560 65.245 66.015 ;
        RECT 65.425 65.365 65.675 65.845 ;
        RECT 65.845 65.560 66.105 66.015 ;
        RECT 66.285 65.365 66.545 65.845 ;
        RECT 66.715 65.560 66.975 66.015 ;
        RECT 67.145 65.365 67.445 65.845 ;
        RECT 67.705 65.365 69.375 66.135 ;
        RECT 70.005 65.365 70.295 66.090 ;
        RECT 70.990 66.085 71.220 67.075 ;
        RECT 70.555 65.915 71.220 66.085 ;
        RECT 70.555 65.625 70.725 65.915 ;
        RECT 70.895 65.365 71.225 65.745 ;
        RECT 71.395 65.625 71.620 67.745 ;
        RECT 71.835 67.415 72.165 67.915 ;
        RECT 72.335 67.245 72.505 67.745 ;
        RECT 72.740 67.530 73.570 67.700 ;
        RECT 73.810 67.535 74.190 67.915 ;
        RECT 71.810 67.075 72.505 67.245 ;
        RECT 71.810 66.105 71.980 67.075 ;
        RECT 72.150 66.285 72.560 66.905 ;
        RECT 72.730 66.855 73.230 67.235 ;
        RECT 71.810 65.915 72.505 66.105 ;
        RECT 72.730 65.985 72.950 66.855 ;
        RECT 73.400 66.685 73.570 67.530 ;
        RECT 74.370 67.365 74.540 67.655 ;
        RECT 74.710 67.535 75.040 67.915 ;
        RECT 75.510 67.445 76.140 67.695 ;
        RECT 76.320 67.535 76.740 67.915 ;
        RECT 75.970 67.365 76.140 67.445 ;
        RECT 76.940 67.365 77.180 67.655 ;
        RECT 73.740 67.115 75.110 67.365 ;
        RECT 73.740 66.855 73.990 67.115 ;
        RECT 74.500 66.685 74.750 66.845 ;
        RECT 73.400 66.515 74.750 66.685 ;
        RECT 73.400 66.475 73.820 66.515 ;
        RECT 73.130 65.925 73.480 66.295 ;
        RECT 71.835 65.365 72.165 65.745 ;
        RECT 72.335 65.585 72.505 65.915 ;
        RECT 73.650 65.745 73.820 66.475 ;
        RECT 74.920 66.345 75.110 67.115 ;
        RECT 73.990 66.015 74.400 66.345 ;
        RECT 74.690 66.005 75.110 66.345 ;
        RECT 75.280 66.935 75.800 67.245 ;
        RECT 75.970 67.195 77.180 67.365 ;
        RECT 77.410 67.225 77.740 67.915 ;
        RECT 75.280 66.175 75.450 66.935 ;
        RECT 75.620 66.345 75.800 66.755 ;
        RECT 75.970 66.685 76.140 67.195 ;
        RECT 77.910 67.045 78.080 67.655 ;
        RECT 78.350 67.195 78.680 67.705 ;
        RECT 77.910 67.025 78.230 67.045 ;
        RECT 76.310 66.855 78.230 67.025 ;
        RECT 75.970 66.515 77.870 66.685 ;
        RECT 76.200 66.175 76.530 66.295 ;
        RECT 75.280 66.005 76.530 66.175 ;
        RECT 72.805 65.545 73.820 65.745 ;
        RECT 73.990 65.365 74.400 65.805 ;
        RECT 74.690 65.575 74.940 66.005 ;
        RECT 75.140 65.365 75.460 65.825 ;
        RECT 76.700 65.755 76.870 66.515 ;
        RECT 77.540 66.455 77.870 66.515 ;
        RECT 77.060 66.285 77.390 66.345 ;
        RECT 77.060 66.015 77.720 66.285 ;
        RECT 78.040 65.960 78.230 66.855 ;
        RECT 76.020 65.585 76.870 65.755 ;
        RECT 77.070 65.365 77.730 65.845 ;
        RECT 77.910 65.630 78.230 65.960 ;
        RECT 78.430 66.605 78.680 67.195 ;
        RECT 78.860 67.115 79.145 67.915 ;
        RECT 79.325 67.575 79.580 67.605 ;
        RECT 79.325 67.405 79.665 67.575 ;
        RECT 79.325 66.935 79.580 67.405 ;
        RECT 78.430 66.275 79.230 66.605 ;
        RECT 78.430 65.625 78.680 66.275 ;
        RECT 79.400 66.075 79.580 66.935 ;
        RECT 80.125 66.825 81.795 67.915 ;
        RECT 78.860 65.365 79.145 65.825 ;
        RECT 79.325 65.545 79.580 66.075 ;
        RECT 80.125 66.135 80.875 66.655 ;
        RECT 81.045 66.305 81.795 66.825 ;
        RECT 82.630 66.945 82.960 67.745 ;
        RECT 83.130 67.115 83.460 67.915 ;
        RECT 83.760 66.945 84.090 67.745 ;
        RECT 84.735 67.115 84.985 67.915 ;
        RECT 82.630 66.775 85.065 66.945 ;
        RECT 85.255 66.775 85.425 67.915 ;
        RECT 85.595 66.775 85.935 67.745 ;
        RECT 86.310 66.945 86.640 67.745 ;
        RECT 86.810 67.115 87.140 67.915 ;
        RECT 87.440 66.945 87.770 67.745 ;
        RECT 88.415 67.115 88.665 67.915 ;
        RECT 86.310 66.775 88.745 66.945 ;
        RECT 88.935 66.775 89.105 67.915 ;
        RECT 89.275 66.775 89.615 67.745 ;
        RECT 89.990 66.945 90.320 67.745 ;
        RECT 90.490 67.115 90.820 67.915 ;
        RECT 91.120 66.945 91.450 67.745 ;
        RECT 92.095 67.115 92.345 67.915 ;
        RECT 89.990 66.775 92.425 66.945 ;
        RECT 92.615 66.775 92.785 67.915 ;
        RECT 92.955 66.775 93.295 67.745 ;
        RECT 93.465 66.825 95.135 67.915 ;
        RECT 82.425 66.355 82.775 66.605 ;
        RECT 82.960 66.145 83.130 66.775 ;
        RECT 83.300 66.355 83.630 66.555 ;
        RECT 83.800 66.355 84.130 66.555 ;
        RECT 84.300 66.355 84.720 66.555 ;
        RECT 84.895 66.525 85.065 66.775 ;
        RECT 84.895 66.355 85.590 66.525 ;
        RECT 80.125 65.365 81.795 66.135 ;
        RECT 82.630 65.535 83.130 66.145 ;
        RECT 83.760 66.015 84.985 66.185 ;
        RECT 85.760 66.165 85.935 66.775 ;
        RECT 86.105 66.355 86.455 66.605 ;
        RECT 83.760 65.535 84.090 66.015 ;
        RECT 84.260 65.365 84.485 65.825 ;
        RECT 84.655 65.535 84.985 66.015 ;
        RECT 85.175 65.365 85.425 66.165 ;
        RECT 85.595 65.535 85.935 66.165 ;
        RECT 86.640 66.145 86.810 66.775 ;
        RECT 86.980 66.355 87.310 66.555 ;
        RECT 87.480 66.355 87.810 66.555 ;
        RECT 87.980 66.355 88.400 66.555 ;
        RECT 88.575 66.525 88.745 66.775 ;
        RECT 88.575 66.355 89.270 66.525 ;
        RECT 86.310 65.535 86.810 66.145 ;
        RECT 87.440 66.015 88.665 66.185 ;
        RECT 89.440 66.165 89.615 66.775 ;
        RECT 89.785 66.355 90.135 66.605 ;
        RECT 87.440 65.535 87.770 66.015 ;
        RECT 87.940 65.365 88.165 65.825 ;
        RECT 88.335 65.535 88.665 66.015 ;
        RECT 88.855 65.365 89.105 66.165 ;
        RECT 89.275 65.535 89.615 66.165 ;
        RECT 90.320 66.145 90.490 66.775 ;
        RECT 90.660 66.355 90.990 66.555 ;
        RECT 91.160 66.355 91.490 66.555 ;
        RECT 91.660 66.355 92.080 66.555 ;
        RECT 92.255 66.525 92.425 66.775 ;
        RECT 92.255 66.355 92.950 66.525 ;
        RECT 89.990 65.535 90.490 66.145 ;
        RECT 91.120 66.015 92.345 66.185 ;
        RECT 93.120 66.165 93.295 66.775 ;
        RECT 91.120 65.535 91.450 66.015 ;
        RECT 91.620 65.365 91.845 65.825 ;
        RECT 92.015 65.535 92.345 66.015 ;
        RECT 92.535 65.365 92.785 66.165 ;
        RECT 92.955 65.535 93.295 66.165 ;
        RECT 93.465 66.135 94.215 66.655 ;
        RECT 94.385 66.305 95.135 66.825 ;
        RECT 95.765 66.750 96.055 67.915 ;
        RECT 96.230 66.775 96.565 67.745 ;
        RECT 96.735 66.775 96.905 67.915 ;
        RECT 97.075 67.575 99.105 67.745 ;
        RECT 93.465 65.365 95.135 66.135 ;
        RECT 96.230 66.105 96.400 66.775 ;
        RECT 97.075 66.605 97.245 67.575 ;
        RECT 96.570 66.275 96.825 66.605 ;
        RECT 97.050 66.275 97.245 66.605 ;
        RECT 97.415 67.235 98.540 67.405 ;
        RECT 96.655 66.105 96.825 66.275 ;
        RECT 97.415 66.105 97.585 67.235 ;
        RECT 95.765 65.365 96.055 66.090 ;
        RECT 96.230 65.535 96.485 66.105 ;
        RECT 96.655 65.935 97.585 66.105 ;
        RECT 97.755 66.895 98.765 67.065 ;
        RECT 97.755 66.095 97.925 66.895 ;
        RECT 97.410 65.900 97.585 65.935 ;
        RECT 96.655 65.365 96.985 65.765 ;
        RECT 97.410 65.535 97.940 65.900 ;
        RECT 98.130 65.875 98.405 66.695 ;
        RECT 98.125 65.705 98.405 65.875 ;
        RECT 98.130 65.535 98.405 65.705 ;
        RECT 98.575 65.535 98.765 66.895 ;
        RECT 98.935 66.910 99.105 67.575 ;
        RECT 99.275 67.155 99.445 67.915 ;
        RECT 99.680 67.155 100.195 67.565 ;
        RECT 98.935 66.720 99.685 66.910 ;
        RECT 99.855 66.345 100.195 67.155 ;
        RECT 100.365 66.825 103.875 67.915 ;
        RECT 104.045 66.825 105.255 67.915 ;
        RECT 98.965 66.175 100.195 66.345 ;
        RECT 98.945 65.365 99.455 65.900 ;
        RECT 99.675 65.570 99.920 66.175 ;
        RECT 100.365 66.135 102.015 66.655 ;
        RECT 102.185 66.305 103.875 66.825 ;
        RECT 100.365 65.365 103.875 66.135 ;
        RECT 104.045 66.115 104.565 66.655 ;
        RECT 104.735 66.285 105.255 66.825 ;
        RECT 105.515 66.985 105.685 67.745 ;
        RECT 105.865 67.155 106.195 67.915 ;
        RECT 105.515 66.815 106.180 66.985 ;
        RECT 106.365 66.840 106.635 67.745 ;
        RECT 106.895 67.245 107.065 67.745 ;
        RECT 107.235 67.415 107.565 67.915 ;
        RECT 106.895 67.075 107.560 67.245 ;
        RECT 106.010 66.670 106.180 66.815 ;
        RECT 105.445 66.265 105.775 66.635 ;
        RECT 106.010 66.340 106.295 66.670 ;
        RECT 104.045 65.365 105.255 66.115 ;
        RECT 106.010 66.085 106.180 66.340 ;
        RECT 105.515 65.915 106.180 66.085 ;
        RECT 106.465 66.040 106.635 66.840 ;
        RECT 106.810 66.255 107.160 66.905 ;
        RECT 107.330 66.085 107.560 67.075 ;
        RECT 105.515 65.535 105.685 65.915 ;
        RECT 105.865 65.365 106.195 65.745 ;
        RECT 106.375 65.535 106.635 66.040 ;
        RECT 106.895 65.915 107.560 66.085 ;
        RECT 106.895 65.625 107.065 65.915 ;
        RECT 107.235 65.365 107.565 65.745 ;
        RECT 107.735 65.625 107.960 67.745 ;
        RECT 108.175 67.415 108.505 67.915 ;
        RECT 108.675 67.245 108.845 67.745 ;
        RECT 109.080 67.530 109.910 67.700 ;
        RECT 110.150 67.535 110.530 67.915 ;
        RECT 108.150 67.075 108.845 67.245 ;
        RECT 108.150 66.105 108.320 67.075 ;
        RECT 108.490 66.285 108.900 66.905 ;
        RECT 109.070 66.855 109.570 67.235 ;
        RECT 108.150 65.915 108.845 66.105 ;
        RECT 109.070 65.985 109.290 66.855 ;
        RECT 109.740 66.685 109.910 67.530 ;
        RECT 110.710 67.365 110.880 67.655 ;
        RECT 111.050 67.535 111.380 67.915 ;
        RECT 111.850 67.445 112.480 67.695 ;
        RECT 112.660 67.535 113.080 67.915 ;
        RECT 112.310 67.365 112.480 67.445 ;
        RECT 113.280 67.365 113.520 67.655 ;
        RECT 110.080 67.115 111.450 67.365 ;
        RECT 110.080 66.855 110.330 67.115 ;
        RECT 110.840 66.685 111.090 66.845 ;
        RECT 109.740 66.515 111.090 66.685 ;
        RECT 109.740 66.475 110.160 66.515 ;
        RECT 109.470 65.925 109.820 66.295 ;
        RECT 108.175 65.365 108.505 65.745 ;
        RECT 108.675 65.585 108.845 65.915 ;
        RECT 109.990 65.745 110.160 66.475 ;
        RECT 111.260 66.345 111.450 67.115 ;
        RECT 110.330 66.015 110.740 66.345 ;
        RECT 111.030 66.005 111.450 66.345 ;
        RECT 111.620 66.935 112.140 67.245 ;
        RECT 112.310 67.195 113.520 67.365 ;
        RECT 113.750 67.225 114.080 67.915 ;
        RECT 111.620 66.175 111.790 66.935 ;
        RECT 111.960 66.345 112.140 66.755 ;
        RECT 112.310 66.685 112.480 67.195 ;
        RECT 114.250 67.045 114.420 67.655 ;
        RECT 114.690 67.195 115.020 67.705 ;
        RECT 114.250 67.025 114.570 67.045 ;
        RECT 112.650 66.855 114.570 67.025 ;
        RECT 112.310 66.515 114.210 66.685 ;
        RECT 112.540 66.175 112.870 66.295 ;
        RECT 111.620 66.005 112.870 66.175 ;
        RECT 109.145 65.545 110.160 65.745 ;
        RECT 110.330 65.365 110.740 65.805 ;
        RECT 111.030 65.575 111.280 66.005 ;
        RECT 111.480 65.365 111.800 65.825 ;
        RECT 113.040 65.755 113.210 66.515 ;
        RECT 113.880 66.455 114.210 66.515 ;
        RECT 113.400 66.285 113.730 66.345 ;
        RECT 113.400 66.015 114.060 66.285 ;
        RECT 114.380 65.960 114.570 66.855 ;
        RECT 112.360 65.585 113.210 65.755 ;
        RECT 113.410 65.365 114.070 65.845 ;
        RECT 114.250 65.630 114.570 65.960 ;
        RECT 114.770 66.605 115.020 67.195 ;
        RECT 115.200 67.115 115.485 67.915 ;
        RECT 115.665 66.935 115.920 67.605 ;
        RECT 114.770 66.275 115.570 66.605 ;
        RECT 114.770 65.625 115.020 66.275 ;
        RECT 115.740 66.075 115.920 66.935 ;
        RECT 117.385 66.825 118.595 67.915 ;
        RECT 117.385 66.285 117.905 66.825 ;
        RECT 118.075 66.115 118.595 66.655 ;
        RECT 115.665 65.875 115.920 66.075 ;
        RECT 115.200 65.365 115.485 65.825 ;
        RECT 115.665 65.705 116.005 65.875 ;
        RECT 115.665 65.545 115.920 65.705 ;
        RECT 117.385 65.365 118.595 66.115 ;
        RECT 5.520 65.195 118.680 65.365 ;
        RECT 5.605 64.445 6.815 65.195 ;
        RECT 6.985 64.650 12.330 65.195 ;
        RECT 5.605 63.905 6.125 64.445 ;
        RECT 6.295 63.735 6.815 64.275 ;
        RECT 8.570 63.820 8.910 64.650 ;
        RECT 13.425 64.455 13.810 65.025 ;
        RECT 13.980 64.735 14.305 65.195 ;
        RECT 14.825 64.565 15.105 65.025 ;
        RECT 5.605 62.645 6.815 63.735 ;
        RECT 10.390 63.080 10.740 64.330 ;
        RECT 13.425 63.785 13.705 64.455 ;
        RECT 13.980 64.395 15.105 64.565 ;
        RECT 13.980 64.285 14.430 64.395 ;
        RECT 13.875 63.955 14.430 64.285 ;
        RECT 15.295 64.225 15.695 65.025 ;
        RECT 16.095 64.735 16.365 65.195 ;
        RECT 16.535 64.565 16.820 65.025 ;
        RECT 6.985 62.645 12.330 63.080 ;
        RECT 13.425 62.815 13.810 63.785 ;
        RECT 13.980 63.495 14.430 63.955 ;
        RECT 14.600 63.665 15.695 64.225 ;
        RECT 13.980 63.275 15.105 63.495 ;
        RECT 13.980 62.645 14.305 63.105 ;
        RECT 14.825 62.815 15.105 63.275 ;
        RECT 15.295 62.815 15.695 63.665 ;
        RECT 15.865 64.395 16.820 64.565 ;
        RECT 17.105 64.425 20.615 65.195 ;
        RECT 15.865 63.495 16.075 64.395 ;
        RECT 16.245 63.665 16.935 64.225 ;
        RECT 17.105 63.905 18.755 64.425 ;
        RECT 21.910 64.415 22.410 65.025 ;
        RECT 18.925 63.735 20.615 64.255 ;
        RECT 21.705 63.955 22.055 64.205 ;
        RECT 22.240 63.785 22.410 64.415 ;
        RECT 23.040 64.545 23.370 65.025 ;
        RECT 23.540 64.735 23.765 65.195 ;
        RECT 23.935 64.545 24.265 65.025 ;
        RECT 23.040 64.375 24.265 64.545 ;
        RECT 24.455 64.395 24.705 65.195 ;
        RECT 24.875 64.395 25.215 65.025 ;
        RECT 22.580 64.005 22.910 64.205 ;
        RECT 23.080 64.005 23.410 64.205 ;
        RECT 23.580 64.005 24.000 64.205 ;
        RECT 24.175 64.035 24.870 64.205 ;
        RECT 24.175 63.785 24.345 64.035 ;
        RECT 25.040 63.785 25.215 64.395 ;
        RECT 15.865 63.275 16.820 63.495 ;
        RECT 16.095 62.645 16.365 63.105 ;
        RECT 16.535 62.815 16.820 63.275 ;
        RECT 17.105 62.645 20.615 63.735 ;
        RECT 21.910 63.615 24.345 63.785 ;
        RECT 21.910 62.815 22.240 63.615 ;
        RECT 22.410 62.645 22.740 63.445 ;
        RECT 23.040 62.815 23.370 63.615 ;
        RECT 24.015 62.645 24.265 63.445 ;
        RECT 24.535 62.645 24.705 63.785 ;
        RECT 24.875 62.815 25.215 63.785 ;
        RECT 26.305 64.520 26.565 65.025 ;
        RECT 26.745 64.815 27.075 65.195 ;
        RECT 27.255 64.645 27.425 65.025 ;
        RECT 26.305 63.720 26.475 64.520 ;
        RECT 26.760 64.475 27.425 64.645 ;
        RECT 27.775 64.645 27.945 65.025 ;
        RECT 28.125 64.815 28.455 65.195 ;
        RECT 27.775 64.475 28.440 64.645 ;
        RECT 28.635 64.520 28.895 65.025 ;
        RECT 26.760 64.220 26.930 64.475 ;
        RECT 26.645 63.890 26.930 64.220 ;
        RECT 27.165 63.925 27.495 64.295 ;
        RECT 27.705 63.925 28.035 64.295 ;
        RECT 28.270 64.220 28.440 64.475 ;
        RECT 26.760 63.745 26.930 63.890 ;
        RECT 28.270 63.890 28.555 64.220 ;
        RECT 28.270 63.745 28.440 63.890 ;
        RECT 26.305 62.815 26.575 63.720 ;
        RECT 26.760 63.575 27.425 63.745 ;
        RECT 26.745 62.645 27.075 63.405 ;
        RECT 27.255 62.815 27.425 63.575 ;
        RECT 27.775 63.575 28.440 63.745 ;
        RECT 28.725 63.720 28.895 64.520 ;
        RECT 29.065 64.425 30.735 65.195 ;
        RECT 31.365 64.470 31.655 65.195 ;
        RECT 29.065 63.905 29.815 64.425 ;
        RECT 32.345 64.375 32.555 65.195 ;
        RECT 32.725 64.395 33.055 65.025 ;
        RECT 29.985 63.735 30.735 64.255 ;
        RECT 27.775 62.815 27.945 63.575 ;
        RECT 28.125 62.645 28.455 63.405 ;
        RECT 28.625 62.815 28.895 63.720 ;
        RECT 29.065 62.645 30.735 63.735 ;
        RECT 31.365 62.645 31.655 63.810 ;
        RECT 32.725 63.795 32.975 64.395 ;
        RECT 33.225 64.375 33.455 65.195 ;
        RECT 33.665 64.425 35.335 65.195 ;
        RECT 35.505 64.520 35.765 65.025 ;
        RECT 35.945 64.815 36.275 65.195 ;
        RECT 36.455 64.645 36.625 65.025 ;
        RECT 33.145 63.955 33.475 64.205 ;
        RECT 33.665 63.905 34.415 64.425 ;
        RECT 32.345 62.645 32.555 63.785 ;
        RECT 32.725 62.815 33.055 63.795 ;
        RECT 33.225 62.645 33.455 63.785 ;
        RECT 34.585 63.735 35.335 64.255 ;
        RECT 33.665 62.645 35.335 63.735 ;
        RECT 35.505 63.720 35.675 64.520 ;
        RECT 35.960 64.475 36.625 64.645 ;
        RECT 35.960 64.220 36.130 64.475 ;
        RECT 36.885 64.425 38.555 65.195 ;
        RECT 35.845 63.890 36.130 64.220 ;
        RECT 36.365 63.925 36.695 64.295 ;
        RECT 36.885 63.905 37.635 64.425 ;
        RECT 39.245 64.375 39.455 65.195 ;
        RECT 39.625 64.395 39.955 65.025 ;
        RECT 35.960 63.745 36.130 63.890 ;
        RECT 35.505 62.815 35.775 63.720 ;
        RECT 35.960 63.575 36.625 63.745 ;
        RECT 37.805 63.735 38.555 64.255 ;
        RECT 39.625 63.795 39.875 64.395 ;
        RECT 40.125 64.375 40.355 65.195 ;
        RECT 40.565 64.425 42.235 65.195 ;
        RECT 42.955 64.645 43.125 64.935 ;
        RECT 43.295 64.815 43.625 65.195 ;
        RECT 42.955 64.475 43.620 64.645 ;
        RECT 40.045 63.955 40.375 64.205 ;
        RECT 40.565 63.905 41.315 64.425 ;
        RECT 35.945 62.645 36.275 63.405 ;
        RECT 36.455 62.815 36.625 63.575 ;
        RECT 36.885 62.645 38.555 63.735 ;
        RECT 39.245 62.645 39.455 63.785 ;
        RECT 39.625 62.815 39.955 63.795 ;
        RECT 40.125 62.645 40.355 63.785 ;
        RECT 41.485 63.735 42.235 64.255 ;
        RECT 40.565 62.645 42.235 63.735 ;
        RECT 42.870 63.655 43.220 64.305 ;
        RECT 43.390 63.485 43.620 64.475 ;
        RECT 42.955 63.315 43.620 63.485 ;
        RECT 42.955 62.815 43.125 63.315 ;
        RECT 43.295 62.645 43.625 63.145 ;
        RECT 43.795 62.815 44.020 64.935 ;
        RECT 44.235 64.815 44.565 65.195 ;
        RECT 44.735 64.645 44.905 64.975 ;
        RECT 45.205 64.815 46.220 65.015 ;
        RECT 44.210 64.455 44.905 64.645 ;
        RECT 44.210 63.485 44.380 64.455 ;
        RECT 44.550 63.655 44.960 64.275 ;
        RECT 45.130 63.705 45.350 64.575 ;
        RECT 45.530 64.265 45.880 64.635 ;
        RECT 46.050 64.085 46.220 64.815 ;
        RECT 46.390 64.755 46.800 65.195 ;
        RECT 47.090 64.555 47.340 64.985 ;
        RECT 47.540 64.735 47.860 65.195 ;
        RECT 48.420 64.805 49.270 64.975 ;
        RECT 46.390 64.215 46.800 64.545 ;
        RECT 47.090 64.215 47.510 64.555 ;
        RECT 45.800 64.045 46.220 64.085 ;
        RECT 45.800 63.875 47.150 64.045 ;
        RECT 44.210 63.315 44.905 63.485 ;
        RECT 45.130 63.325 45.630 63.705 ;
        RECT 44.235 62.645 44.565 63.145 ;
        RECT 44.735 62.815 44.905 63.315 ;
        RECT 45.800 63.030 45.970 63.875 ;
        RECT 46.900 63.715 47.150 63.875 ;
        RECT 46.140 63.445 46.390 63.705 ;
        RECT 47.320 63.445 47.510 64.215 ;
        RECT 46.140 63.195 47.510 63.445 ;
        RECT 47.680 64.385 48.930 64.555 ;
        RECT 47.680 63.625 47.850 64.385 ;
        RECT 48.600 64.265 48.930 64.385 ;
        RECT 48.020 63.805 48.200 64.215 ;
        RECT 49.100 64.045 49.270 64.805 ;
        RECT 49.470 64.715 50.130 65.195 ;
        RECT 50.310 64.600 50.630 64.930 ;
        RECT 49.460 64.275 50.120 64.545 ;
        RECT 49.460 64.215 49.790 64.275 ;
        RECT 49.940 64.045 50.270 64.105 ;
        RECT 48.370 63.875 50.270 64.045 ;
        RECT 47.680 63.315 48.200 63.625 ;
        RECT 48.370 63.365 48.540 63.875 ;
        RECT 50.440 63.705 50.630 64.600 ;
        RECT 48.710 63.535 50.630 63.705 ;
        RECT 50.310 63.515 50.630 63.535 ;
        RECT 50.830 64.285 51.080 64.935 ;
        RECT 51.260 64.735 51.545 65.195 ;
        RECT 51.725 64.485 51.980 65.015 ;
        RECT 50.830 63.955 51.630 64.285 ;
        RECT 48.370 63.195 49.580 63.365 ;
        RECT 45.140 62.860 45.970 63.030 ;
        RECT 46.210 62.645 46.590 63.025 ;
        RECT 46.770 62.905 46.940 63.195 ;
        RECT 48.370 63.115 48.540 63.195 ;
        RECT 47.110 62.645 47.440 63.025 ;
        RECT 47.910 62.865 48.540 63.115 ;
        RECT 48.720 62.645 49.140 63.025 ;
        RECT 49.340 62.905 49.580 63.195 ;
        RECT 49.810 62.645 50.140 63.335 ;
        RECT 50.310 62.905 50.480 63.515 ;
        RECT 50.830 63.365 51.080 63.955 ;
        RECT 51.800 63.625 51.980 64.485 ;
        RECT 50.750 62.855 51.080 63.365 ;
        RECT 51.260 62.645 51.545 63.445 ;
        RECT 51.725 63.155 51.980 63.625 ;
        RECT 52.985 64.395 53.325 65.025 ;
        RECT 53.495 64.395 53.745 65.195 ;
        RECT 53.935 64.545 54.265 65.025 ;
        RECT 54.435 64.735 54.660 65.195 ;
        RECT 54.830 64.545 55.160 65.025 ;
        RECT 52.985 63.785 53.160 64.395 ;
        RECT 53.935 64.375 55.160 64.545 ;
        RECT 55.790 64.415 56.290 65.025 ;
        RECT 57.125 64.470 57.415 65.195 ;
        RECT 53.330 64.035 54.025 64.205 ;
        RECT 53.855 63.785 54.025 64.035 ;
        RECT 54.200 64.005 54.620 64.205 ;
        RECT 54.790 64.005 55.120 64.205 ;
        RECT 55.290 64.005 55.620 64.205 ;
        RECT 55.790 63.785 55.960 64.415 ;
        RECT 57.585 64.395 57.925 65.025 ;
        RECT 58.095 64.395 58.345 65.195 ;
        RECT 58.535 64.545 58.865 65.025 ;
        RECT 59.035 64.735 59.260 65.195 ;
        RECT 59.430 64.545 59.760 65.025 ;
        RECT 56.145 63.955 56.495 64.205 ;
        RECT 51.725 62.985 52.065 63.155 ;
        RECT 51.725 62.955 51.980 62.985 ;
        RECT 52.985 62.815 53.325 63.785 ;
        RECT 53.495 62.645 53.665 63.785 ;
        RECT 53.855 63.615 56.290 63.785 ;
        RECT 53.935 62.645 54.185 63.445 ;
        RECT 54.830 62.815 55.160 63.615 ;
        RECT 55.460 62.645 55.790 63.445 ;
        RECT 55.960 62.815 56.290 63.615 ;
        RECT 57.125 62.645 57.415 63.810 ;
        RECT 57.585 63.785 57.760 64.395 ;
        RECT 58.535 64.375 59.760 64.545 ;
        RECT 60.390 64.415 60.890 65.025 ;
        RECT 57.930 64.035 58.625 64.205 ;
        RECT 58.455 63.785 58.625 64.035 ;
        RECT 58.800 64.005 59.220 64.205 ;
        RECT 59.390 64.005 59.720 64.205 ;
        RECT 59.890 64.005 60.220 64.205 ;
        RECT 60.390 63.785 60.560 64.415 ;
        RECT 61.270 64.355 61.530 65.195 ;
        RECT 61.705 64.450 61.960 65.025 ;
        RECT 62.130 64.815 62.460 65.195 ;
        RECT 62.675 64.645 62.845 65.025 ;
        RECT 62.130 64.475 62.845 64.645 ;
        RECT 60.745 63.955 61.095 64.205 ;
        RECT 57.585 62.815 57.925 63.785 ;
        RECT 58.095 62.645 58.265 63.785 ;
        RECT 58.455 63.615 60.890 63.785 ;
        RECT 58.535 62.645 58.785 63.445 ;
        RECT 59.430 62.815 59.760 63.615 ;
        RECT 60.060 62.645 60.390 63.445 ;
        RECT 60.560 62.815 60.890 63.615 ;
        RECT 61.270 62.645 61.530 63.795 ;
        RECT 61.705 63.720 61.875 64.450 ;
        RECT 62.130 64.285 62.300 64.475 ;
        RECT 63.110 64.355 63.370 65.195 ;
        RECT 63.545 64.450 63.800 65.025 ;
        RECT 63.970 64.815 64.300 65.195 ;
        RECT 64.515 64.645 64.685 65.025 ;
        RECT 63.970 64.475 64.685 64.645 ;
        RECT 62.045 63.955 62.300 64.285 ;
        RECT 62.130 63.745 62.300 63.955 ;
        RECT 62.580 63.925 62.935 64.295 ;
        RECT 61.705 62.815 61.960 63.720 ;
        RECT 62.130 63.575 62.845 63.745 ;
        RECT 62.130 62.645 62.460 63.405 ;
        RECT 62.675 62.815 62.845 63.575 ;
        RECT 63.110 62.645 63.370 63.795 ;
        RECT 63.545 63.720 63.715 64.450 ;
        RECT 63.970 64.285 64.140 64.475 ;
        RECT 64.945 64.425 68.455 65.195 ;
        RECT 69.175 64.545 69.345 65.025 ;
        RECT 69.525 64.715 69.765 65.195 ;
        RECT 70.015 64.545 70.185 65.025 ;
        RECT 70.355 64.715 70.685 65.195 ;
        RECT 70.855 64.545 71.025 65.025 ;
        RECT 63.885 63.955 64.140 64.285 ;
        RECT 63.970 63.745 64.140 63.955 ;
        RECT 64.420 63.925 64.775 64.295 ;
        RECT 64.945 63.905 66.595 64.425 ;
        RECT 69.175 64.375 69.810 64.545 ;
        RECT 70.015 64.375 71.025 64.545 ;
        RECT 71.195 64.395 71.525 65.195 ;
        RECT 71.885 64.375 72.115 65.195 ;
        RECT 72.285 64.395 72.615 65.025 ;
        RECT 63.545 62.815 63.800 63.720 ;
        RECT 63.970 63.575 64.685 63.745 ;
        RECT 66.765 63.735 68.455 64.255 ;
        RECT 69.640 64.205 69.810 64.375 ;
        RECT 69.090 63.965 69.470 64.205 ;
        RECT 69.640 64.035 70.140 64.205 ;
        RECT 70.530 64.175 71.025 64.375 ;
        RECT 69.640 63.795 69.810 64.035 ;
        RECT 70.525 64.005 71.025 64.175 ;
        RECT 70.530 63.835 71.025 64.005 ;
        RECT 71.865 63.955 72.195 64.205 ;
        RECT 63.970 62.645 64.300 63.405 ;
        RECT 64.515 62.815 64.685 63.575 ;
        RECT 64.945 62.645 68.455 63.735 ;
        RECT 69.095 63.625 69.810 63.795 ;
        RECT 70.015 63.665 71.025 63.835 ;
        RECT 72.365 63.795 72.615 64.395 ;
        RECT 72.785 64.375 72.995 65.195 ;
        RECT 73.225 64.650 78.570 65.195 ;
        RECT 74.810 63.820 75.150 64.650 ;
        RECT 79.410 64.415 79.910 65.025 ;
        RECT 69.095 62.815 69.425 63.625 ;
        RECT 69.595 62.645 69.835 63.445 ;
        RECT 70.015 62.815 70.185 63.665 ;
        RECT 70.355 62.645 70.685 63.445 ;
        RECT 70.855 62.815 71.025 63.665 ;
        RECT 71.195 62.645 71.525 63.795 ;
        RECT 71.885 62.645 72.115 63.785 ;
        RECT 72.285 62.815 72.615 63.795 ;
        RECT 72.785 62.645 72.995 63.785 ;
        RECT 76.630 63.080 76.980 64.330 ;
        RECT 79.205 63.955 79.555 64.205 ;
        RECT 79.740 63.785 79.910 64.415 ;
        RECT 80.540 64.545 80.870 65.025 ;
        RECT 81.040 64.735 81.265 65.195 ;
        RECT 81.435 64.545 81.765 65.025 ;
        RECT 80.540 64.375 81.765 64.545 ;
        RECT 81.955 64.395 82.205 65.195 ;
        RECT 82.375 64.395 82.715 65.025 ;
        RECT 82.885 64.470 83.175 65.195 ;
        RECT 80.080 64.005 80.410 64.205 ;
        RECT 80.580 64.005 80.910 64.205 ;
        RECT 81.080 64.005 81.500 64.205 ;
        RECT 81.675 64.035 82.370 64.205 ;
        RECT 81.675 63.785 81.845 64.035 ;
        RECT 82.540 63.785 82.715 64.395 ;
        RECT 83.345 64.455 83.730 65.025 ;
        RECT 83.900 64.735 84.225 65.195 ;
        RECT 84.745 64.565 85.025 65.025 ;
        RECT 79.410 63.615 81.845 63.785 ;
        RECT 73.225 62.645 78.570 63.080 ;
        RECT 79.410 62.815 79.740 63.615 ;
        RECT 79.910 62.645 80.240 63.445 ;
        RECT 80.540 62.815 80.870 63.615 ;
        RECT 81.515 62.645 81.765 63.445 ;
        RECT 82.035 62.645 82.205 63.785 ;
        RECT 82.375 62.815 82.715 63.785 ;
        RECT 82.885 62.645 83.175 63.810 ;
        RECT 83.345 63.785 83.625 64.455 ;
        RECT 83.900 64.395 85.025 64.565 ;
        RECT 83.900 64.285 84.350 64.395 ;
        RECT 83.795 63.955 84.350 64.285 ;
        RECT 85.215 64.225 85.615 65.025 ;
        RECT 86.015 64.735 86.285 65.195 ;
        RECT 86.455 64.565 86.740 65.025 ;
        RECT 83.345 62.815 83.730 63.785 ;
        RECT 83.900 63.495 84.350 63.955 ;
        RECT 84.520 63.665 85.615 64.225 ;
        RECT 83.900 63.275 85.025 63.495 ;
        RECT 83.900 62.645 84.225 63.105 ;
        RECT 84.745 62.815 85.025 63.275 ;
        RECT 85.215 62.815 85.615 63.665 ;
        RECT 85.785 64.395 86.740 64.565 ;
        RECT 87.025 64.395 87.365 65.025 ;
        RECT 87.535 64.395 87.785 65.195 ;
        RECT 87.975 64.545 88.305 65.025 ;
        RECT 88.475 64.735 88.700 65.195 ;
        RECT 88.870 64.545 89.200 65.025 ;
        RECT 85.785 63.495 85.995 64.395 ;
        RECT 86.165 63.665 86.855 64.225 ;
        RECT 87.025 63.785 87.200 64.395 ;
        RECT 87.975 64.375 89.200 64.545 ;
        RECT 89.830 64.415 90.330 65.025 ;
        RECT 87.370 64.035 88.065 64.205 ;
        RECT 87.895 63.785 88.065 64.035 ;
        RECT 88.240 64.005 88.660 64.205 ;
        RECT 88.830 64.005 89.160 64.205 ;
        RECT 89.330 64.005 89.660 64.205 ;
        RECT 89.830 63.785 90.000 64.415 ;
        RECT 90.705 64.395 91.045 65.025 ;
        RECT 91.215 64.395 91.465 65.195 ;
        RECT 91.655 64.545 91.985 65.025 ;
        RECT 92.155 64.735 92.380 65.195 ;
        RECT 92.550 64.545 92.880 65.025 ;
        RECT 90.185 63.955 90.535 64.205 ;
        RECT 90.705 63.785 90.880 64.395 ;
        RECT 91.655 64.375 92.880 64.545 ;
        RECT 93.510 64.415 94.010 65.025 ;
        RECT 94.385 64.425 97.895 65.195 ;
        RECT 98.065 64.455 98.450 65.025 ;
        RECT 98.620 64.735 98.945 65.195 ;
        RECT 99.465 64.565 99.745 65.025 ;
        RECT 91.050 64.035 91.745 64.205 ;
        RECT 91.575 63.785 91.745 64.035 ;
        RECT 91.920 64.005 92.340 64.205 ;
        RECT 92.510 64.005 92.840 64.205 ;
        RECT 93.010 64.005 93.340 64.205 ;
        RECT 93.510 63.785 93.680 64.415 ;
        RECT 93.865 63.955 94.215 64.205 ;
        RECT 94.385 63.905 96.035 64.425 ;
        RECT 85.785 63.275 86.740 63.495 ;
        RECT 86.015 62.645 86.285 63.105 ;
        RECT 86.455 62.815 86.740 63.275 ;
        RECT 87.025 62.815 87.365 63.785 ;
        RECT 87.535 62.645 87.705 63.785 ;
        RECT 87.895 63.615 90.330 63.785 ;
        RECT 87.975 62.645 88.225 63.445 ;
        RECT 88.870 62.815 89.200 63.615 ;
        RECT 89.500 62.645 89.830 63.445 ;
        RECT 90.000 62.815 90.330 63.615 ;
        RECT 90.705 62.815 91.045 63.785 ;
        RECT 91.215 62.645 91.385 63.785 ;
        RECT 91.575 63.615 94.010 63.785 ;
        RECT 96.205 63.735 97.895 64.255 ;
        RECT 91.655 62.645 91.905 63.445 ;
        RECT 92.550 62.815 92.880 63.615 ;
        RECT 93.180 62.645 93.510 63.445 ;
        RECT 93.680 62.815 94.010 63.615 ;
        RECT 94.385 62.645 97.895 63.735 ;
        RECT 98.065 63.785 98.345 64.455 ;
        RECT 98.620 64.395 99.745 64.565 ;
        RECT 98.620 64.285 99.070 64.395 ;
        RECT 98.515 63.955 99.070 64.285 ;
        RECT 99.935 64.225 100.335 65.025 ;
        RECT 100.735 64.735 101.005 65.195 ;
        RECT 101.175 64.565 101.460 65.025 ;
        RECT 98.065 62.815 98.450 63.785 ;
        RECT 98.620 63.495 99.070 63.955 ;
        RECT 99.240 63.665 100.335 64.225 ;
        RECT 98.620 63.275 99.745 63.495 ;
        RECT 98.620 62.645 98.945 63.105 ;
        RECT 99.465 62.815 99.745 63.275 ;
        RECT 99.935 62.815 100.335 63.665 ;
        RECT 100.505 64.395 101.460 64.565 ;
        RECT 101.745 64.455 102.130 65.025 ;
        RECT 102.300 64.735 102.625 65.195 ;
        RECT 103.145 64.565 103.425 65.025 ;
        RECT 100.505 63.495 100.715 64.395 ;
        RECT 100.885 63.665 101.575 64.225 ;
        RECT 101.745 63.785 102.025 64.455 ;
        RECT 102.300 64.395 103.425 64.565 ;
        RECT 102.300 64.285 102.750 64.395 ;
        RECT 102.195 63.955 102.750 64.285 ;
        RECT 103.615 64.225 104.015 65.025 ;
        RECT 104.415 64.735 104.685 65.195 ;
        RECT 104.855 64.565 105.140 65.025 ;
        RECT 100.505 63.275 101.460 63.495 ;
        RECT 100.735 62.645 101.005 63.105 ;
        RECT 101.175 62.815 101.460 63.275 ;
        RECT 101.745 62.815 102.130 63.785 ;
        RECT 102.300 63.495 102.750 63.955 ;
        RECT 102.920 63.665 104.015 64.225 ;
        RECT 102.300 63.275 103.425 63.495 ;
        RECT 102.300 62.645 102.625 63.105 ;
        RECT 103.145 62.815 103.425 63.275 ;
        RECT 103.615 62.815 104.015 63.665 ;
        RECT 104.185 64.395 105.140 64.565 ;
        RECT 105.425 64.425 107.095 65.195 ;
        RECT 107.265 64.520 107.525 65.025 ;
        RECT 107.705 64.815 108.035 65.195 ;
        RECT 108.215 64.645 108.385 65.025 ;
        RECT 104.185 63.495 104.395 64.395 ;
        RECT 104.565 63.665 105.255 64.225 ;
        RECT 105.425 63.905 106.175 64.425 ;
        RECT 106.345 63.735 107.095 64.255 ;
        RECT 104.185 63.275 105.140 63.495 ;
        RECT 104.415 62.645 104.685 63.105 ;
        RECT 104.855 62.815 105.140 63.275 ;
        RECT 105.425 62.645 107.095 63.735 ;
        RECT 107.265 63.720 107.435 64.520 ;
        RECT 107.720 64.475 108.385 64.645 ;
        RECT 107.720 64.220 107.890 64.475 ;
        RECT 108.645 64.470 108.935 65.195 ;
        RECT 109.110 64.455 109.365 65.025 ;
        RECT 109.535 64.795 109.865 65.195 ;
        RECT 110.290 64.660 110.820 65.025 ;
        RECT 111.010 64.855 111.285 65.025 ;
        RECT 111.005 64.685 111.285 64.855 ;
        RECT 110.290 64.625 110.465 64.660 ;
        RECT 109.535 64.455 110.465 64.625 ;
        RECT 107.605 63.890 107.890 64.220 ;
        RECT 108.125 63.925 108.455 64.295 ;
        RECT 107.720 63.745 107.890 63.890 ;
        RECT 107.265 62.815 107.535 63.720 ;
        RECT 107.720 63.575 108.385 63.745 ;
        RECT 107.705 62.645 108.035 63.405 ;
        RECT 108.215 62.815 108.385 63.575 ;
        RECT 108.645 62.645 108.935 63.810 ;
        RECT 109.110 63.785 109.280 64.455 ;
        RECT 109.535 64.285 109.705 64.455 ;
        RECT 109.450 63.955 109.705 64.285 ;
        RECT 109.930 63.955 110.125 64.285 ;
        RECT 109.110 62.815 109.445 63.785 ;
        RECT 109.615 62.645 109.785 63.785 ;
        RECT 109.955 62.985 110.125 63.955 ;
        RECT 110.295 63.325 110.465 64.455 ;
        RECT 110.635 63.665 110.805 64.465 ;
        RECT 111.010 63.865 111.285 64.685 ;
        RECT 111.455 63.665 111.645 65.025 ;
        RECT 111.825 64.660 112.335 65.195 ;
        RECT 112.555 64.385 112.800 64.990 ;
        RECT 111.845 64.215 113.075 64.385 ;
        RECT 113.305 64.375 113.515 65.195 ;
        RECT 113.685 64.395 114.015 65.025 ;
        RECT 110.635 63.495 111.645 63.665 ;
        RECT 111.815 63.650 112.565 63.840 ;
        RECT 110.295 63.155 111.420 63.325 ;
        RECT 111.815 62.985 111.985 63.650 ;
        RECT 112.735 63.405 113.075 64.215 ;
        RECT 113.685 63.795 113.935 64.395 ;
        RECT 114.185 64.375 114.415 65.195 ;
        RECT 114.665 64.375 114.895 65.195 ;
        RECT 115.065 64.395 115.395 65.025 ;
        RECT 114.105 63.955 114.435 64.205 ;
        RECT 114.645 63.955 114.975 64.205 ;
        RECT 115.145 63.795 115.395 64.395 ;
        RECT 115.565 64.375 115.775 65.195 ;
        RECT 116.005 64.445 117.215 65.195 ;
        RECT 117.385 64.445 118.595 65.195 ;
        RECT 116.005 63.905 116.525 64.445 ;
        RECT 109.955 62.815 111.985 62.985 ;
        RECT 112.155 62.645 112.325 63.405 ;
        RECT 112.560 62.995 113.075 63.405 ;
        RECT 113.305 62.645 113.515 63.785 ;
        RECT 113.685 62.815 114.015 63.795 ;
        RECT 114.185 62.645 114.415 63.785 ;
        RECT 114.665 62.645 114.895 63.785 ;
        RECT 115.065 62.815 115.395 63.795 ;
        RECT 115.565 62.645 115.775 63.785 ;
        RECT 116.695 63.735 117.215 64.275 ;
        RECT 116.005 62.645 117.215 63.735 ;
        RECT 117.385 63.735 117.905 64.275 ;
        RECT 118.075 63.905 118.595 64.445 ;
        RECT 117.385 62.645 118.595 63.735 ;
        RECT 5.520 62.475 118.680 62.645 ;
        RECT 5.605 61.385 6.815 62.475 ;
        RECT 6.985 61.385 10.495 62.475 ;
        RECT 5.605 60.675 6.125 61.215 ;
        RECT 6.295 60.845 6.815 61.385 ;
        RECT 6.985 60.695 8.635 61.215 ;
        RECT 8.805 60.865 10.495 61.385 ;
        RECT 11.125 61.400 11.395 62.305 ;
        RECT 11.565 61.715 11.895 62.475 ;
        RECT 12.075 61.545 12.245 62.305 ;
        RECT 5.605 59.925 6.815 60.675 ;
        RECT 6.985 59.925 10.495 60.695 ;
        RECT 11.125 60.600 11.295 61.400 ;
        RECT 11.580 61.375 12.245 61.545 ;
        RECT 11.580 61.230 11.750 61.375 ;
        RECT 13.025 61.335 13.235 62.475 ;
        RECT 11.465 60.900 11.750 61.230 ;
        RECT 13.405 61.325 13.735 62.305 ;
        RECT 13.905 61.335 14.135 62.475 ;
        RECT 14.350 61.335 14.685 62.305 ;
        RECT 14.855 61.335 15.025 62.475 ;
        RECT 15.195 62.135 17.225 62.305 ;
        RECT 11.580 60.645 11.750 60.900 ;
        RECT 11.985 60.825 12.315 61.195 ;
        RECT 11.125 60.095 11.385 60.600 ;
        RECT 11.580 60.475 12.245 60.645 ;
        RECT 11.565 59.925 11.895 60.305 ;
        RECT 12.075 60.095 12.245 60.475 ;
        RECT 13.025 59.925 13.235 60.745 ;
        RECT 13.405 60.725 13.655 61.325 ;
        RECT 13.825 60.915 14.155 61.165 ;
        RECT 13.405 60.095 13.735 60.725 ;
        RECT 13.905 59.925 14.135 60.745 ;
        RECT 14.350 60.665 14.520 61.335 ;
        RECT 15.195 61.165 15.365 62.135 ;
        RECT 14.690 60.835 14.945 61.165 ;
        RECT 15.170 60.835 15.365 61.165 ;
        RECT 15.535 61.795 16.660 61.965 ;
        RECT 14.775 60.665 14.945 60.835 ;
        RECT 15.535 60.665 15.705 61.795 ;
        RECT 14.350 60.095 14.605 60.665 ;
        RECT 14.775 60.495 15.705 60.665 ;
        RECT 15.875 61.455 16.885 61.625 ;
        RECT 15.875 60.655 16.045 61.455 ;
        RECT 15.530 60.460 15.705 60.495 ;
        RECT 14.775 59.925 15.105 60.325 ;
        RECT 15.530 60.095 16.060 60.460 ;
        RECT 16.250 60.435 16.525 61.255 ;
        RECT 16.245 60.265 16.525 60.435 ;
        RECT 16.250 60.095 16.525 60.265 ;
        RECT 16.695 60.095 16.885 61.455 ;
        RECT 17.055 61.470 17.225 62.135 ;
        RECT 17.395 61.715 17.565 62.475 ;
        RECT 17.800 61.715 18.315 62.125 ;
        RECT 17.055 61.280 17.805 61.470 ;
        RECT 17.975 60.905 18.315 61.715 ;
        RECT 18.485 61.310 18.775 62.475 ;
        RECT 18.950 61.335 19.285 62.305 ;
        RECT 19.455 61.335 19.625 62.475 ;
        RECT 19.795 62.135 21.825 62.305 ;
        RECT 17.085 60.735 18.315 60.905 ;
        RECT 17.065 59.925 17.575 60.460 ;
        RECT 17.795 60.130 18.040 60.735 ;
        RECT 18.950 60.665 19.120 61.335 ;
        RECT 19.795 61.165 19.965 62.135 ;
        RECT 19.290 60.835 19.545 61.165 ;
        RECT 19.770 60.835 19.965 61.165 ;
        RECT 20.135 61.795 21.260 61.965 ;
        RECT 19.375 60.665 19.545 60.835 ;
        RECT 20.135 60.665 20.305 61.795 ;
        RECT 18.485 59.925 18.775 60.650 ;
        RECT 18.950 60.095 19.205 60.665 ;
        RECT 19.375 60.495 20.305 60.665 ;
        RECT 20.475 61.455 21.485 61.625 ;
        RECT 20.475 60.655 20.645 61.455 ;
        RECT 20.850 61.115 21.125 61.255 ;
        RECT 20.845 60.945 21.125 61.115 ;
        RECT 20.130 60.460 20.305 60.495 ;
        RECT 19.375 59.925 19.705 60.325 ;
        RECT 20.130 60.095 20.660 60.460 ;
        RECT 20.850 60.095 21.125 60.945 ;
        RECT 21.295 60.095 21.485 61.455 ;
        RECT 21.655 61.470 21.825 62.135 ;
        RECT 21.995 61.715 22.165 62.475 ;
        RECT 22.400 61.715 22.915 62.125 ;
        RECT 21.655 61.280 22.405 61.470 ;
        RECT 22.575 60.905 22.915 61.715 ;
        RECT 21.685 60.735 22.915 60.905 ;
        RECT 23.085 61.335 23.470 62.305 ;
        RECT 23.640 62.015 23.965 62.475 ;
        RECT 24.485 61.845 24.765 62.305 ;
        RECT 23.640 61.625 24.765 61.845 ;
        RECT 21.665 59.925 22.175 60.460 ;
        RECT 22.395 60.130 22.640 60.735 ;
        RECT 23.085 60.665 23.365 61.335 ;
        RECT 23.640 61.165 24.090 61.625 ;
        RECT 24.955 61.455 25.355 62.305 ;
        RECT 25.755 62.015 26.025 62.475 ;
        RECT 26.195 61.845 26.480 62.305 ;
        RECT 23.535 60.835 24.090 61.165 ;
        RECT 24.260 60.895 25.355 61.455 ;
        RECT 23.640 60.725 24.090 60.835 ;
        RECT 23.085 60.095 23.470 60.665 ;
        RECT 23.640 60.555 24.765 60.725 ;
        RECT 23.640 59.925 23.965 60.385 ;
        RECT 24.485 60.095 24.765 60.555 ;
        RECT 24.955 60.095 25.355 60.895 ;
        RECT 25.525 61.625 26.480 61.845 ;
        RECT 25.525 60.725 25.735 61.625 ;
        RECT 25.905 60.895 26.595 61.455 ;
        RECT 27.225 61.335 27.610 62.305 ;
        RECT 27.780 62.015 28.105 62.475 ;
        RECT 28.625 61.845 28.905 62.305 ;
        RECT 27.780 61.625 28.905 61.845 ;
        RECT 25.525 60.555 26.480 60.725 ;
        RECT 25.755 59.925 26.025 60.385 ;
        RECT 26.195 60.095 26.480 60.555 ;
        RECT 27.225 60.665 27.505 61.335 ;
        RECT 27.780 61.165 28.230 61.625 ;
        RECT 29.095 61.455 29.495 62.305 ;
        RECT 29.895 62.015 30.165 62.475 ;
        RECT 30.335 61.845 30.620 62.305 ;
        RECT 27.675 60.835 28.230 61.165 ;
        RECT 28.400 60.895 29.495 61.455 ;
        RECT 27.780 60.725 28.230 60.835 ;
        RECT 27.225 60.095 27.610 60.665 ;
        RECT 27.780 60.555 28.905 60.725 ;
        RECT 27.780 59.925 28.105 60.385 ;
        RECT 28.625 60.095 28.905 60.555 ;
        RECT 29.095 60.095 29.495 60.895 ;
        RECT 29.665 61.625 30.620 61.845 ;
        RECT 29.665 60.725 29.875 61.625 ;
        RECT 30.045 60.895 30.735 61.455 ;
        RECT 30.950 61.335 31.245 62.475 ;
        RECT 31.505 61.505 31.835 62.305 ;
        RECT 32.005 61.675 32.175 62.475 ;
        RECT 32.345 61.505 32.675 62.305 ;
        RECT 32.845 61.675 33.015 62.475 ;
        RECT 33.185 61.525 33.515 62.305 ;
        RECT 33.685 62.015 33.855 62.475 ;
        RECT 34.215 61.805 34.385 62.305 ;
        RECT 34.555 61.975 34.885 62.475 ;
        RECT 34.215 61.635 34.880 61.805 ;
        RECT 33.185 61.505 33.955 61.525 ;
        RECT 31.505 61.335 33.955 61.505 ;
        RECT 30.925 60.915 33.435 61.165 ;
        RECT 33.605 60.745 33.955 61.335 ;
        RECT 34.130 60.815 34.480 61.465 ;
        RECT 29.665 60.555 30.620 60.725 ;
        RECT 29.895 59.925 30.165 60.385 ;
        RECT 30.335 60.095 30.620 60.555 ;
        RECT 31.585 60.565 33.955 60.745 ;
        RECT 34.650 60.645 34.880 61.635 ;
        RECT 30.950 59.925 31.215 60.385 ;
        RECT 31.585 60.095 31.755 60.565 ;
        RECT 32.005 59.925 32.175 60.385 ;
        RECT 32.425 60.095 32.595 60.565 ;
        RECT 32.845 59.925 33.015 60.385 ;
        RECT 33.265 60.095 33.435 60.565 ;
        RECT 34.215 60.475 34.880 60.645 ;
        RECT 33.605 59.925 33.855 60.390 ;
        RECT 34.215 60.185 34.385 60.475 ;
        RECT 34.555 59.925 34.885 60.305 ;
        RECT 35.055 60.185 35.280 62.305 ;
        RECT 35.495 61.975 35.825 62.475 ;
        RECT 35.995 61.805 36.165 62.305 ;
        RECT 36.400 62.090 37.230 62.260 ;
        RECT 37.470 62.095 37.850 62.475 ;
        RECT 35.470 61.635 36.165 61.805 ;
        RECT 35.470 60.665 35.640 61.635 ;
        RECT 35.810 60.845 36.220 61.465 ;
        RECT 36.390 61.415 36.890 61.795 ;
        RECT 35.470 60.475 36.165 60.665 ;
        RECT 36.390 60.545 36.610 61.415 ;
        RECT 37.060 61.245 37.230 62.090 ;
        RECT 38.030 61.925 38.200 62.215 ;
        RECT 38.370 62.095 38.700 62.475 ;
        RECT 39.170 62.005 39.800 62.255 ;
        RECT 39.980 62.095 40.400 62.475 ;
        RECT 39.630 61.925 39.800 62.005 ;
        RECT 40.600 61.925 40.840 62.215 ;
        RECT 37.400 61.675 38.770 61.925 ;
        RECT 37.400 61.415 37.650 61.675 ;
        RECT 38.160 61.245 38.410 61.405 ;
        RECT 37.060 61.075 38.410 61.245 ;
        RECT 37.060 61.035 37.480 61.075 ;
        RECT 36.790 60.485 37.140 60.855 ;
        RECT 35.495 59.925 35.825 60.305 ;
        RECT 35.995 60.145 36.165 60.475 ;
        RECT 37.310 60.305 37.480 61.035 ;
        RECT 38.580 60.905 38.770 61.675 ;
        RECT 37.650 60.575 38.060 60.905 ;
        RECT 38.350 60.565 38.770 60.905 ;
        RECT 38.940 61.495 39.460 61.805 ;
        RECT 39.630 61.755 40.840 61.925 ;
        RECT 41.070 61.785 41.400 62.475 ;
        RECT 38.940 60.735 39.110 61.495 ;
        RECT 39.280 60.905 39.460 61.315 ;
        RECT 39.630 61.245 39.800 61.755 ;
        RECT 41.570 61.605 41.740 62.215 ;
        RECT 42.010 61.755 42.340 62.265 ;
        RECT 41.570 61.585 41.890 61.605 ;
        RECT 39.970 61.415 41.890 61.585 ;
        RECT 39.630 61.075 41.530 61.245 ;
        RECT 39.860 60.735 40.190 60.855 ;
        RECT 38.940 60.565 40.190 60.735 ;
        RECT 36.465 60.105 37.480 60.305 ;
        RECT 37.650 59.925 38.060 60.365 ;
        RECT 38.350 60.135 38.600 60.565 ;
        RECT 38.800 59.925 39.120 60.385 ;
        RECT 40.360 60.315 40.530 61.075 ;
        RECT 41.200 61.015 41.530 61.075 ;
        RECT 40.720 60.845 41.050 60.905 ;
        RECT 40.720 60.575 41.380 60.845 ;
        RECT 41.700 60.520 41.890 61.415 ;
        RECT 39.680 60.145 40.530 60.315 ;
        RECT 40.730 59.925 41.390 60.405 ;
        RECT 41.570 60.190 41.890 60.520 ;
        RECT 42.090 61.165 42.340 61.755 ;
        RECT 42.520 61.675 42.805 62.475 ;
        RECT 42.985 61.495 43.240 62.165 ;
        RECT 42.090 60.835 42.890 61.165 ;
        RECT 42.090 60.185 42.340 60.835 ;
        RECT 43.060 60.635 43.240 61.495 ;
        RECT 44.245 61.310 44.535 62.475 ;
        RECT 45.625 61.400 45.895 62.305 ;
        RECT 46.065 61.715 46.395 62.475 ;
        RECT 46.575 61.545 46.745 62.305 ;
        RECT 42.985 60.435 43.240 60.635 ;
        RECT 42.520 59.925 42.805 60.385 ;
        RECT 42.985 60.265 43.325 60.435 ;
        RECT 42.985 60.105 43.240 60.265 ;
        RECT 44.245 59.925 44.535 60.650 ;
        RECT 45.625 60.600 45.795 61.400 ;
        RECT 46.080 61.375 46.745 61.545 ;
        RECT 46.080 61.230 46.250 61.375 ;
        RECT 45.965 60.900 46.250 61.230 ;
        RECT 47.010 61.335 47.345 62.305 ;
        RECT 47.515 61.335 47.685 62.475 ;
        RECT 47.855 62.135 49.885 62.305 ;
        RECT 46.080 60.645 46.250 60.900 ;
        RECT 46.485 60.825 46.815 61.195 ;
        RECT 47.010 60.665 47.180 61.335 ;
        RECT 47.855 61.165 48.025 62.135 ;
        RECT 47.350 60.835 47.605 61.165 ;
        RECT 47.830 60.835 48.025 61.165 ;
        RECT 48.195 61.795 49.320 61.965 ;
        RECT 47.435 60.665 47.605 60.835 ;
        RECT 48.195 60.665 48.365 61.795 ;
        RECT 45.625 60.095 45.885 60.600 ;
        RECT 46.080 60.475 46.745 60.645 ;
        RECT 46.065 59.925 46.395 60.305 ;
        RECT 46.575 60.095 46.745 60.475 ;
        RECT 47.010 60.095 47.265 60.665 ;
        RECT 47.435 60.495 48.365 60.665 ;
        RECT 48.535 61.455 49.545 61.625 ;
        RECT 48.535 60.655 48.705 61.455 ;
        RECT 48.910 60.775 49.185 61.255 ;
        RECT 48.905 60.605 49.185 60.775 ;
        RECT 48.190 60.460 48.365 60.495 ;
        RECT 47.435 59.925 47.765 60.325 ;
        RECT 48.190 60.095 48.720 60.460 ;
        RECT 48.910 60.095 49.185 60.605 ;
        RECT 49.355 60.095 49.545 61.455 ;
        RECT 49.715 61.470 49.885 62.135 ;
        RECT 50.055 61.715 50.225 62.475 ;
        RECT 50.460 61.715 50.975 62.125 ;
        RECT 49.715 61.280 50.465 61.470 ;
        RECT 50.635 60.905 50.975 61.715 ;
        RECT 51.185 61.335 51.415 62.475 ;
        RECT 51.585 61.325 51.915 62.305 ;
        RECT 52.085 61.335 52.295 62.475 ;
        RECT 52.525 62.040 57.870 62.475 ;
        RECT 51.165 60.915 51.495 61.165 ;
        RECT 49.745 60.735 50.975 60.905 ;
        RECT 49.725 59.925 50.235 60.460 ;
        RECT 50.455 60.130 50.700 60.735 ;
        RECT 51.185 59.925 51.415 60.745 ;
        RECT 51.665 60.725 51.915 61.325 ;
        RECT 51.585 60.095 51.915 60.725 ;
        RECT 52.085 59.925 52.295 60.745 ;
        RECT 54.110 60.470 54.450 61.300 ;
        RECT 55.930 60.790 56.280 62.040 ;
        RECT 58.045 61.385 60.635 62.475 ;
        RECT 58.045 60.695 59.255 61.215 ;
        RECT 59.425 60.865 60.635 61.385 ;
        RECT 61.270 61.325 61.530 62.475 ;
        RECT 61.705 61.400 61.960 62.305 ;
        RECT 62.130 61.715 62.460 62.475 ;
        RECT 62.675 61.545 62.845 62.305 ;
        RECT 52.525 59.925 57.870 60.470 ;
        RECT 58.045 59.925 60.635 60.695 ;
        RECT 61.270 59.925 61.530 60.765 ;
        RECT 61.705 60.670 61.875 61.400 ;
        RECT 62.130 61.375 62.845 61.545 ;
        RECT 62.130 61.165 62.300 61.375 ;
        RECT 63.110 61.325 63.370 62.475 ;
        RECT 63.545 61.400 63.800 62.305 ;
        RECT 63.970 61.715 64.300 62.475 ;
        RECT 64.515 61.545 64.685 62.305 ;
        RECT 62.045 60.835 62.300 61.165 ;
        RECT 61.705 60.095 61.960 60.670 ;
        RECT 62.130 60.645 62.300 60.835 ;
        RECT 62.580 60.825 62.935 61.195 ;
        RECT 62.130 60.475 62.845 60.645 ;
        RECT 62.130 59.925 62.460 60.305 ;
        RECT 62.675 60.095 62.845 60.475 ;
        RECT 63.110 59.925 63.370 60.765 ;
        RECT 63.545 60.670 63.715 61.400 ;
        RECT 63.970 61.375 64.685 61.545 ;
        RECT 65.035 61.545 65.205 62.305 ;
        RECT 65.420 61.715 65.750 62.475 ;
        RECT 65.035 61.375 65.750 61.545 ;
        RECT 65.920 61.400 66.175 62.305 ;
        RECT 63.970 61.165 64.140 61.375 ;
        RECT 63.885 60.835 64.140 61.165 ;
        RECT 63.545 60.095 63.800 60.670 ;
        RECT 63.970 60.645 64.140 60.835 ;
        RECT 64.420 60.825 64.775 61.195 ;
        RECT 64.945 60.825 65.300 61.195 ;
        RECT 65.580 61.165 65.750 61.375 ;
        RECT 65.580 60.835 65.835 61.165 ;
        RECT 65.580 60.645 65.750 60.835 ;
        RECT 66.005 60.670 66.175 61.400 ;
        RECT 66.350 61.325 66.610 62.475 ;
        RECT 66.875 61.545 67.045 62.305 ;
        RECT 67.260 61.715 67.590 62.475 ;
        RECT 66.875 61.375 67.590 61.545 ;
        RECT 67.760 61.400 68.015 62.305 ;
        RECT 66.785 60.825 67.140 61.195 ;
        RECT 67.420 61.165 67.590 61.375 ;
        RECT 67.420 60.835 67.675 61.165 ;
        RECT 63.970 60.475 64.685 60.645 ;
        RECT 63.970 59.925 64.300 60.305 ;
        RECT 64.515 60.095 64.685 60.475 ;
        RECT 65.035 60.475 65.750 60.645 ;
        RECT 65.035 60.095 65.205 60.475 ;
        RECT 65.420 59.925 65.750 60.305 ;
        RECT 65.920 60.095 66.175 60.670 ;
        RECT 66.350 59.925 66.610 60.765 ;
        RECT 67.420 60.645 67.590 60.835 ;
        RECT 67.845 60.670 68.015 61.400 ;
        RECT 68.190 61.325 68.450 62.475 ;
        RECT 68.625 61.385 69.835 62.475 ;
        RECT 66.875 60.475 67.590 60.645 ;
        RECT 66.875 60.095 67.045 60.475 ;
        RECT 67.260 59.925 67.590 60.305 ;
        RECT 67.760 60.095 68.015 60.670 ;
        RECT 68.190 59.925 68.450 60.765 ;
        RECT 68.625 60.675 69.145 61.215 ;
        RECT 69.315 60.845 69.835 61.385 ;
        RECT 70.005 61.310 70.295 62.475 ;
        RECT 70.465 61.385 72.135 62.475 ;
        RECT 70.465 60.695 71.215 61.215 ;
        RECT 71.385 60.865 72.135 61.385 ;
        RECT 72.305 61.400 72.575 62.305 ;
        RECT 72.745 61.715 73.075 62.475 ;
        RECT 73.255 61.545 73.425 62.305 ;
        RECT 68.625 59.925 69.835 60.675 ;
        RECT 70.005 59.925 70.295 60.650 ;
        RECT 70.465 59.925 72.135 60.695 ;
        RECT 72.305 60.600 72.475 61.400 ;
        RECT 72.760 61.375 73.425 61.545 ;
        RECT 73.685 61.385 75.355 62.475 ;
        RECT 72.760 61.230 72.930 61.375 ;
        RECT 72.645 60.900 72.930 61.230 ;
        RECT 72.760 60.645 72.930 60.900 ;
        RECT 73.165 60.825 73.495 61.195 ;
        RECT 73.685 60.695 74.435 61.215 ;
        RECT 74.605 60.865 75.355 61.385 ;
        RECT 75.990 61.335 76.325 62.305 ;
        RECT 76.495 61.335 76.665 62.475 ;
        RECT 76.835 62.135 78.865 62.305 ;
        RECT 72.305 60.095 72.565 60.600 ;
        RECT 72.760 60.475 73.425 60.645 ;
        RECT 72.745 59.925 73.075 60.305 ;
        RECT 73.255 60.095 73.425 60.475 ;
        RECT 73.685 59.925 75.355 60.695 ;
        RECT 75.990 60.665 76.160 61.335 ;
        RECT 76.835 61.165 77.005 62.135 ;
        RECT 76.330 60.835 76.585 61.165 ;
        RECT 76.810 60.835 77.005 61.165 ;
        RECT 77.175 61.795 78.300 61.965 ;
        RECT 76.415 60.665 76.585 60.835 ;
        RECT 77.175 60.665 77.345 61.795 ;
        RECT 75.990 60.095 76.245 60.665 ;
        RECT 76.415 60.495 77.345 60.665 ;
        RECT 77.515 61.455 78.525 61.625 ;
        RECT 77.515 60.655 77.685 61.455 ;
        RECT 77.170 60.460 77.345 60.495 ;
        RECT 76.415 59.925 76.745 60.325 ;
        RECT 77.170 60.095 77.700 60.460 ;
        RECT 77.890 60.435 78.165 61.255 ;
        RECT 77.885 60.265 78.165 60.435 ;
        RECT 77.890 60.095 78.165 60.265 ;
        RECT 78.335 60.095 78.525 61.455 ;
        RECT 78.695 61.470 78.865 62.135 ;
        RECT 79.035 61.715 79.205 62.475 ;
        RECT 79.440 61.715 79.955 62.125 ;
        RECT 78.695 61.280 79.445 61.470 ;
        RECT 79.615 60.905 79.955 61.715 ;
        RECT 78.725 60.735 79.955 60.905 ;
        RECT 80.125 61.715 80.640 62.125 ;
        RECT 80.875 61.715 81.045 62.475 ;
        RECT 81.215 62.135 83.245 62.305 ;
        RECT 80.125 60.905 80.465 61.715 ;
        RECT 81.215 61.470 81.385 62.135 ;
        RECT 81.780 61.795 82.905 61.965 ;
        RECT 80.635 61.280 81.385 61.470 ;
        RECT 81.555 61.455 82.565 61.625 ;
        RECT 80.125 60.735 81.355 60.905 ;
        RECT 78.705 59.925 79.215 60.460 ;
        RECT 79.435 60.130 79.680 60.735 ;
        RECT 80.400 60.130 80.645 60.735 ;
        RECT 80.865 59.925 81.375 60.460 ;
        RECT 81.555 60.095 81.745 61.455 ;
        RECT 81.915 61.115 82.190 61.255 ;
        RECT 81.915 60.945 82.195 61.115 ;
        RECT 81.915 60.095 82.190 60.945 ;
        RECT 82.395 60.655 82.565 61.455 ;
        RECT 82.735 60.665 82.905 61.795 ;
        RECT 83.075 61.165 83.245 62.135 ;
        RECT 83.415 61.335 83.585 62.475 ;
        RECT 83.755 61.335 84.090 62.305 ;
        RECT 84.355 61.545 84.525 62.305 ;
        RECT 84.705 61.715 85.035 62.475 ;
        RECT 84.355 61.375 85.020 61.545 ;
        RECT 85.205 61.400 85.475 62.305 ;
        RECT 83.075 60.835 83.270 61.165 ;
        RECT 83.495 60.835 83.750 61.165 ;
        RECT 83.495 60.665 83.665 60.835 ;
        RECT 83.920 60.665 84.090 61.335 ;
        RECT 84.850 61.230 85.020 61.375 ;
        RECT 84.285 60.825 84.615 61.195 ;
        RECT 84.850 60.900 85.135 61.230 ;
        RECT 82.735 60.495 83.665 60.665 ;
        RECT 82.735 60.460 82.910 60.495 ;
        RECT 82.380 60.095 82.910 60.460 ;
        RECT 83.335 59.925 83.665 60.325 ;
        RECT 83.835 60.095 84.090 60.665 ;
        RECT 84.850 60.645 85.020 60.900 ;
        RECT 84.355 60.475 85.020 60.645 ;
        RECT 85.305 60.600 85.475 61.400 ;
        RECT 85.645 61.715 86.160 62.125 ;
        RECT 86.395 61.715 86.565 62.475 ;
        RECT 86.735 62.135 88.765 62.305 ;
        RECT 85.645 60.905 85.985 61.715 ;
        RECT 86.735 61.470 86.905 62.135 ;
        RECT 87.300 61.795 88.425 61.965 ;
        RECT 86.155 61.280 86.905 61.470 ;
        RECT 87.075 61.455 88.085 61.625 ;
        RECT 85.645 60.735 86.875 60.905 ;
        RECT 84.355 60.095 84.525 60.475 ;
        RECT 84.705 59.925 85.035 60.305 ;
        RECT 85.215 60.095 85.475 60.600 ;
        RECT 85.920 60.130 86.165 60.735 ;
        RECT 86.385 59.925 86.895 60.460 ;
        RECT 87.075 60.095 87.265 61.455 ;
        RECT 87.435 60.435 87.710 61.255 ;
        RECT 87.915 60.655 88.085 61.455 ;
        RECT 88.255 60.665 88.425 61.795 ;
        RECT 88.595 61.165 88.765 62.135 ;
        RECT 88.935 61.335 89.105 62.475 ;
        RECT 89.275 61.335 89.610 62.305 ;
        RECT 88.595 60.835 88.790 61.165 ;
        RECT 89.015 60.835 89.270 61.165 ;
        RECT 89.015 60.665 89.185 60.835 ;
        RECT 89.440 60.665 89.610 61.335 ;
        RECT 88.255 60.495 89.185 60.665 ;
        RECT 88.255 60.460 88.430 60.495 ;
        RECT 87.435 60.265 87.715 60.435 ;
        RECT 87.435 60.095 87.710 60.265 ;
        RECT 87.900 60.095 88.430 60.460 ;
        RECT 88.855 59.925 89.185 60.325 ;
        RECT 89.355 60.095 89.610 60.665 ;
        RECT 89.785 61.335 90.170 62.305 ;
        RECT 90.340 62.015 90.665 62.475 ;
        RECT 91.185 61.845 91.465 62.305 ;
        RECT 90.340 61.625 91.465 61.845 ;
        RECT 89.785 60.665 90.065 61.335 ;
        RECT 90.340 61.165 90.790 61.625 ;
        RECT 91.655 61.455 92.055 62.305 ;
        RECT 92.455 62.015 92.725 62.475 ;
        RECT 92.895 61.845 93.180 62.305 ;
        RECT 90.235 60.835 90.790 61.165 ;
        RECT 90.960 60.895 92.055 61.455 ;
        RECT 90.340 60.725 90.790 60.835 ;
        RECT 89.785 60.095 90.170 60.665 ;
        RECT 90.340 60.555 91.465 60.725 ;
        RECT 90.340 59.925 90.665 60.385 ;
        RECT 91.185 60.095 91.465 60.555 ;
        RECT 91.655 60.095 92.055 60.895 ;
        RECT 92.225 61.625 93.180 61.845 ;
        RECT 92.225 60.725 92.435 61.625 ;
        RECT 92.605 60.895 93.295 61.455 ;
        RECT 93.465 61.385 95.135 62.475 ;
        RECT 92.225 60.555 93.180 60.725 ;
        RECT 92.455 59.925 92.725 60.385 ;
        RECT 92.895 60.095 93.180 60.555 ;
        RECT 93.465 60.695 94.215 61.215 ;
        RECT 94.385 60.865 95.135 61.385 ;
        RECT 95.765 61.310 96.055 62.475 ;
        RECT 96.225 61.715 96.740 62.125 ;
        RECT 96.975 61.715 97.145 62.475 ;
        RECT 97.315 62.135 99.345 62.305 ;
        RECT 96.225 60.905 96.565 61.715 ;
        RECT 97.315 61.470 97.485 62.135 ;
        RECT 97.880 61.795 99.005 61.965 ;
        RECT 96.735 61.280 97.485 61.470 ;
        RECT 97.655 61.455 98.665 61.625 ;
        RECT 96.225 60.735 97.455 60.905 ;
        RECT 93.465 59.925 95.135 60.695 ;
        RECT 95.765 59.925 96.055 60.650 ;
        RECT 96.500 60.130 96.745 60.735 ;
        RECT 96.965 59.925 97.475 60.460 ;
        RECT 97.655 60.095 97.845 61.455 ;
        RECT 98.015 60.775 98.290 61.255 ;
        RECT 98.015 60.605 98.295 60.775 ;
        RECT 98.495 60.655 98.665 61.455 ;
        RECT 98.835 60.665 99.005 61.795 ;
        RECT 99.175 61.165 99.345 62.135 ;
        RECT 99.515 61.335 99.685 62.475 ;
        RECT 99.855 61.335 100.190 62.305 ;
        RECT 100.365 61.385 101.575 62.475 ;
        RECT 99.175 60.835 99.370 61.165 ;
        RECT 99.595 60.835 99.850 61.165 ;
        RECT 99.595 60.665 99.765 60.835 ;
        RECT 100.020 60.665 100.190 61.335 ;
        RECT 98.015 60.095 98.290 60.605 ;
        RECT 98.835 60.495 99.765 60.665 ;
        RECT 98.835 60.460 99.010 60.495 ;
        RECT 98.480 60.095 99.010 60.460 ;
        RECT 99.435 59.925 99.765 60.325 ;
        RECT 99.935 60.095 100.190 60.665 ;
        RECT 100.365 60.675 100.885 61.215 ;
        RECT 101.055 60.845 101.575 61.385 ;
        RECT 101.745 61.715 102.260 62.125 ;
        RECT 102.495 61.715 102.665 62.475 ;
        RECT 102.835 62.135 104.865 62.305 ;
        RECT 101.745 60.905 102.085 61.715 ;
        RECT 102.835 61.470 103.005 62.135 ;
        RECT 103.400 61.795 104.525 61.965 ;
        RECT 102.255 61.280 103.005 61.470 ;
        RECT 103.175 61.455 104.185 61.625 ;
        RECT 101.745 60.735 102.975 60.905 ;
        RECT 100.365 59.925 101.575 60.675 ;
        RECT 102.020 60.130 102.265 60.735 ;
        RECT 102.485 59.925 102.995 60.460 ;
        RECT 103.175 60.095 103.365 61.455 ;
        RECT 103.535 60.775 103.810 61.255 ;
        RECT 103.535 60.605 103.815 60.775 ;
        RECT 104.015 60.655 104.185 61.455 ;
        RECT 104.355 60.665 104.525 61.795 ;
        RECT 104.695 61.165 104.865 62.135 ;
        RECT 105.035 61.335 105.205 62.475 ;
        RECT 105.375 61.335 105.710 62.305 ;
        RECT 105.975 61.805 106.145 62.305 ;
        RECT 106.315 61.975 106.645 62.475 ;
        RECT 105.975 61.635 106.640 61.805 ;
        RECT 104.695 60.835 104.890 61.165 ;
        RECT 105.115 60.835 105.370 61.165 ;
        RECT 105.115 60.665 105.285 60.835 ;
        RECT 105.540 60.665 105.710 61.335 ;
        RECT 105.890 60.815 106.240 61.465 ;
        RECT 103.535 60.095 103.810 60.605 ;
        RECT 104.355 60.495 105.285 60.665 ;
        RECT 104.355 60.460 104.530 60.495 ;
        RECT 104.000 60.095 104.530 60.460 ;
        RECT 104.955 59.925 105.285 60.325 ;
        RECT 105.455 60.095 105.710 60.665 ;
        RECT 106.410 60.645 106.640 61.635 ;
        RECT 105.975 60.475 106.640 60.645 ;
        RECT 105.975 60.185 106.145 60.475 ;
        RECT 106.315 59.925 106.645 60.305 ;
        RECT 106.815 60.185 107.040 62.305 ;
        RECT 107.255 61.975 107.585 62.475 ;
        RECT 107.755 61.805 107.925 62.305 ;
        RECT 108.160 62.090 108.990 62.260 ;
        RECT 109.230 62.095 109.610 62.475 ;
        RECT 107.230 61.635 107.925 61.805 ;
        RECT 107.230 60.665 107.400 61.635 ;
        RECT 107.570 60.845 107.980 61.465 ;
        RECT 108.150 61.415 108.650 61.795 ;
        RECT 107.230 60.475 107.925 60.665 ;
        RECT 108.150 60.545 108.370 61.415 ;
        RECT 108.820 61.245 108.990 62.090 ;
        RECT 109.790 61.925 109.960 62.215 ;
        RECT 110.130 62.095 110.460 62.475 ;
        RECT 110.930 62.005 111.560 62.255 ;
        RECT 111.740 62.095 112.160 62.475 ;
        RECT 111.390 61.925 111.560 62.005 ;
        RECT 112.360 61.925 112.600 62.215 ;
        RECT 109.160 61.675 110.530 61.925 ;
        RECT 109.160 61.415 109.410 61.675 ;
        RECT 109.920 61.245 110.170 61.405 ;
        RECT 108.820 61.075 110.170 61.245 ;
        RECT 108.820 61.035 109.240 61.075 ;
        RECT 108.550 60.485 108.900 60.855 ;
        RECT 107.255 59.925 107.585 60.305 ;
        RECT 107.755 60.145 107.925 60.475 ;
        RECT 109.070 60.305 109.240 61.035 ;
        RECT 110.340 60.905 110.530 61.675 ;
        RECT 109.410 60.575 109.820 60.905 ;
        RECT 110.110 60.565 110.530 60.905 ;
        RECT 110.700 61.495 111.220 61.805 ;
        RECT 111.390 61.755 112.600 61.925 ;
        RECT 112.830 61.785 113.160 62.475 ;
        RECT 110.700 60.735 110.870 61.495 ;
        RECT 111.040 60.905 111.220 61.315 ;
        RECT 111.390 61.245 111.560 61.755 ;
        RECT 113.330 61.605 113.500 62.215 ;
        RECT 113.770 61.755 114.100 62.265 ;
        RECT 113.330 61.585 113.650 61.605 ;
        RECT 111.730 61.415 113.650 61.585 ;
        RECT 111.390 61.075 113.290 61.245 ;
        RECT 111.620 60.735 111.950 60.855 ;
        RECT 110.700 60.565 111.950 60.735 ;
        RECT 108.225 60.105 109.240 60.305 ;
        RECT 109.410 59.925 109.820 60.365 ;
        RECT 110.110 60.135 110.360 60.565 ;
        RECT 110.560 59.925 110.880 60.385 ;
        RECT 112.120 60.315 112.290 61.075 ;
        RECT 112.960 61.015 113.290 61.075 ;
        RECT 112.480 60.845 112.810 60.905 ;
        RECT 112.480 60.575 113.140 60.845 ;
        RECT 113.460 60.520 113.650 61.415 ;
        RECT 111.440 60.145 112.290 60.315 ;
        RECT 112.490 59.925 113.150 60.405 ;
        RECT 113.330 60.190 113.650 60.520 ;
        RECT 113.850 61.165 114.100 61.755 ;
        RECT 114.280 61.675 114.565 62.475 ;
        RECT 114.745 62.135 115.000 62.165 ;
        RECT 114.745 61.965 115.085 62.135 ;
        RECT 114.745 61.495 115.000 61.965 ;
        RECT 113.850 60.835 114.650 61.165 ;
        RECT 113.850 60.185 114.100 60.835 ;
        RECT 114.820 60.635 115.000 61.495 ;
        RECT 115.545 61.385 117.215 62.475 ;
        RECT 114.280 59.925 114.565 60.385 ;
        RECT 114.745 60.105 115.000 60.635 ;
        RECT 115.545 60.695 116.295 61.215 ;
        RECT 116.465 60.865 117.215 61.385 ;
        RECT 117.385 61.385 118.595 62.475 ;
        RECT 117.385 60.845 117.905 61.385 ;
        RECT 115.545 59.925 117.215 60.695 ;
        RECT 118.075 60.675 118.595 61.215 ;
        RECT 117.385 59.925 118.595 60.675 ;
        RECT 5.520 59.755 118.680 59.925 ;
        RECT 5.605 59.005 6.815 59.755 ;
        RECT 5.605 58.465 6.125 59.005 ;
        RECT 6.985 58.985 8.655 59.755 ;
        RECT 9.375 59.205 9.545 59.585 ;
        RECT 9.725 59.375 10.055 59.755 ;
        RECT 9.375 59.035 10.040 59.205 ;
        RECT 10.235 59.080 10.495 59.585 ;
        RECT 6.295 58.295 6.815 58.835 ;
        RECT 6.985 58.465 7.735 58.985 ;
        RECT 7.905 58.295 8.655 58.815 ;
        RECT 9.305 58.485 9.635 58.855 ;
        RECT 9.870 58.780 10.040 59.035 ;
        RECT 9.870 58.450 10.155 58.780 ;
        RECT 9.870 58.305 10.040 58.450 ;
        RECT 5.605 57.205 6.815 58.295 ;
        RECT 6.985 57.205 8.655 58.295 ;
        RECT 9.375 58.135 10.040 58.305 ;
        RECT 10.325 58.280 10.495 59.080 ;
        RECT 10.670 59.205 10.925 59.495 ;
        RECT 11.095 59.375 11.425 59.755 ;
        RECT 10.670 59.035 11.420 59.205 ;
        RECT 9.375 57.375 9.545 58.135 ;
        RECT 9.725 57.205 10.055 57.965 ;
        RECT 10.225 57.375 10.495 58.280 ;
        RECT 10.670 58.215 11.020 58.865 ;
        RECT 11.190 58.045 11.420 59.035 ;
        RECT 10.670 57.875 11.420 58.045 ;
        RECT 10.670 57.375 10.925 57.875 ;
        RECT 11.095 57.205 11.425 57.705 ;
        RECT 11.595 57.375 11.765 59.495 ;
        RECT 12.125 59.395 12.455 59.755 ;
        RECT 12.625 59.365 13.120 59.535 ;
        RECT 13.325 59.365 14.180 59.535 ;
        RECT 11.995 58.175 12.455 59.225 ;
        RECT 11.935 57.390 12.260 58.175 ;
        RECT 12.625 58.005 12.795 59.365 ;
        RECT 12.965 58.455 13.315 59.075 ;
        RECT 13.485 58.855 13.840 59.075 ;
        RECT 13.485 58.265 13.655 58.855 ;
        RECT 14.010 58.655 14.180 59.365 ;
        RECT 15.055 59.295 15.385 59.755 ;
        RECT 15.595 59.395 15.945 59.565 ;
        RECT 14.385 58.825 15.175 59.075 ;
        RECT 15.595 59.005 15.855 59.395 ;
        RECT 16.165 59.305 17.115 59.585 ;
        RECT 17.285 59.315 17.475 59.755 ;
        RECT 17.645 59.375 18.715 59.545 ;
        RECT 15.345 58.655 15.515 58.835 ;
        RECT 12.625 57.835 13.020 58.005 ;
        RECT 13.190 57.875 13.655 58.265 ;
        RECT 13.825 58.485 15.515 58.655 ;
        RECT 12.850 57.705 13.020 57.835 ;
        RECT 13.825 57.705 13.995 58.485 ;
        RECT 15.685 58.315 15.855 59.005 ;
        RECT 14.355 58.145 15.855 58.315 ;
        RECT 16.045 58.345 16.255 59.135 ;
        RECT 16.425 58.515 16.775 59.135 ;
        RECT 16.945 58.525 17.115 59.305 ;
        RECT 17.645 59.145 17.815 59.375 ;
        RECT 17.285 58.975 17.815 59.145 ;
        RECT 17.285 58.695 17.505 58.975 ;
        RECT 17.985 58.805 18.225 59.205 ;
        RECT 16.945 58.355 17.350 58.525 ;
        RECT 17.685 58.435 18.225 58.805 ;
        RECT 18.395 59.020 18.715 59.375 ;
        RECT 18.960 59.295 19.265 59.755 ;
        RECT 19.435 59.045 19.690 59.575 ;
        RECT 18.395 58.845 18.720 59.020 ;
        RECT 18.395 58.545 19.310 58.845 ;
        RECT 18.570 58.515 19.310 58.545 ;
        RECT 16.045 58.185 16.720 58.345 ;
        RECT 17.180 58.265 17.350 58.355 ;
        RECT 16.045 58.175 17.010 58.185 ;
        RECT 15.685 58.005 15.855 58.145 ;
        RECT 12.430 57.205 12.680 57.665 ;
        RECT 12.850 57.375 13.100 57.705 ;
        RECT 13.315 57.375 13.995 57.705 ;
        RECT 14.165 57.805 15.240 57.975 ;
        RECT 15.685 57.835 16.245 58.005 ;
        RECT 16.550 57.885 17.010 58.175 ;
        RECT 17.180 58.095 18.400 58.265 ;
        RECT 14.165 57.465 14.335 57.805 ;
        RECT 14.570 57.205 14.900 57.635 ;
        RECT 15.070 57.465 15.240 57.805 ;
        RECT 15.535 57.205 15.905 57.665 ;
        RECT 16.075 57.375 16.245 57.835 ;
        RECT 17.180 57.715 17.350 58.095 ;
        RECT 18.570 57.925 18.740 58.515 ;
        RECT 19.480 58.395 19.690 59.045 ;
        RECT 19.955 59.105 20.125 59.585 ;
        RECT 20.305 59.275 20.545 59.755 ;
        RECT 20.795 59.105 20.965 59.585 ;
        RECT 21.135 59.275 21.465 59.755 ;
        RECT 21.635 59.105 21.805 59.585 ;
        RECT 19.955 58.935 20.590 59.105 ;
        RECT 20.795 58.935 21.805 59.105 ;
        RECT 21.975 58.955 22.305 59.755 ;
        RECT 22.900 58.945 23.145 59.550 ;
        RECT 23.365 59.220 23.875 59.755 ;
        RECT 20.420 58.765 20.590 58.935 ;
        RECT 21.305 58.905 21.805 58.935 ;
        RECT 19.870 58.525 20.250 58.765 ;
        RECT 20.420 58.595 20.920 58.765 ;
        RECT 16.480 57.375 17.350 57.715 ;
        RECT 17.940 57.755 18.740 57.925 ;
        RECT 17.520 57.205 17.770 57.665 ;
        RECT 17.940 57.465 18.110 57.755 ;
        RECT 18.290 57.205 18.620 57.585 ;
        RECT 18.960 57.205 19.265 58.345 ;
        RECT 19.435 57.515 19.690 58.395 ;
        RECT 20.420 58.355 20.590 58.595 ;
        RECT 21.310 58.395 21.805 58.905 ;
        RECT 19.875 58.185 20.590 58.355 ;
        RECT 20.795 58.225 21.805 58.395 ;
        RECT 22.625 58.775 23.855 58.945 ;
        RECT 19.875 57.375 20.205 58.185 ;
        RECT 20.375 57.205 20.615 58.005 ;
        RECT 20.795 57.375 20.965 58.225 ;
        RECT 21.135 57.205 21.465 58.005 ;
        RECT 21.635 57.375 21.805 58.225 ;
        RECT 21.975 57.205 22.305 58.355 ;
        RECT 22.625 57.965 22.965 58.775 ;
        RECT 23.135 58.210 23.885 58.400 ;
        RECT 22.625 57.555 23.140 57.965 ;
        RECT 23.375 57.205 23.545 57.965 ;
        RECT 23.715 57.545 23.885 58.210 ;
        RECT 24.055 58.225 24.245 59.585 ;
        RECT 24.415 59.415 24.690 59.585 ;
        RECT 24.415 59.245 24.695 59.415 ;
        RECT 24.415 58.425 24.690 59.245 ;
        RECT 24.880 59.220 25.410 59.585 ;
        RECT 25.835 59.355 26.165 59.755 ;
        RECT 25.235 59.185 25.410 59.220 ;
        RECT 24.895 58.225 25.065 59.025 ;
        RECT 24.055 58.055 25.065 58.225 ;
        RECT 25.235 59.015 26.165 59.185 ;
        RECT 26.335 59.015 26.590 59.585 ;
        RECT 25.235 57.885 25.405 59.015 ;
        RECT 25.995 58.845 26.165 59.015 ;
        RECT 24.280 57.715 25.405 57.885 ;
        RECT 25.575 58.515 25.770 58.845 ;
        RECT 25.995 58.515 26.250 58.845 ;
        RECT 25.575 57.545 25.745 58.515 ;
        RECT 26.420 58.345 26.590 59.015 ;
        RECT 23.715 57.375 25.745 57.545 ;
        RECT 25.915 57.205 26.085 58.345 ;
        RECT 26.255 57.375 26.590 58.345 ;
        RECT 27.230 59.015 27.485 59.585 ;
        RECT 27.655 59.355 27.985 59.755 ;
        RECT 28.410 59.220 28.940 59.585 ;
        RECT 28.410 59.185 28.585 59.220 ;
        RECT 27.655 59.015 28.585 59.185 ;
        RECT 29.130 59.075 29.405 59.585 ;
        RECT 27.230 58.345 27.400 59.015 ;
        RECT 27.655 58.845 27.825 59.015 ;
        RECT 27.570 58.515 27.825 58.845 ;
        RECT 28.050 58.515 28.245 58.845 ;
        RECT 27.230 57.375 27.565 58.345 ;
        RECT 27.735 57.205 27.905 58.345 ;
        RECT 28.075 57.545 28.245 58.515 ;
        RECT 28.415 57.885 28.585 59.015 ;
        RECT 28.755 58.225 28.925 59.025 ;
        RECT 29.125 58.905 29.405 59.075 ;
        RECT 29.130 58.425 29.405 58.905 ;
        RECT 29.575 58.225 29.765 59.585 ;
        RECT 29.945 59.220 30.455 59.755 ;
        RECT 30.675 58.945 30.920 59.550 ;
        RECT 31.365 59.030 31.655 59.755 ;
        RECT 31.825 59.245 32.130 59.755 ;
        RECT 29.965 58.775 31.195 58.945 ;
        RECT 28.755 58.055 29.765 58.225 ;
        RECT 29.935 58.210 30.685 58.400 ;
        RECT 28.415 57.715 29.540 57.885 ;
        RECT 29.935 57.545 30.105 58.210 ;
        RECT 30.855 57.965 31.195 58.775 ;
        RECT 31.825 58.515 32.140 59.075 ;
        RECT 32.310 58.765 32.560 59.575 ;
        RECT 32.730 59.230 32.990 59.755 ;
        RECT 33.170 58.765 33.420 59.575 ;
        RECT 33.590 59.195 33.850 59.755 ;
        RECT 34.020 59.105 34.280 59.560 ;
        RECT 34.450 59.275 34.710 59.755 ;
        RECT 34.880 59.105 35.140 59.560 ;
        RECT 35.310 59.275 35.570 59.755 ;
        RECT 35.740 59.105 36.000 59.560 ;
        RECT 36.170 59.275 36.415 59.755 ;
        RECT 36.585 59.105 36.860 59.560 ;
        RECT 37.030 59.275 37.275 59.755 ;
        RECT 37.445 59.105 37.705 59.560 ;
        RECT 37.885 59.275 38.135 59.755 ;
        RECT 38.305 59.105 38.565 59.560 ;
        RECT 38.745 59.275 38.995 59.755 ;
        RECT 39.165 59.105 39.425 59.560 ;
        RECT 39.605 59.275 39.865 59.755 ;
        RECT 40.035 59.105 40.295 59.560 ;
        RECT 40.465 59.275 40.765 59.755 ;
        RECT 41.025 59.210 46.370 59.755 ;
        RECT 34.020 58.935 40.765 59.105 ;
        RECT 32.310 58.515 39.430 58.765 ;
        RECT 28.075 57.375 30.105 57.545 ;
        RECT 30.275 57.205 30.445 57.965 ;
        RECT 30.680 57.555 31.195 57.965 ;
        RECT 31.365 57.205 31.655 58.370 ;
        RECT 31.835 57.205 32.130 58.015 ;
        RECT 32.310 57.375 32.555 58.515 ;
        RECT 32.730 57.205 32.990 58.015 ;
        RECT 33.170 57.380 33.420 58.515 ;
        RECT 39.600 58.345 40.765 58.935 ;
        RECT 42.610 58.380 42.950 59.210 ;
        RECT 46.545 59.080 46.805 59.585 ;
        RECT 46.985 59.375 47.315 59.755 ;
        RECT 47.495 59.205 47.665 59.585 ;
        RECT 34.020 58.120 40.765 58.345 ;
        RECT 34.020 58.105 39.425 58.120 ;
        RECT 33.590 57.210 33.850 58.005 ;
        RECT 34.020 57.380 34.280 58.105 ;
        RECT 34.450 57.210 34.710 57.935 ;
        RECT 34.880 57.380 35.140 58.105 ;
        RECT 35.310 57.210 35.570 57.935 ;
        RECT 35.740 57.380 36.000 58.105 ;
        RECT 36.170 57.210 36.430 57.935 ;
        RECT 36.600 57.380 36.860 58.105 ;
        RECT 37.030 57.210 37.275 57.935 ;
        RECT 37.445 57.380 37.705 58.105 ;
        RECT 37.890 57.210 38.135 57.935 ;
        RECT 38.305 57.380 38.565 58.105 ;
        RECT 38.750 57.210 38.995 57.935 ;
        RECT 39.165 57.380 39.425 58.105 ;
        RECT 39.610 57.210 39.865 57.935 ;
        RECT 40.035 57.380 40.325 58.120 ;
        RECT 33.590 57.205 39.865 57.210 ;
        RECT 40.495 57.205 40.765 57.950 ;
        RECT 44.430 57.640 44.780 58.890 ;
        RECT 46.545 58.280 46.715 59.080 ;
        RECT 47.000 59.035 47.665 59.205 ;
        RECT 47.000 58.780 47.170 59.035 ;
        RECT 47.925 58.985 49.595 59.755 ;
        RECT 49.765 59.080 50.025 59.585 ;
        RECT 50.205 59.375 50.535 59.755 ;
        RECT 50.715 59.205 50.885 59.585 ;
        RECT 46.885 58.450 47.170 58.780 ;
        RECT 47.405 58.485 47.735 58.855 ;
        RECT 47.925 58.465 48.675 58.985 ;
        RECT 47.000 58.305 47.170 58.450 ;
        RECT 41.025 57.205 46.370 57.640 ;
        RECT 46.545 57.375 46.815 58.280 ;
        RECT 47.000 58.135 47.665 58.305 ;
        RECT 48.845 58.295 49.595 58.815 ;
        RECT 46.985 57.205 47.315 57.965 ;
        RECT 47.495 57.375 47.665 58.135 ;
        RECT 47.925 57.205 49.595 58.295 ;
        RECT 49.765 58.280 49.935 59.080 ;
        RECT 50.220 59.035 50.885 59.205 ;
        RECT 50.220 58.780 50.390 59.035 ;
        RECT 51.150 59.015 51.405 59.585 ;
        RECT 51.575 59.355 51.905 59.755 ;
        RECT 52.330 59.220 52.860 59.585 ;
        RECT 53.050 59.415 53.325 59.585 ;
        RECT 53.045 59.245 53.325 59.415 ;
        RECT 52.330 59.185 52.505 59.220 ;
        RECT 51.575 59.015 52.505 59.185 ;
        RECT 50.105 58.450 50.390 58.780 ;
        RECT 50.625 58.485 50.955 58.855 ;
        RECT 50.220 58.305 50.390 58.450 ;
        RECT 51.150 58.345 51.320 59.015 ;
        RECT 51.575 58.845 51.745 59.015 ;
        RECT 51.490 58.515 51.745 58.845 ;
        RECT 51.970 58.515 52.165 58.845 ;
        RECT 49.765 57.375 50.035 58.280 ;
        RECT 50.220 58.135 50.885 58.305 ;
        RECT 50.205 57.205 50.535 57.965 ;
        RECT 50.715 57.375 50.885 58.135 ;
        RECT 51.150 57.375 51.485 58.345 ;
        RECT 51.655 57.205 51.825 58.345 ;
        RECT 51.995 57.545 52.165 58.515 ;
        RECT 52.335 57.885 52.505 59.015 ;
        RECT 52.675 58.225 52.845 59.025 ;
        RECT 53.050 58.425 53.325 59.245 ;
        RECT 53.495 58.225 53.685 59.585 ;
        RECT 53.865 59.220 54.375 59.755 ;
        RECT 54.595 58.945 54.840 59.550 ;
        RECT 55.285 58.985 56.955 59.755 ;
        RECT 57.125 59.030 57.415 59.755 ;
        RECT 57.585 59.210 62.930 59.755 ;
        RECT 63.565 59.255 63.865 59.585 ;
        RECT 64.035 59.275 64.310 59.755 ;
        RECT 53.885 58.775 55.115 58.945 ;
        RECT 52.675 58.055 53.685 58.225 ;
        RECT 53.855 58.210 54.605 58.400 ;
        RECT 52.335 57.715 53.460 57.885 ;
        RECT 53.855 57.545 54.025 58.210 ;
        RECT 54.775 57.965 55.115 58.775 ;
        RECT 55.285 58.465 56.035 58.985 ;
        RECT 56.205 58.295 56.955 58.815 ;
        RECT 59.170 58.380 59.510 59.210 ;
        RECT 51.995 57.375 54.025 57.545 ;
        RECT 54.195 57.205 54.365 57.965 ;
        RECT 54.600 57.555 55.115 57.965 ;
        RECT 55.285 57.205 56.955 58.295 ;
        RECT 57.125 57.205 57.415 58.370 ;
        RECT 60.990 57.640 61.340 58.890 ;
        RECT 63.565 58.345 63.735 59.255 ;
        RECT 64.490 59.105 64.785 59.495 ;
        RECT 64.955 59.275 65.210 59.755 ;
        RECT 65.385 59.105 65.645 59.495 ;
        RECT 65.815 59.275 66.095 59.755 ;
        RECT 66.415 59.105 66.585 59.585 ;
        RECT 66.765 59.275 67.005 59.755 ;
        RECT 67.255 59.105 67.425 59.585 ;
        RECT 67.595 59.275 67.925 59.755 ;
        RECT 68.095 59.105 68.265 59.585 ;
        RECT 63.905 58.515 64.255 59.085 ;
        RECT 64.490 58.935 66.140 59.105 ;
        RECT 66.415 58.935 67.050 59.105 ;
        RECT 67.255 58.935 68.265 59.105 ;
        RECT 68.435 58.955 68.765 59.755 ;
        RECT 69.090 59.205 69.345 59.495 ;
        RECT 69.515 59.375 69.845 59.755 ;
        RECT 69.090 59.035 69.840 59.205 ;
        RECT 64.425 58.595 65.565 58.765 ;
        RECT 64.425 58.345 64.595 58.595 ;
        RECT 65.735 58.425 66.140 58.935 ;
        RECT 66.880 58.765 67.050 58.935 ;
        RECT 67.765 58.905 68.265 58.935 ;
        RECT 66.330 58.525 66.710 58.765 ;
        RECT 66.880 58.595 67.380 58.765 ;
        RECT 63.565 58.175 64.595 58.345 ;
        RECT 65.385 58.255 66.140 58.425 ;
        RECT 66.880 58.355 67.050 58.595 ;
        RECT 67.770 58.395 68.265 58.905 ;
        RECT 57.585 57.205 62.930 57.640 ;
        RECT 63.565 57.375 63.875 58.175 ;
        RECT 65.385 58.005 65.645 58.255 ;
        RECT 66.335 58.185 67.050 58.355 ;
        RECT 67.255 58.225 68.265 58.395 ;
        RECT 64.045 57.205 64.355 58.005 ;
        RECT 64.525 57.835 65.645 58.005 ;
        RECT 64.525 57.375 64.785 57.835 ;
        RECT 64.955 57.205 65.210 57.665 ;
        RECT 65.385 57.375 65.645 57.835 ;
        RECT 65.815 57.205 66.100 58.075 ;
        RECT 66.335 57.375 66.665 58.185 ;
        RECT 66.835 57.205 67.075 58.005 ;
        RECT 67.255 57.375 67.425 58.225 ;
        RECT 67.595 57.205 67.925 58.005 ;
        RECT 68.095 57.375 68.265 58.225 ;
        RECT 68.435 57.205 68.765 58.355 ;
        RECT 69.090 58.215 69.440 58.865 ;
        RECT 69.610 58.045 69.840 59.035 ;
        RECT 69.090 57.875 69.840 58.045 ;
        RECT 69.090 57.375 69.345 57.875 ;
        RECT 69.515 57.205 69.845 57.705 ;
        RECT 70.015 57.375 70.185 59.495 ;
        RECT 70.545 59.395 70.875 59.755 ;
        RECT 71.045 59.365 71.540 59.535 ;
        RECT 71.745 59.365 72.600 59.535 ;
        RECT 70.415 58.175 70.875 59.225 ;
        RECT 70.355 57.390 70.680 58.175 ;
        RECT 71.045 58.005 71.215 59.365 ;
        RECT 71.385 58.455 71.735 59.075 ;
        RECT 71.905 58.855 72.260 59.075 ;
        RECT 71.905 58.265 72.075 58.855 ;
        RECT 72.430 58.655 72.600 59.365 ;
        RECT 73.475 59.295 73.805 59.755 ;
        RECT 74.015 59.395 74.365 59.565 ;
        RECT 72.805 58.825 73.595 59.075 ;
        RECT 74.015 59.005 74.275 59.395 ;
        RECT 74.585 59.305 75.535 59.585 ;
        RECT 75.705 59.315 75.895 59.755 ;
        RECT 76.065 59.375 77.135 59.545 ;
        RECT 73.765 58.655 73.935 58.835 ;
        RECT 71.045 57.835 71.440 58.005 ;
        RECT 71.610 57.875 72.075 58.265 ;
        RECT 72.245 58.485 73.935 58.655 ;
        RECT 71.270 57.705 71.440 57.835 ;
        RECT 72.245 57.705 72.415 58.485 ;
        RECT 74.105 58.315 74.275 59.005 ;
        RECT 72.775 58.145 74.275 58.315 ;
        RECT 74.465 58.345 74.675 59.135 ;
        RECT 74.845 58.515 75.195 59.135 ;
        RECT 75.365 58.525 75.535 59.305 ;
        RECT 76.065 59.145 76.235 59.375 ;
        RECT 75.705 58.975 76.235 59.145 ;
        RECT 75.705 58.695 75.925 58.975 ;
        RECT 76.405 58.805 76.645 59.205 ;
        RECT 75.365 58.355 75.770 58.525 ;
        RECT 76.105 58.435 76.645 58.805 ;
        RECT 76.815 59.020 77.135 59.375 ;
        RECT 77.380 59.295 77.685 59.755 ;
        RECT 77.855 59.045 78.110 59.575 ;
        RECT 76.815 58.845 77.140 59.020 ;
        RECT 76.815 58.545 77.730 58.845 ;
        RECT 76.990 58.515 77.730 58.545 ;
        RECT 74.465 58.185 75.140 58.345 ;
        RECT 75.600 58.265 75.770 58.355 ;
        RECT 74.465 58.175 75.430 58.185 ;
        RECT 74.105 58.005 74.275 58.145 ;
        RECT 70.850 57.205 71.100 57.665 ;
        RECT 71.270 57.375 71.520 57.705 ;
        RECT 71.735 57.375 72.415 57.705 ;
        RECT 72.585 57.805 73.660 57.975 ;
        RECT 74.105 57.835 74.665 58.005 ;
        RECT 74.970 57.885 75.430 58.175 ;
        RECT 75.600 58.095 76.820 58.265 ;
        RECT 72.585 57.465 72.755 57.805 ;
        RECT 72.990 57.205 73.320 57.635 ;
        RECT 73.490 57.465 73.660 57.805 ;
        RECT 73.955 57.205 74.325 57.665 ;
        RECT 74.495 57.375 74.665 57.835 ;
        RECT 75.600 57.715 75.770 58.095 ;
        RECT 76.990 57.925 77.160 58.515 ;
        RECT 77.900 58.395 78.110 59.045 ;
        RECT 74.900 57.375 75.770 57.715 ;
        RECT 76.360 57.755 77.160 57.925 ;
        RECT 75.940 57.205 76.190 57.665 ;
        RECT 76.360 57.465 76.530 57.755 ;
        RECT 76.710 57.205 77.040 57.585 ;
        RECT 77.380 57.205 77.685 58.345 ;
        RECT 77.855 57.515 78.110 58.395 ;
        RECT 78.285 59.080 78.545 59.585 ;
        RECT 78.725 59.375 79.055 59.755 ;
        RECT 79.235 59.205 79.405 59.585 ;
        RECT 78.285 58.280 78.455 59.080 ;
        RECT 78.740 59.035 79.405 59.205 ;
        RECT 78.740 58.780 78.910 59.035 ;
        RECT 79.665 58.985 81.335 59.755 ;
        RECT 78.625 58.450 78.910 58.780 ;
        RECT 79.145 58.485 79.475 58.855 ;
        RECT 79.665 58.465 80.415 58.985 ;
        RECT 81.545 58.935 81.775 59.755 ;
        RECT 81.945 58.955 82.275 59.585 ;
        RECT 78.740 58.305 78.910 58.450 ;
        RECT 78.285 57.375 78.555 58.280 ;
        RECT 78.740 58.135 79.405 58.305 ;
        RECT 80.585 58.295 81.335 58.815 ;
        RECT 81.525 58.515 81.855 58.765 ;
        RECT 82.025 58.355 82.275 58.955 ;
        RECT 82.445 58.935 82.655 59.755 ;
        RECT 82.885 59.030 83.175 59.755 ;
        RECT 83.345 59.015 83.730 59.585 ;
        RECT 83.900 59.295 84.225 59.755 ;
        RECT 84.745 59.125 85.025 59.585 ;
        RECT 78.725 57.205 79.055 57.965 ;
        RECT 79.235 57.375 79.405 58.135 ;
        RECT 79.665 57.205 81.335 58.295 ;
        RECT 81.545 57.205 81.775 58.345 ;
        RECT 81.945 57.375 82.275 58.355 ;
        RECT 82.445 57.205 82.655 58.345 ;
        RECT 82.885 57.205 83.175 58.370 ;
        RECT 83.345 58.345 83.625 59.015 ;
        RECT 83.900 58.955 85.025 59.125 ;
        RECT 83.900 58.845 84.350 58.955 ;
        RECT 83.795 58.515 84.350 58.845 ;
        RECT 85.215 58.785 85.615 59.585 ;
        RECT 86.015 59.295 86.285 59.755 ;
        RECT 86.455 59.125 86.740 59.585 ;
        RECT 83.345 57.375 83.730 58.345 ;
        RECT 83.900 58.055 84.350 58.515 ;
        RECT 84.520 58.225 85.615 58.785 ;
        RECT 83.900 57.835 85.025 58.055 ;
        RECT 83.900 57.205 84.225 57.665 ;
        RECT 84.745 57.375 85.025 57.835 ;
        RECT 85.215 57.375 85.615 58.225 ;
        RECT 85.785 58.955 86.740 59.125 ;
        RECT 87.950 59.205 88.205 59.495 ;
        RECT 88.375 59.375 88.705 59.755 ;
        RECT 87.950 59.035 88.700 59.205 ;
        RECT 85.785 58.055 85.995 58.955 ;
        RECT 86.165 58.225 86.855 58.785 ;
        RECT 87.950 58.215 88.300 58.865 ;
        RECT 85.785 57.835 86.740 58.055 ;
        RECT 88.470 58.045 88.700 59.035 ;
        RECT 86.015 57.205 86.285 57.665 ;
        RECT 86.455 57.375 86.740 57.835 ;
        RECT 87.950 57.875 88.700 58.045 ;
        RECT 87.950 57.375 88.205 57.875 ;
        RECT 88.375 57.205 88.705 57.705 ;
        RECT 88.875 57.375 89.045 59.495 ;
        RECT 89.405 59.395 89.735 59.755 ;
        RECT 89.905 59.365 90.400 59.535 ;
        RECT 90.605 59.365 91.460 59.535 ;
        RECT 89.275 58.175 89.735 59.225 ;
        RECT 89.215 57.390 89.540 58.175 ;
        RECT 89.905 58.005 90.075 59.365 ;
        RECT 90.245 58.455 90.595 59.075 ;
        RECT 90.765 58.855 91.120 59.075 ;
        RECT 90.765 58.265 90.935 58.855 ;
        RECT 91.290 58.655 91.460 59.365 ;
        RECT 92.335 59.295 92.665 59.755 ;
        RECT 92.875 59.395 93.225 59.565 ;
        RECT 91.665 58.825 92.455 59.075 ;
        RECT 92.875 59.005 93.135 59.395 ;
        RECT 93.445 59.305 94.395 59.585 ;
        RECT 94.565 59.315 94.755 59.755 ;
        RECT 94.925 59.375 95.995 59.545 ;
        RECT 92.625 58.655 92.795 58.835 ;
        RECT 89.905 57.835 90.300 58.005 ;
        RECT 90.470 57.875 90.935 58.265 ;
        RECT 91.105 58.485 92.795 58.655 ;
        RECT 90.130 57.705 90.300 57.835 ;
        RECT 91.105 57.705 91.275 58.485 ;
        RECT 92.965 58.315 93.135 59.005 ;
        RECT 91.635 58.145 93.135 58.315 ;
        RECT 93.325 58.345 93.535 59.135 ;
        RECT 93.705 58.515 94.055 59.135 ;
        RECT 94.225 58.525 94.395 59.305 ;
        RECT 94.925 59.145 95.095 59.375 ;
        RECT 94.565 58.975 95.095 59.145 ;
        RECT 94.565 58.695 94.785 58.975 ;
        RECT 95.265 58.805 95.505 59.205 ;
        RECT 94.225 58.355 94.630 58.525 ;
        RECT 94.965 58.435 95.505 58.805 ;
        RECT 95.675 59.020 95.995 59.375 ;
        RECT 96.240 59.295 96.545 59.755 ;
        RECT 96.715 59.045 96.970 59.575 ;
        RECT 95.675 58.845 96.000 59.020 ;
        RECT 95.675 58.545 96.590 58.845 ;
        RECT 95.850 58.515 96.590 58.545 ;
        RECT 93.325 58.185 94.000 58.345 ;
        RECT 94.460 58.265 94.630 58.355 ;
        RECT 93.325 58.175 94.290 58.185 ;
        RECT 92.965 58.005 93.135 58.145 ;
        RECT 89.710 57.205 89.960 57.665 ;
        RECT 90.130 57.375 90.380 57.705 ;
        RECT 90.595 57.375 91.275 57.705 ;
        RECT 91.445 57.805 92.520 57.975 ;
        RECT 92.965 57.835 93.525 58.005 ;
        RECT 93.830 57.885 94.290 58.175 ;
        RECT 94.460 58.095 95.680 58.265 ;
        RECT 91.445 57.465 91.615 57.805 ;
        RECT 91.850 57.205 92.180 57.635 ;
        RECT 92.350 57.465 92.520 57.805 ;
        RECT 92.815 57.205 93.185 57.665 ;
        RECT 93.355 57.375 93.525 57.835 ;
        RECT 94.460 57.715 94.630 58.095 ;
        RECT 95.850 57.925 96.020 58.515 ;
        RECT 96.760 58.395 96.970 59.045 ;
        RECT 93.760 57.375 94.630 57.715 ;
        RECT 95.220 57.755 96.020 57.925 ;
        RECT 94.800 57.205 95.050 57.665 ;
        RECT 95.220 57.465 95.390 57.755 ;
        RECT 95.570 57.205 95.900 57.585 ;
        RECT 96.240 57.205 96.545 58.345 ;
        RECT 96.715 57.515 96.970 58.395 ;
        RECT 97.150 59.045 97.405 59.575 ;
        RECT 97.575 59.295 97.880 59.755 ;
        RECT 98.125 59.375 99.195 59.545 ;
        RECT 97.150 58.395 97.360 59.045 ;
        RECT 98.125 59.020 98.445 59.375 ;
        RECT 98.120 58.845 98.445 59.020 ;
        RECT 97.530 58.545 98.445 58.845 ;
        RECT 98.615 58.805 98.855 59.205 ;
        RECT 99.025 59.145 99.195 59.375 ;
        RECT 99.365 59.315 99.555 59.755 ;
        RECT 99.725 59.305 100.675 59.585 ;
        RECT 100.895 59.395 101.245 59.565 ;
        RECT 99.025 58.975 99.555 59.145 ;
        RECT 97.530 58.515 98.270 58.545 ;
        RECT 97.150 57.515 97.405 58.395 ;
        RECT 97.575 57.205 97.880 58.345 ;
        RECT 98.100 57.925 98.270 58.515 ;
        RECT 98.615 58.435 99.155 58.805 ;
        RECT 99.335 58.695 99.555 58.975 ;
        RECT 99.725 58.525 99.895 59.305 ;
        RECT 99.490 58.355 99.895 58.525 ;
        RECT 100.065 58.515 100.415 59.135 ;
        RECT 99.490 58.265 99.660 58.355 ;
        RECT 100.585 58.345 100.795 59.135 ;
        RECT 98.440 58.095 99.660 58.265 ;
        RECT 100.120 58.185 100.795 58.345 ;
        RECT 98.100 57.755 98.900 57.925 ;
        RECT 98.220 57.205 98.550 57.585 ;
        RECT 98.730 57.465 98.900 57.755 ;
        RECT 99.490 57.715 99.660 58.095 ;
        RECT 99.830 58.175 100.795 58.185 ;
        RECT 100.985 59.005 101.245 59.395 ;
        RECT 101.455 59.295 101.785 59.755 ;
        RECT 102.660 59.365 103.515 59.535 ;
        RECT 103.720 59.365 104.215 59.535 ;
        RECT 104.385 59.395 104.715 59.755 ;
        RECT 100.985 58.315 101.155 59.005 ;
        RECT 101.325 58.655 101.495 58.835 ;
        RECT 101.665 58.825 102.455 59.075 ;
        RECT 102.660 58.655 102.830 59.365 ;
        RECT 103.000 58.855 103.355 59.075 ;
        RECT 101.325 58.485 103.015 58.655 ;
        RECT 99.830 57.885 100.290 58.175 ;
        RECT 100.985 58.145 102.485 58.315 ;
        RECT 100.985 58.005 101.155 58.145 ;
        RECT 100.595 57.835 101.155 58.005 ;
        RECT 99.070 57.205 99.320 57.665 ;
        RECT 99.490 57.375 100.360 57.715 ;
        RECT 100.595 57.375 100.765 57.835 ;
        RECT 101.600 57.805 102.675 57.975 ;
        RECT 100.935 57.205 101.305 57.665 ;
        RECT 101.600 57.465 101.770 57.805 ;
        RECT 101.940 57.205 102.270 57.635 ;
        RECT 102.505 57.465 102.675 57.805 ;
        RECT 102.845 57.705 103.015 58.485 ;
        RECT 103.185 58.265 103.355 58.855 ;
        RECT 103.525 58.455 103.875 59.075 ;
        RECT 103.185 57.875 103.650 58.265 ;
        RECT 104.045 58.005 104.215 59.365 ;
        RECT 104.385 58.175 104.845 59.225 ;
        RECT 103.820 57.835 104.215 58.005 ;
        RECT 103.820 57.705 103.990 57.835 ;
        RECT 102.845 57.375 103.525 57.705 ;
        RECT 103.740 57.375 103.990 57.705 ;
        RECT 104.160 57.205 104.410 57.665 ;
        RECT 104.580 57.390 104.905 58.175 ;
        RECT 105.075 57.375 105.245 59.495 ;
        RECT 105.415 59.375 105.745 59.755 ;
        RECT 105.915 59.205 106.170 59.495 ;
        RECT 105.420 59.035 106.170 59.205 ;
        RECT 106.435 59.205 106.605 59.585 ;
        RECT 106.785 59.375 107.115 59.755 ;
        RECT 106.435 59.035 107.100 59.205 ;
        RECT 107.295 59.080 107.555 59.585 ;
        RECT 105.420 58.045 105.650 59.035 ;
        RECT 105.820 58.215 106.170 58.865 ;
        RECT 106.365 58.485 106.695 58.855 ;
        RECT 106.930 58.780 107.100 59.035 ;
        RECT 106.930 58.450 107.215 58.780 ;
        RECT 106.930 58.305 107.100 58.450 ;
        RECT 106.435 58.135 107.100 58.305 ;
        RECT 107.385 58.280 107.555 59.080 ;
        RECT 108.645 59.030 108.935 59.755 ;
        RECT 109.105 59.210 114.450 59.755 ;
        RECT 110.690 58.380 111.030 59.210 ;
        RECT 114.625 58.985 117.215 59.755 ;
        RECT 117.385 59.005 118.595 59.755 ;
        RECT 105.420 57.875 106.170 58.045 ;
        RECT 105.415 57.205 105.745 57.705 ;
        RECT 105.915 57.375 106.170 57.875 ;
        RECT 106.435 57.375 106.605 58.135 ;
        RECT 106.785 57.205 107.115 57.965 ;
        RECT 107.285 57.375 107.555 58.280 ;
        RECT 108.645 57.205 108.935 58.370 ;
        RECT 112.510 57.640 112.860 58.890 ;
        RECT 114.625 58.465 115.835 58.985 ;
        RECT 116.005 58.295 117.215 58.815 ;
        RECT 109.105 57.205 114.450 57.640 ;
        RECT 114.625 57.205 117.215 58.295 ;
        RECT 117.385 58.295 117.905 58.835 ;
        RECT 118.075 58.465 118.595 59.005 ;
        RECT 117.385 57.205 118.595 58.295 ;
        RECT 5.520 57.035 118.680 57.205 ;
        RECT 5.605 55.945 6.815 57.035 ;
        RECT 6.985 55.945 8.195 57.035 ;
        RECT 8.370 56.365 8.625 56.865 ;
        RECT 8.795 56.535 9.125 57.035 ;
        RECT 8.370 56.195 9.120 56.365 ;
        RECT 5.605 55.235 6.125 55.775 ;
        RECT 6.295 55.405 6.815 55.945 ;
        RECT 6.985 55.235 7.505 55.775 ;
        RECT 7.675 55.405 8.195 55.945 ;
        RECT 8.370 55.375 8.720 56.025 ;
        RECT 5.605 54.485 6.815 55.235 ;
        RECT 6.985 54.485 8.195 55.235 ;
        RECT 8.890 55.205 9.120 56.195 ;
        RECT 8.370 55.035 9.120 55.205 ;
        RECT 8.370 54.745 8.625 55.035 ;
        RECT 8.795 54.485 9.125 54.865 ;
        RECT 9.295 54.745 9.465 56.865 ;
        RECT 9.635 56.065 9.960 56.850 ;
        RECT 10.130 56.575 10.380 57.035 ;
        RECT 10.550 56.535 10.800 56.865 ;
        RECT 11.015 56.535 11.695 56.865 ;
        RECT 10.550 56.405 10.720 56.535 ;
        RECT 10.325 56.235 10.720 56.405 ;
        RECT 9.695 55.015 10.155 56.065 ;
        RECT 10.325 54.875 10.495 56.235 ;
        RECT 10.890 55.975 11.355 56.365 ;
        RECT 10.665 55.165 11.015 55.785 ;
        RECT 11.185 55.385 11.355 55.975 ;
        RECT 11.525 55.755 11.695 56.535 ;
        RECT 11.865 56.435 12.035 56.775 ;
        RECT 12.270 56.605 12.600 57.035 ;
        RECT 12.770 56.435 12.940 56.775 ;
        RECT 13.235 56.575 13.605 57.035 ;
        RECT 11.865 56.265 12.940 56.435 ;
        RECT 13.775 56.405 13.945 56.865 ;
        RECT 14.180 56.525 15.050 56.865 ;
        RECT 15.220 56.575 15.470 57.035 ;
        RECT 13.385 56.235 13.945 56.405 ;
        RECT 13.385 56.095 13.555 56.235 ;
        RECT 12.055 55.925 13.555 56.095 ;
        RECT 14.250 56.065 14.710 56.355 ;
        RECT 11.525 55.585 13.215 55.755 ;
        RECT 11.185 55.165 11.540 55.385 ;
        RECT 11.710 54.875 11.880 55.585 ;
        RECT 12.085 55.165 12.875 55.415 ;
        RECT 13.045 55.405 13.215 55.585 ;
        RECT 13.385 55.235 13.555 55.925 ;
        RECT 9.825 54.485 10.155 54.845 ;
        RECT 10.325 54.705 10.820 54.875 ;
        RECT 11.025 54.705 11.880 54.875 ;
        RECT 12.755 54.485 13.085 54.945 ;
        RECT 13.295 54.845 13.555 55.235 ;
        RECT 13.745 56.055 14.710 56.065 ;
        RECT 14.880 56.145 15.050 56.525 ;
        RECT 15.640 56.485 15.810 56.775 ;
        RECT 15.990 56.655 16.320 57.035 ;
        RECT 15.640 56.315 16.440 56.485 ;
        RECT 13.745 55.895 14.420 56.055 ;
        RECT 14.880 55.975 16.100 56.145 ;
        RECT 13.745 55.105 13.955 55.895 ;
        RECT 14.880 55.885 15.050 55.975 ;
        RECT 14.125 55.105 14.475 55.725 ;
        RECT 14.645 55.715 15.050 55.885 ;
        RECT 14.645 54.935 14.815 55.715 ;
        RECT 14.985 55.265 15.205 55.545 ;
        RECT 15.385 55.435 15.925 55.805 ;
        RECT 16.270 55.725 16.440 56.315 ;
        RECT 16.660 55.895 16.965 57.035 ;
        RECT 17.135 55.845 17.390 56.725 ;
        RECT 18.485 55.870 18.775 57.035 ;
        RECT 18.945 55.895 19.330 56.865 ;
        RECT 19.500 56.575 19.825 57.035 ;
        RECT 20.345 56.405 20.625 56.865 ;
        RECT 19.500 56.185 20.625 56.405 ;
        RECT 16.270 55.695 17.010 55.725 ;
        RECT 14.985 55.095 15.515 55.265 ;
        RECT 13.295 54.675 13.645 54.845 ;
        RECT 13.865 54.655 14.815 54.935 ;
        RECT 14.985 54.485 15.175 54.925 ;
        RECT 15.345 54.865 15.515 55.095 ;
        RECT 15.685 55.035 15.925 55.435 ;
        RECT 16.095 55.395 17.010 55.695 ;
        RECT 16.095 55.220 16.420 55.395 ;
        RECT 16.095 54.865 16.415 55.220 ;
        RECT 17.180 55.195 17.390 55.845 ;
        RECT 18.945 55.225 19.225 55.895 ;
        RECT 19.500 55.725 19.950 56.185 ;
        RECT 20.815 56.015 21.215 56.865 ;
        RECT 21.615 56.575 21.885 57.035 ;
        RECT 22.055 56.405 22.340 56.865 ;
        RECT 19.395 55.395 19.950 55.725 ;
        RECT 20.120 55.455 21.215 56.015 ;
        RECT 19.500 55.285 19.950 55.395 ;
        RECT 15.345 54.695 16.415 54.865 ;
        RECT 16.660 54.485 16.965 54.945 ;
        RECT 17.135 54.665 17.390 55.195 ;
        RECT 18.485 54.485 18.775 55.210 ;
        RECT 18.945 54.655 19.330 55.225 ;
        RECT 19.500 55.115 20.625 55.285 ;
        RECT 19.500 54.485 19.825 54.945 ;
        RECT 20.345 54.655 20.625 55.115 ;
        RECT 20.815 54.655 21.215 55.455 ;
        RECT 21.385 56.185 22.340 56.405 ;
        RECT 21.385 55.285 21.595 56.185 ;
        RECT 21.765 55.455 22.455 56.015 ;
        RECT 22.625 55.895 23.010 56.865 ;
        RECT 23.180 56.575 23.505 57.035 ;
        RECT 24.025 56.405 24.305 56.865 ;
        RECT 23.180 56.185 24.305 56.405 ;
        RECT 21.385 55.115 22.340 55.285 ;
        RECT 21.615 54.485 21.885 54.945 ;
        RECT 22.055 54.655 22.340 55.115 ;
        RECT 22.625 55.225 22.905 55.895 ;
        RECT 23.180 55.725 23.630 56.185 ;
        RECT 24.495 56.015 24.895 56.865 ;
        RECT 25.295 56.575 25.565 57.035 ;
        RECT 25.735 56.405 26.020 56.865 ;
        RECT 23.075 55.395 23.630 55.725 ;
        RECT 23.800 55.455 24.895 56.015 ;
        RECT 23.180 55.285 23.630 55.395 ;
        RECT 22.625 54.655 23.010 55.225 ;
        RECT 23.180 55.115 24.305 55.285 ;
        RECT 23.180 54.485 23.505 54.945 ;
        RECT 24.025 54.655 24.305 55.115 ;
        RECT 24.495 54.655 24.895 55.455 ;
        RECT 25.065 56.185 26.020 56.405 ;
        RECT 26.395 56.365 26.565 56.865 ;
        RECT 26.735 56.535 27.065 57.035 ;
        RECT 26.395 56.195 27.060 56.365 ;
        RECT 25.065 55.285 25.275 56.185 ;
        RECT 25.445 55.455 26.135 56.015 ;
        RECT 26.310 55.375 26.660 56.025 ;
        RECT 25.065 55.115 26.020 55.285 ;
        RECT 26.830 55.205 27.060 56.195 ;
        RECT 25.295 54.485 25.565 54.945 ;
        RECT 25.735 54.655 26.020 55.115 ;
        RECT 26.395 55.035 27.060 55.205 ;
        RECT 26.395 54.745 26.565 55.035 ;
        RECT 26.735 54.485 27.065 54.865 ;
        RECT 27.235 54.745 27.460 56.865 ;
        RECT 27.675 56.535 28.005 57.035 ;
        RECT 28.175 56.365 28.345 56.865 ;
        RECT 28.580 56.650 29.410 56.820 ;
        RECT 29.650 56.655 30.030 57.035 ;
        RECT 27.650 56.195 28.345 56.365 ;
        RECT 27.650 55.225 27.820 56.195 ;
        RECT 27.990 55.405 28.400 56.025 ;
        RECT 28.570 55.975 29.070 56.355 ;
        RECT 27.650 55.035 28.345 55.225 ;
        RECT 28.570 55.105 28.790 55.975 ;
        RECT 29.240 55.805 29.410 56.650 ;
        RECT 30.210 56.485 30.380 56.775 ;
        RECT 30.550 56.655 30.880 57.035 ;
        RECT 31.350 56.565 31.980 56.815 ;
        RECT 32.160 56.655 32.580 57.035 ;
        RECT 31.810 56.485 31.980 56.565 ;
        RECT 32.780 56.485 33.020 56.775 ;
        RECT 29.580 56.235 30.950 56.485 ;
        RECT 29.580 55.975 29.830 56.235 ;
        RECT 30.340 55.805 30.590 55.965 ;
        RECT 29.240 55.635 30.590 55.805 ;
        RECT 29.240 55.595 29.660 55.635 ;
        RECT 28.970 55.045 29.320 55.415 ;
        RECT 27.675 54.485 28.005 54.865 ;
        RECT 28.175 54.705 28.345 55.035 ;
        RECT 29.490 54.865 29.660 55.595 ;
        RECT 30.760 55.465 30.950 56.235 ;
        RECT 29.830 55.135 30.240 55.465 ;
        RECT 30.530 55.125 30.950 55.465 ;
        RECT 31.120 56.055 31.640 56.365 ;
        RECT 31.810 56.315 33.020 56.485 ;
        RECT 33.250 56.345 33.580 57.035 ;
        RECT 31.120 55.295 31.290 56.055 ;
        RECT 31.460 55.465 31.640 55.875 ;
        RECT 31.810 55.805 31.980 56.315 ;
        RECT 33.750 56.165 33.920 56.775 ;
        RECT 34.190 56.315 34.520 56.825 ;
        RECT 33.750 56.145 34.070 56.165 ;
        RECT 32.150 55.975 34.070 56.145 ;
        RECT 31.810 55.635 33.710 55.805 ;
        RECT 32.040 55.295 32.370 55.415 ;
        RECT 31.120 55.125 32.370 55.295 ;
        RECT 28.645 54.665 29.660 54.865 ;
        RECT 29.830 54.485 30.240 54.925 ;
        RECT 30.530 54.695 30.780 55.125 ;
        RECT 30.980 54.485 31.300 54.945 ;
        RECT 32.540 54.875 32.710 55.635 ;
        RECT 33.380 55.575 33.710 55.635 ;
        RECT 32.900 55.405 33.230 55.465 ;
        RECT 32.900 55.135 33.560 55.405 ;
        RECT 33.880 55.080 34.070 55.975 ;
        RECT 31.860 54.705 32.710 54.875 ;
        RECT 32.910 54.485 33.570 54.965 ;
        RECT 33.750 54.750 34.070 55.080 ;
        RECT 34.270 55.725 34.520 56.315 ;
        RECT 34.700 56.235 34.985 57.035 ;
        RECT 35.165 56.055 35.420 56.725 ;
        RECT 35.240 56.015 35.420 56.055 ;
        RECT 35.240 55.845 35.505 56.015 ;
        RECT 35.970 55.895 36.305 56.865 ;
        RECT 36.475 55.895 36.645 57.035 ;
        RECT 36.815 56.695 38.845 56.865 ;
        RECT 34.270 55.395 35.070 55.725 ;
        RECT 34.270 54.745 34.520 55.395 ;
        RECT 35.240 55.195 35.420 55.845 ;
        RECT 34.700 54.485 34.985 54.945 ;
        RECT 35.165 54.665 35.420 55.195 ;
        RECT 35.970 55.225 36.140 55.895 ;
        RECT 36.815 55.725 36.985 56.695 ;
        RECT 36.310 55.395 36.565 55.725 ;
        RECT 36.790 55.395 36.985 55.725 ;
        RECT 37.155 56.355 38.280 56.525 ;
        RECT 36.395 55.225 36.565 55.395 ;
        RECT 37.155 55.225 37.325 56.355 ;
        RECT 35.970 54.655 36.225 55.225 ;
        RECT 36.395 55.055 37.325 55.225 ;
        RECT 37.495 56.015 38.505 56.185 ;
        RECT 37.495 55.215 37.665 56.015 ;
        RECT 37.870 55.675 38.145 55.815 ;
        RECT 37.865 55.505 38.145 55.675 ;
        RECT 37.150 55.020 37.325 55.055 ;
        RECT 36.395 54.485 36.725 54.885 ;
        RECT 37.150 54.655 37.680 55.020 ;
        RECT 37.870 54.655 38.145 55.505 ;
        RECT 38.315 54.655 38.505 56.015 ;
        RECT 38.675 56.030 38.845 56.695 ;
        RECT 39.015 56.275 39.185 57.035 ;
        RECT 39.420 56.275 39.935 56.685 ;
        RECT 38.675 55.840 39.425 56.030 ;
        RECT 39.595 55.465 39.935 56.275 ;
        RECT 40.105 55.945 43.615 57.035 ;
        RECT 38.705 55.295 39.935 55.465 ;
        RECT 38.685 54.485 39.195 55.020 ;
        RECT 39.415 54.690 39.660 55.295 ;
        RECT 40.105 55.255 41.755 55.775 ;
        RECT 41.925 55.425 43.615 55.945 ;
        RECT 44.245 55.870 44.535 57.035 ;
        RECT 45.665 55.895 45.895 57.035 ;
        RECT 46.065 55.885 46.395 56.865 ;
        RECT 46.565 55.895 46.775 57.035 ;
        RECT 47.045 55.895 47.275 57.035 ;
        RECT 47.445 55.885 47.775 56.865 ;
        RECT 47.945 55.895 48.155 57.035 ;
        RECT 48.475 56.365 48.645 56.865 ;
        RECT 48.815 56.535 49.145 57.035 ;
        RECT 48.475 56.195 49.140 56.365 ;
        RECT 45.645 55.475 45.975 55.725 ;
        RECT 40.105 54.485 43.615 55.255 ;
        RECT 44.245 54.485 44.535 55.210 ;
        RECT 45.665 54.485 45.895 55.305 ;
        RECT 46.145 55.285 46.395 55.885 ;
        RECT 47.025 55.475 47.355 55.725 ;
        RECT 46.065 54.655 46.395 55.285 ;
        RECT 46.565 54.485 46.775 55.305 ;
        RECT 47.045 54.485 47.275 55.305 ;
        RECT 47.525 55.285 47.775 55.885 ;
        RECT 48.390 55.375 48.740 56.025 ;
        RECT 47.445 54.655 47.775 55.285 ;
        RECT 47.945 54.485 48.155 55.305 ;
        RECT 48.910 55.205 49.140 56.195 ;
        RECT 48.475 55.035 49.140 55.205 ;
        RECT 48.475 54.745 48.645 55.035 ;
        RECT 48.815 54.485 49.145 54.865 ;
        RECT 49.315 54.745 49.540 56.865 ;
        RECT 49.755 56.535 50.085 57.035 ;
        RECT 50.255 56.365 50.425 56.865 ;
        RECT 50.660 56.650 51.490 56.820 ;
        RECT 51.730 56.655 52.110 57.035 ;
        RECT 49.730 56.195 50.425 56.365 ;
        RECT 49.730 55.225 49.900 56.195 ;
        RECT 50.070 55.405 50.480 56.025 ;
        RECT 50.650 55.975 51.150 56.355 ;
        RECT 49.730 55.035 50.425 55.225 ;
        RECT 50.650 55.105 50.870 55.975 ;
        RECT 51.320 55.805 51.490 56.650 ;
        RECT 52.290 56.485 52.460 56.775 ;
        RECT 52.630 56.655 52.960 57.035 ;
        RECT 53.430 56.565 54.060 56.815 ;
        RECT 54.240 56.655 54.660 57.035 ;
        RECT 53.890 56.485 54.060 56.565 ;
        RECT 54.860 56.485 55.100 56.775 ;
        RECT 51.660 56.235 53.030 56.485 ;
        RECT 51.660 55.975 51.910 56.235 ;
        RECT 52.420 55.805 52.670 55.965 ;
        RECT 51.320 55.635 52.670 55.805 ;
        RECT 51.320 55.595 51.740 55.635 ;
        RECT 51.050 55.045 51.400 55.415 ;
        RECT 49.755 54.485 50.085 54.865 ;
        RECT 50.255 54.705 50.425 55.035 ;
        RECT 51.570 54.865 51.740 55.595 ;
        RECT 52.840 55.465 53.030 56.235 ;
        RECT 51.910 55.135 52.320 55.465 ;
        RECT 52.610 55.125 53.030 55.465 ;
        RECT 53.200 56.055 53.720 56.365 ;
        RECT 53.890 56.315 55.100 56.485 ;
        RECT 55.330 56.345 55.660 57.035 ;
        RECT 53.200 55.295 53.370 56.055 ;
        RECT 53.540 55.465 53.720 55.875 ;
        RECT 53.890 55.805 54.060 56.315 ;
        RECT 55.830 56.165 56.000 56.775 ;
        RECT 56.270 56.315 56.600 56.825 ;
        RECT 55.830 56.145 56.150 56.165 ;
        RECT 54.230 55.975 56.150 56.145 ;
        RECT 53.890 55.635 55.790 55.805 ;
        RECT 54.120 55.295 54.450 55.415 ;
        RECT 53.200 55.125 54.450 55.295 ;
        RECT 50.725 54.665 51.740 54.865 ;
        RECT 51.910 54.485 52.320 54.925 ;
        RECT 52.610 54.695 52.860 55.125 ;
        RECT 53.060 54.485 53.380 54.945 ;
        RECT 54.620 54.875 54.790 55.635 ;
        RECT 55.460 55.575 55.790 55.635 ;
        RECT 54.980 55.405 55.310 55.465 ;
        RECT 54.980 55.135 55.640 55.405 ;
        RECT 55.960 55.080 56.150 55.975 ;
        RECT 53.940 54.705 54.790 54.875 ;
        RECT 54.990 54.485 55.650 54.965 ;
        RECT 55.830 54.750 56.150 55.080 ;
        RECT 56.350 55.725 56.600 56.315 ;
        RECT 56.780 56.235 57.065 57.035 ;
        RECT 57.245 56.695 57.500 56.725 ;
        RECT 57.245 56.525 57.585 56.695 ;
        RECT 57.245 56.055 57.500 56.525 ;
        RECT 56.350 55.395 57.150 55.725 ;
        RECT 56.350 54.745 56.600 55.395 ;
        RECT 57.320 55.195 57.500 56.055 ;
        RECT 58.045 55.945 59.715 57.035 ;
        RECT 56.780 54.485 57.065 54.945 ;
        RECT 57.245 54.665 57.500 55.195 ;
        RECT 58.045 55.255 58.795 55.775 ;
        RECT 58.965 55.425 59.715 55.945 ;
        RECT 59.885 56.445 60.585 56.865 ;
        RECT 60.785 56.675 61.115 57.035 ;
        RECT 61.285 56.445 61.615 56.845 ;
        RECT 59.885 56.215 61.615 56.445 ;
        RECT 59.885 55.335 60.090 56.215 ;
        RECT 60.260 55.475 60.590 56.015 ;
        RECT 60.765 55.725 61.090 56.015 ;
        RECT 61.285 55.995 61.615 56.215 ;
        RECT 61.785 55.725 61.955 56.650 ;
        RECT 62.135 55.975 62.465 57.035 ;
        RECT 62.700 56.165 62.985 57.035 ;
        RECT 63.155 56.405 63.415 56.865 ;
        RECT 63.590 56.575 63.845 57.035 ;
        RECT 64.015 56.405 64.275 56.865 ;
        RECT 63.155 56.235 64.275 56.405 ;
        RECT 64.445 56.235 64.755 57.035 ;
        RECT 63.155 55.985 63.415 56.235 ;
        RECT 64.925 56.065 65.235 56.865 ;
        RECT 62.660 55.815 63.415 55.985 ;
        RECT 64.205 55.895 65.235 56.065 ;
        RECT 60.765 55.395 61.260 55.725 ;
        RECT 61.580 55.395 61.955 55.725 ;
        RECT 62.165 55.395 62.475 55.725 ;
        RECT 58.045 54.485 59.715 55.255 ;
        RECT 59.885 55.245 60.115 55.335 ;
        RECT 62.660 55.305 63.065 55.815 ;
        RECT 64.205 55.645 64.375 55.895 ;
        RECT 63.235 55.475 64.375 55.645 ;
        RECT 59.885 54.655 60.595 55.245 ;
        RECT 61.105 55.015 62.465 55.225 ;
        RECT 62.660 55.135 64.310 55.305 ;
        RECT 64.545 55.155 64.895 55.725 ;
        RECT 61.105 54.655 61.435 55.015 ;
        RECT 61.635 54.485 61.965 54.845 ;
        RECT 62.135 54.655 62.465 55.015 ;
        RECT 62.705 54.485 62.985 54.965 ;
        RECT 63.155 54.745 63.415 55.135 ;
        RECT 63.590 54.485 63.845 54.965 ;
        RECT 64.015 54.745 64.310 55.135 ;
        RECT 65.065 54.985 65.235 55.895 ;
        RECT 64.490 54.485 64.765 54.965 ;
        RECT 64.935 54.655 65.235 54.985 ;
        RECT 65.405 56.065 65.715 56.865 ;
        RECT 65.885 56.235 66.195 57.035 ;
        RECT 66.365 56.405 66.625 56.865 ;
        RECT 66.795 56.575 67.050 57.035 ;
        RECT 67.225 56.405 67.485 56.865 ;
        RECT 66.365 56.235 67.485 56.405 ;
        RECT 65.405 55.895 66.435 56.065 ;
        RECT 65.405 54.985 65.575 55.895 ;
        RECT 65.745 55.155 66.095 55.725 ;
        RECT 66.265 55.645 66.435 55.895 ;
        RECT 67.225 55.985 67.485 56.235 ;
        RECT 67.655 56.165 67.940 57.035 ;
        RECT 67.225 55.815 67.980 55.985 ;
        RECT 68.165 55.945 69.835 57.035 ;
        RECT 66.265 55.475 67.405 55.645 ;
        RECT 67.575 55.305 67.980 55.815 ;
        RECT 66.330 55.135 67.980 55.305 ;
        RECT 68.165 55.255 68.915 55.775 ;
        RECT 69.085 55.425 69.835 55.945 ;
        RECT 70.005 55.870 70.295 57.035 ;
        RECT 70.475 56.055 70.805 56.865 ;
        RECT 70.975 56.235 71.215 57.035 ;
        RECT 70.475 55.885 71.190 56.055 ;
        RECT 70.470 55.475 70.850 55.715 ;
        RECT 71.020 55.645 71.190 55.885 ;
        RECT 71.395 56.015 71.565 56.865 ;
        RECT 71.735 56.235 72.065 57.035 ;
        RECT 72.235 56.015 72.405 56.865 ;
        RECT 71.395 55.845 72.405 56.015 ;
        RECT 72.575 55.885 72.905 57.035 ;
        RECT 73.725 55.895 73.955 57.035 ;
        RECT 74.125 55.885 74.455 56.865 ;
        RECT 74.625 55.895 74.835 57.035 ;
        RECT 75.065 55.945 76.735 57.035 ;
        RECT 76.910 56.365 77.165 56.865 ;
        RECT 77.335 56.535 77.665 57.035 ;
        RECT 76.910 56.195 77.660 56.365 ;
        RECT 71.910 55.675 72.405 55.845 ;
        RECT 71.020 55.475 71.520 55.645 ;
        RECT 71.905 55.505 72.405 55.675 ;
        RECT 71.020 55.305 71.190 55.475 ;
        RECT 71.910 55.305 72.405 55.505 ;
        RECT 73.705 55.475 74.035 55.725 ;
        RECT 65.405 54.655 65.705 54.985 ;
        RECT 65.875 54.485 66.150 54.965 ;
        RECT 66.330 54.745 66.625 55.135 ;
        RECT 66.795 54.485 67.050 54.965 ;
        RECT 67.225 54.745 67.485 55.135 ;
        RECT 67.655 54.485 67.935 54.965 ;
        RECT 68.165 54.485 69.835 55.255 ;
        RECT 70.005 54.485 70.295 55.210 ;
        RECT 70.555 55.135 71.190 55.305 ;
        RECT 71.395 55.135 72.405 55.305 ;
        RECT 70.555 54.655 70.725 55.135 ;
        RECT 70.905 54.485 71.145 54.965 ;
        RECT 71.395 54.655 71.565 55.135 ;
        RECT 71.735 54.485 72.065 54.965 ;
        RECT 72.235 54.655 72.405 55.135 ;
        RECT 72.575 54.485 72.905 55.285 ;
        RECT 73.725 54.485 73.955 55.305 ;
        RECT 74.205 55.285 74.455 55.885 ;
        RECT 74.125 54.655 74.455 55.285 ;
        RECT 74.625 54.485 74.835 55.305 ;
        RECT 75.065 55.255 75.815 55.775 ;
        RECT 75.985 55.425 76.735 55.945 ;
        RECT 76.910 55.375 77.260 56.025 ;
        RECT 75.065 54.485 76.735 55.255 ;
        RECT 77.430 55.205 77.660 56.195 ;
        RECT 76.910 55.035 77.660 55.205 ;
        RECT 76.910 54.745 77.165 55.035 ;
        RECT 77.335 54.485 77.665 54.865 ;
        RECT 77.835 54.745 78.005 56.865 ;
        RECT 78.175 56.065 78.500 56.850 ;
        RECT 78.670 56.575 78.920 57.035 ;
        RECT 79.090 56.535 79.340 56.865 ;
        RECT 79.555 56.535 80.235 56.865 ;
        RECT 79.090 56.405 79.260 56.535 ;
        RECT 78.865 56.235 79.260 56.405 ;
        RECT 78.235 55.015 78.695 56.065 ;
        RECT 78.865 54.875 79.035 56.235 ;
        RECT 79.430 55.975 79.895 56.365 ;
        RECT 79.205 55.165 79.555 55.785 ;
        RECT 79.725 55.385 79.895 55.975 ;
        RECT 80.065 55.755 80.235 56.535 ;
        RECT 80.405 56.435 80.575 56.775 ;
        RECT 80.810 56.605 81.140 57.035 ;
        RECT 81.310 56.435 81.480 56.775 ;
        RECT 81.775 56.575 82.145 57.035 ;
        RECT 80.405 56.265 81.480 56.435 ;
        RECT 82.315 56.405 82.485 56.865 ;
        RECT 82.720 56.525 83.590 56.865 ;
        RECT 83.760 56.575 84.010 57.035 ;
        RECT 81.925 56.235 82.485 56.405 ;
        RECT 81.925 56.095 82.095 56.235 ;
        RECT 80.595 55.925 82.095 56.095 ;
        RECT 82.790 56.065 83.250 56.355 ;
        RECT 80.065 55.585 81.755 55.755 ;
        RECT 79.725 55.165 80.080 55.385 ;
        RECT 80.250 54.875 80.420 55.585 ;
        RECT 80.625 55.165 81.415 55.415 ;
        RECT 81.585 55.405 81.755 55.585 ;
        RECT 81.925 55.235 82.095 55.925 ;
        RECT 78.365 54.485 78.695 54.845 ;
        RECT 78.865 54.705 79.360 54.875 ;
        RECT 79.565 54.705 80.420 54.875 ;
        RECT 81.295 54.485 81.625 54.945 ;
        RECT 81.835 54.845 82.095 55.235 ;
        RECT 82.285 56.055 83.250 56.065 ;
        RECT 83.420 56.145 83.590 56.525 ;
        RECT 84.180 56.485 84.350 56.775 ;
        RECT 84.530 56.655 84.860 57.035 ;
        RECT 84.180 56.315 84.980 56.485 ;
        RECT 82.285 55.895 82.960 56.055 ;
        RECT 83.420 55.975 84.640 56.145 ;
        RECT 82.285 55.105 82.495 55.895 ;
        RECT 83.420 55.885 83.590 55.975 ;
        RECT 82.665 55.105 83.015 55.725 ;
        RECT 83.185 55.715 83.590 55.885 ;
        RECT 83.185 54.935 83.355 55.715 ;
        RECT 83.525 55.265 83.745 55.545 ;
        RECT 83.925 55.435 84.465 55.805 ;
        RECT 84.810 55.725 84.980 56.315 ;
        RECT 85.200 55.895 85.505 57.035 ;
        RECT 85.675 55.845 85.930 56.725 ;
        RECT 87.140 56.405 87.425 56.865 ;
        RECT 87.595 56.575 87.865 57.035 ;
        RECT 87.140 56.185 88.095 56.405 ;
        RECT 84.810 55.695 85.550 55.725 ;
        RECT 83.525 55.095 84.055 55.265 ;
        RECT 81.835 54.675 82.185 54.845 ;
        RECT 82.405 54.655 83.355 54.935 ;
        RECT 83.525 54.485 83.715 54.925 ;
        RECT 83.885 54.865 84.055 55.095 ;
        RECT 84.225 55.035 84.465 55.435 ;
        RECT 84.635 55.395 85.550 55.695 ;
        RECT 84.635 55.220 84.960 55.395 ;
        RECT 84.635 54.865 84.955 55.220 ;
        RECT 85.720 55.195 85.930 55.845 ;
        RECT 87.025 55.455 87.715 56.015 ;
        RECT 87.885 55.285 88.095 56.185 ;
        RECT 83.885 54.695 84.955 54.865 ;
        RECT 85.200 54.485 85.505 54.945 ;
        RECT 85.675 54.665 85.930 55.195 ;
        RECT 87.140 55.115 88.095 55.285 ;
        RECT 88.265 56.015 88.665 56.865 ;
        RECT 88.855 56.405 89.135 56.865 ;
        RECT 89.655 56.575 89.980 57.035 ;
        RECT 88.855 56.185 89.980 56.405 ;
        RECT 88.265 55.455 89.360 56.015 ;
        RECT 89.530 55.725 89.980 56.185 ;
        RECT 90.150 55.895 90.535 56.865 ;
        RECT 87.140 54.655 87.425 55.115 ;
        RECT 87.595 54.485 87.865 54.945 ;
        RECT 88.265 54.655 88.665 55.455 ;
        RECT 89.530 55.395 90.085 55.725 ;
        RECT 89.530 55.285 89.980 55.395 ;
        RECT 88.855 55.115 89.980 55.285 ;
        RECT 90.255 55.225 90.535 55.895 ;
        RECT 88.855 54.655 89.135 55.115 ;
        RECT 89.655 54.485 89.980 54.945 ;
        RECT 90.150 54.655 90.535 55.225 ;
        RECT 90.705 55.895 91.090 56.865 ;
        RECT 91.260 56.575 91.585 57.035 ;
        RECT 92.105 56.405 92.385 56.865 ;
        RECT 91.260 56.185 92.385 56.405 ;
        RECT 90.705 55.225 90.985 55.895 ;
        RECT 91.260 55.725 91.710 56.185 ;
        RECT 92.575 56.015 92.975 56.865 ;
        RECT 93.375 56.575 93.645 57.035 ;
        RECT 93.815 56.405 94.100 56.865 ;
        RECT 91.155 55.395 91.710 55.725 ;
        RECT 91.880 55.455 92.975 56.015 ;
        RECT 91.260 55.285 91.710 55.395 ;
        RECT 90.705 54.655 91.090 55.225 ;
        RECT 91.260 55.115 92.385 55.285 ;
        RECT 91.260 54.485 91.585 54.945 ;
        RECT 92.105 54.655 92.385 55.115 ;
        RECT 92.575 54.655 92.975 55.455 ;
        RECT 93.145 56.185 94.100 56.405 ;
        RECT 93.145 55.285 93.355 56.185 ;
        RECT 93.525 55.455 94.215 56.015 ;
        RECT 94.445 55.895 94.655 57.035 ;
        RECT 94.825 55.885 95.155 56.865 ;
        RECT 95.325 55.895 95.555 57.035 ;
        RECT 93.145 55.115 94.100 55.285 ;
        RECT 93.375 54.485 93.645 54.945 ;
        RECT 93.815 54.655 94.100 55.115 ;
        RECT 94.445 54.485 94.655 55.305 ;
        RECT 94.825 55.285 95.075 55.885 ;
        RECT 95.765 55.870 96.055 57.035 ;
        RECT 96.270 55.895 96.565 57.035 ;
        RECT 96.825 56.065 97.155 56.865 ;
        RECT 97.325 56.235 97.495 57.035 ;
        RECT 97.665 56.065 97.995 56.865 ;
        RECT 98.165 56.235 98.335 57.035 ;
        RECT 98.505 56.085 98.835 56.865 ;
        RECT 99.005 56.575 99.175 57.035 ;
        RECT 99.535 56.105 99.705 56.865 ;
        RECT 99.885 56.275 100.215 57.035 ;
        RECT 98.505 56.065 99.275 56.085 ;
        RECT 96.825 55.895 99.275 56.065 ;
        RECT 99.535 55.935 100.200 56.105 ;
        RECT 100.385 55.960 100.655 56.865 ;
        RECT 95.245 55.475 95.575 55.725 ;
        RECT 96.245 55.475 98.755 55.725 ;
        RECT 98.925 55.305 99.275 55.895 ;
        RECT 100.030 55.790 100.200 55.935 ;
        RECT 99.465 55.385 99.795 55.755 ;
        RECT 100.030 55.460 100.315 55.790 ;
        RECT 94.825 54.655 95.155 55.285 ;
        RECT 95.325 54.485 95.555 55.305 ;
        RECT 95.765 54.485 96.055 55.210 ;
        RECT 96.905 55.125 99.275 55.305 ;
        RECT 100.030 55.205 100.200 55.460 ;
        RECT 96.270 54.485 96.535 54.945 ;
        RECT 96.905 54.655 97.075 55.125 ;
        RECT 97.325 54.485 97.495 54.945 ;
        RECT 97.745 54.655 97.915 55.125 ;
        RECT 98.165 54.485 98.335 54.945 ;
        RECT 98.585 54.655 98.755 55.125 ;
        RECT 99.535 55.035 100.200 55.205 ;
        RECT 100.485 55.160 100.655 55.960 ;
        RECT 98.925 54.485 99.175 54.950 ;
        RECT 99.535 54.655 99.705 55.035 ;
        RECT 99.885 54.485 100.215 54.865 ;
        RECT 100.395 54.655 100.655 55.160 ;
        RECT 100.830 55.845 101.085 56.725 ;
        RECT 101.255 55.895 101.560 57.035 ;
        RECT 101.900 56.655 102.230 57.035 ;
        RECT 102.410 56.485 102.580 56.775 ;
        RECT 102.750 56.575 103.000 57.035 ;
        RECT 101.780 56.315 102.580 56.485 ;
        RECT 103.170 56.525 104.040 56.865 ;
        RECT 100.830 55.195 101.040 55.845 ;
        RECT 101.780 55.725 101.950 56.315 ;
        RECT 103.170 56.145 103.340 56.525 ;
        RECT 104.275 56.405 104.445 56.865 ;
        RECT 104.615 56.575 104.985 57.035 ;
        RECT 105.280 56.435 105.450 56.775 ;
        RECT 105.620 56.605 105.950 57.035 ;
        RECT 106.185 56.435 106.355 56.775 ;
        RECT 102.120 55.975 103.340 56.145 ;
        RECT 103.510 56.065 103.970 56.355 ;
        RECT 104.275 56.235 104.835 56.405 ;
        RECT 105.280 56.265 106.355 56.435 ;
        RECT 106.525 56.535 107.205 56.865 ;
        RECT 107.420 56.535 107.670 56.865 ;
        RECT 107.840 56.575 108.090 57.035 ;
        RECT 104.665 56.095 104.835 56.235 ;
        RECT 103.510 56.055 104.475 56.065 ;
        RECT 103.170 55.885 103.340 55.975 ;
        RECT 103.800 55.895 104.475 56.055 ;
        RECT 101.210 55.695 101.950 55.725 ;
        RECT 101.210 55.395 102.125 55.695 ;
        RECT 101.800 55.220 102.125 55.395 ;
        RECT 100.830 54.665 101.085 55.195 ;
        RECT 101.255 54.485 101.560 54.945 ;
        RECT 101.805 54.865 102.125 55.220 ;
        RECT 102.295 55.435 102.835 55.805 ;
        RECT 103.170 55.715 103.575 55.885 ;
        RECT 102.295 55.035 102.535 55.435 ;
        RECT 103.015 55.265 103.235 55.545 ;
        RECT 102.705 55.095 103.235 55.265 ;
        RECT 102.705 54.865 102.875 55.095 ;
        RECT 103.405 54.935 103.575 55.715 ;
        RECT 103.745 55.105 104.095 55.725 ;
        RECT 104.265 55.105 104.475 55.895 ;
        RECT 104.665 55.925 106.165 56.095 ;
        RECT 104.665 55.235 104.835 55.925 ;
        RECT 106.525 55.755 106.695 56.535 ;
        RECT 107.500 56.405 107.670 56.535 ;
        RECT 105.005 55.585 106.695 55.755 ;
        RECT 106.865 55.975 107.330 56.365 ;
        RECT 107.500 56.235 107.895 56.405 ;
        RECT 105.005 55.405 105.175 55.585 ;
        RECT 101.805 54.695 102.875 54.865 ;
        RECT 103.045 54.485 103.235 54.925 ;
        RECT 103.405 54.655 104.355 54.935 ;
        RECT 104.665 54.845 104.925 55.235 ;
        RECT 105.345 55.165 106.135 55.415 ;
        RECT 104.575 54.675 104.925 54.845 ;
        RECT 105.135 54.485 105.465 54.945 ;
        RECT 106.340 54.875 106.510 55.585 ;
        RECT 106.865 55.385 107.035 55.975 ;
        RECT 106.680 55.165 107.035 55.385 ;
        RECT 107.205 55.165 107.555 55.785 ;
        RECT 107.725 54.875 107.895 56.235 ;
        RECT 108.260 56.065 108.585 56.850 ;
        RECT 108.065 55.015 108.525 56.065 ;
        RECT 106.340 54.705 107.195 54.875 ;
        RECT 107.400 54.705 107.895 54.875 ;
        RECT 108.065 54.485 108.395 54.845 ;
        RECT 108.755 54.745 108.925 56.865 ;
        RECT 109.095 56.535 109.425 57.035 ;
        RECT 109.595 56.365 109.850 56.865 ;
        RECT 110.025 56.600 115.370 57.035 ;
        RECT 109.100 56.195 109.850 56.365 ;
        RECT 109.100 55.205 109.330 56.195 ;
        RECT 109.500 55.375 109.850 56.025 ;
        RECT 109.100 55.035 109.850 55.205 ;
        RECT 109.095 54.485 109.425 54.865 ;
        RECT 109.595 54.745 109.850 55.035 ;
        RECT 111.610 55.030 111.950 55.860 ;
        RECT 113.430 55.350 113.780 56.600 ;
        RECT 115.545 55.945 117.215 57.035 ;
        RECT 115.545 55.255 116.295 55.775 ;
        RECT 116.465 55.425 117.215 55.945 ;
        RECT 117.385 55.945 118.595 57.035 ;
        RECT 117.385 55.405 117.905 55.945 ;
        RECT 110.025 54.485 115.370 55.030 ;
        RECT 115.545 54.485 117.215 55.255 ;
        RECT 118.075 55.235 118.595 55.775 ;
        RECT 117.385 54.485 118.595 55.235 ;
        RECT 5.520 54.315 118.680 54.485 ;
        RECT 5.605 53.565 6.815 54.315 ;
        RECT 5.605 53.025 6.125 53.565 ;
        RECT 6.985 53.545 9.575 54.315 ;
        RECT 9.745 53.815 10.005 54.145 ;
        RECT 10.215 53.835 10.490 54.315 ;
        RECT 6.295 52.855 6.815 53.395 ;
        RECT 6.985 53.025 8.195 53.545 ;
        RECT 8.365 52.855 9.575 53.375 ;
        RECT 5.605 51.765 6.815 52.855 ;
        RECT 6.985 51.765 9.575 52.855 ;
        RECT 9.745 52.905 9.915 53.815 ;
        RECT 10.700 53.745 10.905 54.145 ;
        RECT 11.075 53.915 11.410 54.315 ;
        RECT 10.085 53.075 10.445 53.655 ;
        RECT 10.700 53.575 11.385 53.745 ;
        RECT 10.625 52.905 10.875 53.405 ;
        RECT 9.745 52.735 10.875 52.905 ;
        RECT 9.745 51.965 10.015 52.735 ;
        RECT 11.045 52.545 11.385 53.575 ;
        RECT 10.185 51.765 10.515 52.545 ;
        RECT 10.720 52.370 11.385 52.545 ;
        RECT 11.585 53.640 11.845 54.145 ;
        RECT 12.025 53.935 12.355 54.315 ;
        RECT 12.535 53.765 12.705 54.145 ;
        RECT 11.585 52.840 11.755 53.640 ;
        RECT 12.040 53.595 12.705 53.765 ;
        RECT 13.080 53.685 13.365 54.145 ;
        RECT 13.535 53.855 13.805 54.315 ;
        RECT 12.040 53.340 12.210 53.595 ;
        RECT 13.080 53.515 14.035 53.685 ;
        RECT 11.925 53.010 12.210 53.340 ;
        RECT 12.445 53.045 12.775 53.415 ;
        RECT 12.040 52.865 12.210 53.010 ;
        RECT 10.720 51.965 10.905 52.370 ;
        RECT 11.075 51.765 11.410 52.190 ;
        RECT 11.585 51.935 11.855 52.840 ;
        RECT 12.040 52.695 12.705 52.865 ;
        RECT 12.965 52.785 13.655 53.345 ;
        RECT 12.025 51.765 12.355 52.525 ;
        RECT 12.535 51.935 12.705 52.695 ;
        RECT 13.825 52.615 14.035 53.515 ;
        RECT 13.080 52.395 14.035 52.615 ;
        RECT 14.205 53.345 14.605 54.145 ;
        RECT 14.795 53.685 15.075 54.145 ;
        RECT 15.595 53.855 15.920 54.315 ;
        RECT 14.795 53.515 15.920 53.685 ;
        RECT 16.090 53.575 16.475 54.145 ;
        RECT 15.470 53.405 15.920 53.515 ;
        RECT 14.205 52.785 15.300 53.345 ;
        RECT 15.470 53.075 16.025 53.405 ;
        RECT 13.080 51.935 13.365 52.395 ;
        RECT 13.535 51.765 13.805 52.225 ;
        RECT 14.205 51.935 14.605 52.785 ;
        RECT 15.470 52.615 15.920 53.075 ;
        RECT 16.195 52.905 16.475 53.575 ;
        RECT 16.920 53.505 17.165 54.110 ;
        RECT 17.385 53.780 17.895 54.315 ;
        RECT 14.795 52.395 15.920 52.615 ;
        RECT 14.795 51.935 15.075 52.395 ;
        RECT 15.595 51.765 15.920 52.225 ;
        RECT 16.090 51.935 16.475 52.905 ;
        RECT 16.645 53.335 17.875 53.505 ;
        RECT 16.645 52.525 16.985 53.335 ;
        RECT 17.155 52.770 17.905 52.960 ;
        RECT 16.645 52.115 17.160 52.525 ;
        RECT 17.395 51.765 17.565 52.525 ;
        RECT 17.735 52.105 17.905 52.770 ;
        RECT 18.075 52.785 18.265 54.145 ;
        RECT 18.435 53.295 18.710 54.145 ;
        RECT 18.900 53.780 19.430 54.145 ;
        RECT 19.855 53.915 20.185 54.315 ;
        RECT 19.255 53.745 19.430 53.780 ;
        RECT 18.435 53.125 18.715 53.295 ;
        RECT 18.435 52.985 18.710 53.125 ;
        RECT 18.915 52.785 19.085 53.585 ;
        RECT 18.075 52.615 19.085 52.785 ;
        RECT 19.255 53.575 20.185 53.745 ;
        RECT 20.355 53.575 20.610 54.145 ;
        RECT 21.250 53.765 21.505 54.055 ;
        RECT 21.675 53.935 22.005 54.315 ;
        RECT 21.250 53.595 22.000 53.765 ;
        RECT 19.255 52.445 19.425 53.575 ;
        RECT 20.015 53.405 20.185 53.575 ;
        RECT 18.300 52.275 19.425 52.445 ;
        RECT 19.595 53.075 19.790 53.405 ;
        RECT 20.015 53.075 20.270 53.405 ;
        RECT 19.595 52.105 19.765 53.075 ;
        RECT 20.440 52.905 20.610 53.575 ;
        RECT 17.735 51.935 19.765 52.105 ;
        RECT 19.935 51.765 20.105 52.905 ;
        RECT 20.275 51.935 20.610 52.905 ;
        RECT 21.250 52.775 21.600 53.425 ;
        RECT 21.770 52.605 22.000 53.595 ;
        RECT 21.250 52.435 22.000 52.605 ;
        RECT 21.250 51.935 21.505 52.435 ;
        RECT 21.675 51.765 22.005 52.265 ;
        RECT 22.175 51.935 22.345 54.055 ;
        RECT 22.705 53.955 23.035 54.315 ;
        RECT 23.205 53.925 23.700 54.095 ;
        RECT 23.905 53.925 24.760 54.095 ;
        RECT 22.575 52.735 23.035 53.785 ;
        RECT 22.515 51.950 22.840 52.735 ;
        RECT 23.205 52.565 23.375 53.925 ;
        RECT 23.545 53.015 23.895 53.635 ;
        RECT 24.065 53.415 24.420 53.635 ;
        RECT 24.065 52.825 24.235 53.415 ;
        RECT 24.590 53.215 24.760 53.925 ;
        RECT 25.635 53.855 25.965 54.315 ;
        RECT 26.175 53.955 26.525 54.125 ;
        RECT 24.965 53.385 25.755 53.635 ;
        RECT 26.175 53.565 26.435 53.955 ;
        RECT 26.745 53.865 27.695 54.145 ;
        RECT 27.865 53.875 28.055 54.315 ;
        RECT 28.225 53.935 29.295 54.105 ;
        RECT 25.925 53.215 26.095 53.395 ;
        RECT 23.205 52.395 23.600 52.565 ;
        RECT 23.770 52.435 24.235 52.825 ;
        RECT 24.405 53.045 26.095 53.215 ;
        RECT 23.430 52.265 23.600 52.395 ;
        RECT 24.405 52.265 24.575 53.045 ;
        RECT 26.265 52.875 26.435 53.565 ;
        RECT 24.935 52.705 26.435 52.875 ;
        RECT 26.625 52.905 26.835 53.695 ;
        RECT 27.005 53.075 27.355 53.695 ;
        RECT 27.525 53.085 27.695 53.865 ;
        RECT 28.225 53.705 28.395 53.935 ;
        RECT 27.865 53.535 28.395 53.705 ;
        RECT 27.865 53.255 28.085 53.535 ;
        RECT 28.565 53.365 28.805 53.765 ;
        RECT 27.525 52.915 27.930 53.085 ;
        RECT 28.265 52.995 28.805 53.365 ;
        RECT 28.975 53.580 29.295 53.935 ;
        RECT 29.540 53.855 29.845 54.315 ;
        RECT 30.015 53.605 30.270 54.135 ;
        RECT 28.975 53.405 29.300 53.580 ;
        RECT 28.975 53.105 29.890 53.405 ;
        RECT 29.150 53.075 29.890 53.105 ;
        RECT 26.625 52.745 27.300 52.905 ;
        RECT 27.760 52.825 27.930 52.915 ;
        RECT 26.625 52.735 27.590 52.745 ;
        RECT 26.265 52.565 26.435 52.705 ;
        RECT 23.010 51.765 23.260 52.225 ;
        RECT 23.430 51.935 23.680 52.265 ;
        RECT 23.895 51.935 24.575 52.265 ;
        RECT 24.745 52.365 25.820 52.535 ;
        RECT 26.265 52.395 26.825 52.565 ;
        RECT 27.130 52.445 27.590 52.735 ;
        RECT 27.760 52.655 28.980 52.825 ;
        RECT 24.745 52.025 24.915 52.365 ;
        RECT 25.150 51.765 25.480 52.195 ;
        RECT 25.650 52.025 25.820 52.365 ;
        RECT 26.115 51.765 26.485 52.225 ;
        RECT 26.655 51.935 26.825 52.395 ;
        RECT 27.760 52.275 27.930 52.655 ;
        RECT 29.150 52.485 29.320 53.075 ;
        RECT 30.060 52.955 30.270 53.605 ;
        RECT 31.365 53.590 31.655 54.315 ;
        RECT 31.825 53.545 35.335 54.315 ;
        RECT 35.965 53.640 36.225 54.145 ;
        RECT 36.405 53.935 36.735 54.315 ;
        RECT 36.915 53.765 37.085 54.145 ;
        RECT 31.825 53.025 33.475 53.545 ;
        RECT 27.060 51.935 27.930 52.275 ;
        RECT 28.520 52.315 29.320 52.485 ;
        RECT 28.100 51.765 28.350 52.225 ;
        RECT 28.520 52.025 28.690 52.315 ;
        RECT 28.870 51.765 29.200 52.145 ;
        RECT 29.540 51.765 29.845 52.905 ;
        RECT 30.015 52.075 30.270 52.955 ;
        RECT 31.365 51.765 31.655 52.930 ;
        RECT 33.645 52.855 35.335 53.375 ;
        RECT 31.825 51.765 35.335 52.855 ;
        RECT 35.965 52.840 36.135 53.640 ;
        RECT 36.420 53.595 37.085 53.765 ;
        RECT 36.420 53.340 36.590 53.595 ;
        RECT 37.810 53.575 38.065 54.145 ;
        RECT 38.235 53.915 38.565 54.315 ;
        RECT 38.990 53.780 39.520 54.145 ;
        RECT 38.990 53.745 39.165 53.780 ;
        RECT 38.235 53.575 39.165 53.745 ;
        RECT 36.305 53.010 36.590 53.340 ;
        RECT 36.825 53.045 37.155 53.415 ;
        RECT 36.420 52.865 36.590 53.010 ;
        RECT 37.810 52.905 37.980 53.575 ;
        RECT 38.235 53.405 38.405 53.575 ;
        RECT 38.150 53.075 38.405 53.405 ;
        RECT 38.630 53.075 38.825 53.405 ;
        RECT 35.965 51.935 36.235 52.840 ;
        RECT 36.420 52.695 37.085 52.865 ;
        RECT 36.405 51.765 36.735 52.525 ;
        RECT 36.915 51.935 37.085 52.695 ;
        RECT 37.810 51.935 38.145 52.905 ;
        RECT 38.315 51.765 38.485 52.905 ;
        RECT 38.655 52.105 38.825 53.075 ;
        RECT 38.995 52.445 39.165 53.575 ;
        RECT 39.335 52.785 39.505 53.585 ;
        RECT 39.710 53.295 39.985 54.145 ;
        RECT 39.705 53.125 39.985 53.295 ;
        RECT 39.710 52.985 39.985 53.125 ;
        RECT 40.155 52.785 40.345 54.145 ;
        RECT 40.525 53.780 41.035 54.315 ;
        RECT 41.255 53.505 41.500 54.110 ;
        RECT 41.945 53.565 43.155 54.315 ;
        RECT 43.415 53.765 43.585 54.055 ;
        RECT 43.755 53.935 44.085 54.315 ;
        RECT 43.415 53.595 44.080 53.765 ;
        RECT 40.545 53.335 41.775 53.505 ;
        RECT 39.335 52.615 40.345 52.785 ;
        RECT 40.515 52.770 41.265 52.960 ;
        RECT 38.995 52.275 40.120 52.445 ;
        RECT 40.515 52.105 40.685 52.770 ;
        RECT 41.435 52.525 41.775 53.335 ;
        RECT 41.945 53.025 42.465 53.565 ;
        RECT 42.635 52.855 43.155 53.395 ;
        RECT 38.655 51.935 40.685 52.105 ;
        RECT 40.855 51.765 41.025 52.525 ;
        RECT 41.260 52.115 41.775 52.525 ;
        RECT 41.945 51.765 43.155 52.855 ;
        RECT 43.330 52.775 43.680 53.425 ;
        RECT 43.850 52.605 44.080 53.595 ;
        RECT 43.415 52.435 44.080 52.605 ;
        RECT 43.415 51.935 43.585 52.435 ;
        RECT 43.755 51.765 44.085 52.265 ;
        RECT 44.255 51.935 44.480 54.055 ;
        RECT 44.695 53.935 45.025 54.315 ;
        RECT 45.195 53.765 45.365 54.095 ;
        RECT 45.665 53.935 46.680 54.135 ;
        RECT 44.670 53.575 45.365 53.765 ;
        RECT 44.670 52.605 44.840 53.575 ;
        RECT 45.010 52.775 45.420 53.395 ;
        RECT 45.590 52.825 45.810 53.695 ;
        RECT 45.990 53.385 46.340 53.755 ;
        RECT 46.510 53.205 46.680 53.935 ;
        RECT 46.850 53.875 47.260 54.315 ;
        RECT 47.550 53.675 47.800 54.105 ;
        RECT 48.000 53.855 48.320 54.315 ;
        RECT 48.880 53.925 49.730 54.095 ;
        RECT 46.850 53.335 47.260 53.665 ;
        RECT 47.550 53.335 47.970 53.675 ;
        RECT 46.260 53.165 46.680 53.205 ;
        RECT 46.260 52.995 47.610 53.165 ;
        RECT 44.670 52.435 45.365 52.605 ;
        RECT 45.590 52.445 46.090 52.825 ;
        RECT 44.695 51.765 45.025 52.265 ;
        RECT 45.195 51.935 45.365 52.435 ;
        RECT 46.260 52.150 46.430 52.995 ;
        RECT 47.360 52.835 47.610 52.995 ;
        RECT 46.600 52.565 46.850 52.825 ;
        RECT 47.780 52.565 47.970 53.335 ;
        RECT 46.600 52.315 47.970 52.565 ;
        RECT 48.140 53.505 49.390 53.675 ;
        RECT 48.140 52.745 48.310 53.505 ;
        RECT 49.060 53.385 49.390 53.505 ;
        RECT 48.480 52.925 48.660 53.335 ;
        RECT 49.560 53.165 49.730 53.925 ;
        RECT 49.930 53.835 50.590 54.315 ;
        RECT 50.770 53.720 51.090 54.050 ;
        RECT 49.920 53.395 50.580 53.665 ;
        RECT 49.920 53.335 50.250 53.395 ;
        RECT 50.400 53.165 50.730 53.225 ;
        RECT 48.830 52.995 50.730 53.165 ;
        RECT 48.140 52.435 48.660 52.745 ;
        RECT 48.830 52.485 49.000 52.995 ;
        RECT 50.900 52.825 51.090 53.720 ;
        RECT 49.170 52.655 51.090 52.825 ;
        RECT 50.770 52.635 51.090 52.655 ;
        RECT 51.290 53.405 51.540 54.055 ;
        RECT 51.720 53.855 52.005 54.315 ;
        RECT 52.185 53.635 52.440 54.135 ;
        RECT 52.185 53.605 52.525 53.635 ;
        RECT 52.260 53.465 52.525 53.605 ;
        RECT 52.990 53.575 53.245 54.145 ;
        RECT 53.415 53.915 53.745 54.315 ;
        RECT 54.170 53.780 54.700 54.145 ;
        RECT 54.890 53.975 55.165 54.145 ;
        RECT 54.885 53.805 55.165 53.975 ;
        RECT 54.170 53.745 54.345 53.780 ;
        RECT 53.415 53.575 54.345 53.745 ;
        RECT 51.290 53.075 52.090 53.405 ;
        RECT 48.830 52.315 50.040 52.485 ;
        RECT 45.600 51.980 46.430 52.150 ;
        RECT 46.670 51.765 47.050 52.145 ;
        RECT 47.230 52.025 47.400 52.315 ;
        RECT 48.830 52.235 49.000 52.315 ;
        RECT 47.570 51.765 47.900 52.145 ;
        RECT 48.370 51.985 49.000 52.235 ;
        RECT 49.180 51.765 49.600 52.145 ;
        RECT 49.800 52.025 50.040 52.315 ;
        RECT 50.270 51.765 50.600 52.455 ;
        RECT 50.770 52.025 50.940 52.635 ;
        RECT 51.290 52.485 51.540 53.075 ;
        RECT 52.260 52.745 52.440 53.465 ;
        RECT 51.210 51.975 51.540 52.485 ;
        RECT 51.720 51.765 52.005 52.565 ;
        RECT 52.185 52.075 52.440 52.745 ;
        RECT 52.990 52.905 53.160 53.575 ;
        RECT 53.415 53.405 53.585 53.575 ;
        RECT 53.330 53.075 53.585 53.405 ;
        RECT 53.810 53.075 54.005 53.405 ;
        RECT 52.990 51.935 53.325 52.905 ;
        RECT 53.495 51.765 53.665 52.905 ;
        RECT 53.835 52.105 54.005 53.075 ;
        RECT 54.175 52.445 54.345 53.575 ;
        RECT 54.515 52.785 54.685 53.585 ;
        RECT 54.890 52.985 55.165 53.805 ;
        RECT 55.335 52.785 55.525 54.145 ;
        RECT 55.705 53.780 56.215 54.315 ;
        RECT 56.435 53.505 56.680 54.110 ;
        RECT 57.125 53.590 57.415 54.315 ;
        RECT 57.585 53.545 61.095 54.315 ;
        RECT 61.355 53.765 61.525 54.145 ;
        RECT 61.740 53.935 62.070 54.315 ;
        RECT 61.355 53.595 62.070 53.765 ;
        RECT 55.725 53.335 56.955 53.505 ;
        RECT 54.515 52.615 55.525 52.785 ;
        RECT 55.695 52.770 56.445 52.960 ;
        RECT 54.175 52.275 55.300 52.445 ;
        RECT 55.695 52.105 55.865 52.770 ;
        RECT 56.615 52.525 56.955 53.335 ;
        RECT 57.585 53.025 59.235 53.545 ;
        RECT 53.835 51.935 55.865 52.105 ;
        RECT 56.035 51.765 56.205 52.525 ;
        RECT 56.440 52.115 56.955 52.525 ;
        RECT 57.125 51.765 57.415 52.930 ;
        RECT 59.405 52.855 61.095 53.375 ;
        RECT 61.265 53.045 61.620 53.415 ;
        RECT 61.900 53.405 62.070 53.595 ;
        RECT 62.240 53.570 62.495 54.145 ;
        RECT 61.900 53.075 62.155 53.405 ;
        RECT 61.900 52.865 62.070 53.075 ;
        RECT 57.585 51.765 61.095 52.855 ;
        RECT 61.355 52.695 62.070 52.865 ;
        RECT 62.325 52.840 62.495 53.570 ;
        RECT 62.670 53.475 62.930 54.315 ;
        RECT 63.195 53.765 63.365 54.145 ;
        RECT 63.580 53.935 63.910 54.315 ;
        RECT 63.195 53.595 63.910 53.765 ;
        RECT 63.105 53.045 63.460 53.415 ;
        RECT 63.740 53.405 63.910 53.595 ;
        RECT 64.080 53.570 64.335 54.145 ;
        RECT 63.740 53.075 63.995 53.405 ;
        RECT 61.355 51.935 61.525 52.695 ;
        RECT 61.740 51.765 62.070 52.525 ;
        RECT 62.240 51.935 62.495 52.840 ;
        RECT 62.670 51.765 62.930 52.915 ;
        RECT 63.740 52.865 63.910 53.075 ;
        RECT 63.195 52.695 63.910 52.865 ;
        RECT 64.165 52.840 64.335 53.570 ;
        RECT 64.510 53.475 64.770 54.315 ;
        RECT 64.945 53.770 70.290 54.315 ;
        RECT 70.465 53.770 75.810 54.315 ;
        RECT 75.985 53.770 81.330 54.315 ;
        RECT 66.530 52.940 66.870 53.770 ;
        RECT 63.195 51.935 63.365 52.695 ;
        RECT 63.580 51.765 63.910 52.525 ;
        RECT 64.080 51.935 64.335 52.840 ;
        RECT 64.510 51.765 64.770 52.915 ;
        RECT 68.350 52.200 68.700 53.450 ;
        RECT 72.050 52.940 72.390 53.770 ;
        RECT 73.870 52.200 74.220 53.450 ;
        RECT 77.570 52.940 77.910 53.770 ;
        RECT 81.505 53.565 82.715 54.315 ;
        RECT 82.885 53.590 83.175 54.315 ;
        RECT 83.345 53.770 88.690 54.315 ;
        RECT 88.865 53.805 89.170 54.315 ;
        RECT 79.390 52.200 79.740 53.450 ;
        RECT 81.505 53.025 82.025 53.565 ;
        RECT 82.195 52.855 82.715 53.395 ;
        RECT 84.930 52.940 85.270 53.770 ;
        RECT 64.945 51.765 70.290 52.200 ;
        RECT 70.465 51.765 75.810 52.200 ;
        RECT 75.985 51.765 81.330 52.200 ;
        RECT 81.505 51.765 82.715 52.855 ;
        RECT 82.885 51.765 83.175 52.930 ;
        RECT 86.750 52.200 87.100 53.450 ;
        RECT 88.865 53.075 89.180 53.635 ;
        RECT 89.350 53.325 89.600 54.135 ;
        RECT 89.770 53.790 90.030 54.315 ;
        RECT 90.210 53.325 90.460 54.135 ;
        RECT 90.630 53.755 90.890 54.315 ;
        RECT 91.060 53.665 91.320 54.120 ;
        RECT 91.490 53.835 91.750 54.315 ;
        RECT 91.920 53.665 92.180 54.120 ;
        RECT 92.350 53.835 92.610 54.315 ;
        RECT 92.780 53.665 93.040 54.120 ;
        RECT 93.210 53.835 93.455 54.315 ;
        RECT 93.625 53.665 93.900 54.120 ;
        RECT 94.070 53.835 94.315 54.315 ;
        RECT 94.485 53.665 94.745 54.120 ;
        RECT 94.925 53.835 95.175 54.315 ;
        RECT 95.345 53.665 95.605 54.120 ;
        RECT 95.785 53.835 96.035 54.315 ;
        RECT 96.205 53.665 96.465 54.120 ;
        RECT 96.645 53.835 96.905 54.315 ;
        RECT 97.075 53.665 97.335 54.120 ;
        RECT 97.505 53.835 97.805 54.315 ;
        RECT 91.060 53.495 97.805 53.665 ;
        RECT 89.350 53.075 96.470 53.325 ;
        RECT 83.345 51.765 88.690 52.200 ;
        RECT 88.875 51.765 89.170 52.575 ;
        RECT 89.350 51.935 89.595 53.075 ;
        RECT 89.770 51.765 90.030 52.575 ;
        RECT 90.210 51.940 90.460 53.075 ;
        RECT 96.640 52.905 97.805 53.495 ;
        RECT 98.065 53.565 99.275 54.315 ;
        RECT 98.065 53.025 98.585 53.565 ;
        RECT 99.485 53.495 99.715 54.315 ;
        RECT 99.885 53.515 100.215 54.145 ;
        RECT 91.060 52.680 97.805 52.905 ;
        RECT 98.755 52.855 99.275 53.395 ;
        RECT 99.465 53.075 99.795 53.325 ;
        RECT 99.965 52.915 100.215 53.515 ;
        RECT 100.385 53.495 100.595 54.315 ;
        RECT 100.825 53.545 104.335 54.315 ;
        RECT 100.825 53.025 102.475 53.545 ;
        RECT 105.025 53.495 105.235 54.315 ;
        RECT 105.405 53.515 105.735 54.145 ;
        RECT 91.060 52.665 96.465 52.680 ;
        RECT 90.630 51.770 90.890 52.565 ;
        RECT 91.060 51.940 91.320 52.665 ;
        RECT 91.490 51.770 91.750 52.495 ;
        RECT 91.920 51.940 92.180 52.665 ;
        RECT 92.350 51.770 92.610 52.495 ;
        RECT 92.780 51.940 93.040 52.665 ;
        RECT 93.210 51.770 93.470 52.495 ;
        RECT 93.640 51.940 93.900 52.665 ;
        RECT 94.070 51.770 94.315 52.495 ;
        RECT 94.485 51.940 94.745 52.665 ;
        RECT 94.930 51.770 95.175 52.495 ;
        RECT 95.345 51.940 95.605 52.665 ;
        RECT 95.790 51.770 96.035 52.495 ;
        RECT 96.205 51.940 96.465 52.665 ;
        RECT 96.650 51.770 96.905 52.495 ;
        RECT 97.075 51.940 97.365 52.680 ;
        RECT 90.630 51.765 96.905 51.770 ;
        RECT 97.535 51.765 97.805 52.510 ;
        RECT 98.065 51.765 99.275 52.855 ;
        RECT 99.485 51.765 99.715 52.905 ;
        RECT 99.885 51.935 100.215 52.915 ;
        RECT 100.385 51.765 100.595 52.905 ;
        RECT 102.645 52.855 104.335 53.375 ;
        RECT 105.405 52.915 105.655 53.515 ;
        RECT 105.905 53.495 106.135 54.315 ;
        RECT 106.345 53.545 108.015 54.315 ;
        RECT 108.645 53.590 108.935 54.315 ;
        RECT 109.105 53.770 114.450 54.315 ;
        RECT 105.825 53.075 106.155 53.325 ;
        RECT 106.345 53.025 107.095 53.545 ;
        RECT 100.825 51.765 104.335 52.855 ;
        RECT 105.025 51.765 105.235 52.905 ;
        RECT 105.405 51.935 105.735 52.915 ;
        RECT 105.905 51.765 106.135 52.905 ;
        RECT 107.265 52.855 108.015 53.375 ;
        RECT 110.690 52.940 111.030 53.770 ;
        RECT 114.625 53.545 117.215 54.315 ;
        RECT 117.385 53.565 118.595 54.315 ;
        RECT 106.345 51.765 108.015 52.855 ;
        RECT 108.645 51.765 108.935 52.930 ;
        RECT 112.510 52.200 112.860 53.450 ;
        RECT 114.625 53.025 115.835 53.545 ;
        RECT 116.005 52.855 117.215 53.375 ;
        RECT 109.105 51.765 114.450 52.200 ;
        RECT 114.625 51.765 117.215 52.855 ;
        RECT 117.385 52.855 117.905 53.395 ;
        RECT 118.075 53.025 118.595 53.565 ;
        RECT 117.385 51.765 118.595 52.855 ;
        RECT 5.520 51.595 118.680 51.765 ;
        RECT 5.605 50.505 6.815 51.595 ;
        RECT 6.985 50.505 8.195 51.595 ;
        RECT 8.370 50.925 8.625 51.425 ;
        RECT 8.795 51.095 9.125 51.595 ;
        RECT 8.370 50.755 9.120 50.925 ;
        RECT 5.605 49.795 6.125 50.335 ;
        RECT 6.295 49.965 6.815 50.505 ;
        RECT 6.985 49.795 7.505 50.335 ;
        RECT 7.675 49.965 8.195 50.505 ;
        RECT 8.370 49.935 8.720 50.585 ;
        RECT 5.605 49.045 6.815 49.795 ;
        RECT 6.985 49.045 8.195 49.795 ;
        RECT 8.890 49.765 9.120 50.755 ;
        RECT 8.370 49.595 9.120 49.765 ;
        RECT 8.370 49.305 8.625 49.595 ;
        RECT 8.795 49.045 9.125 49.425 ;
        RECT 9.295 49.305 9.465 51.425 ;
        RECT 9.635 50.625 9.960 51.410 ;
        RECT 10.130 51.135 10.380 51.595 ;
        RECT 10.550 51.095 10.800 51.425 ;
        RECT 11.015 51.095 11.695 51.425 ;
        RECT 10.550 50.965 10.720 51.095 ;
        RECT 10.325 50.795 10.720 50.965 ;
        RECT 9.695 49.575 10.155 50.625 ;
        RECT 10.325 49.435 10.495 50.795 ;
        RECT 10.890 50.535 11.355 50.925 ;
        RECT 10.665 49.725 11.015 50.345 ;
        RECT 11.185 49.945 11.355 50.535 ;
        RECT 11.525 50.315 11.695 51.095 ;
        RECT 11.865 50.995 12.035 51.335 ;
        RECT 12.270 51.165 12.600 51.595 ;
        RECT 12.770 50.995 12.940 51.335 ;
        RECT 13.235 51.135 13.605 51.595 ;
        RECT 11.865 50.825 12.940 50.995 ;
        RECT 13.775 50.965 13.945 51.425 ;
        RECT 14.180 51.085 15.050 51.425 ;
        RECT 15.220 51.135 15.470 51.595 ;
        RECT 13.385 50.795 13.945 50.965 ;
        RECT 13.385 50.655 13.555 50.795 ;
        RECT 12.055 50.485 13.555 50.655 ;
        RECT 14.250 50.625 14.710 50.915 ;
        RECT 11.525 50.145 13.215 50.315 ;
        RECT 11.185 49.725 11.540 49.945 ;
        RECT 11.710 49.435 11.880 50.145 ;
        RECT 12.085 49.725 12.875 49.975 ;
        RECT 13.045 49.965 13.215 50.145 ;
        RECT 13.385 49.795 13.555 50.485 ;
        RECT 9.825 49.045 10.155 49.405 ;
        RECT 10.325 49.265 10.820 49.435 ;
        RECT 11.025 49.265 11.880 49.435 ;
        RECT 12.755 49.045 13.085 49.505 ;
        RECT 13.295 49.405 13.555 49.795 ;
        RECT 13.745 50.615 14.710 50.625 ;
        RECT 14.880 50.705 15.050 51.085 ;
        RECT 15.640 51.045 15.810 51.335 ;
        RECT 15.990 51.215 16.320 51.595 ;
        RECT 15.640 50.875 16.440 51.045 ;
        RECT 13.745 50.455 14.420 50.615 ;
        RECT 14.880 50.535 16.100 50.705 ;
        RECT 13.745 49.665 13.955 50.455 ;
        RECT 14.880 50.445 15.050 50.535 ;
        RECT 14.125 49.665 14.475 50.285 ;
        RECT 14.645 50.275 15.050 50.445 ;
        RECT 14.645 49.495 14.815 50.275 ;
        RECT 14.985 49.825 15.205 50.105 ;
        RECT 15.385 49.995 15.925 50.365 ;
        RECT 16.270 50.285 16.440 50.875 ;
        RECT 16.660 50.455 16.965 51.595 ;
        RECT 17.135 50.405 17.390 51.285 ;
        RECT 18.485 50.430 18.775 51.595 ;
        RECT 19.005 50.455 19.215 51.595 ;
        RECT 19.385 50.445 19.715 51.425 ;
        RECT 19.885 50.455 20.115 51.595 ;
        RECT 20.325 50.505 21.535 51.595 ;
        RECT 16.270 50.255 17.010 50.285 ;
        RECT 14.985 49.655 15.515 49.825 ;
        RECT 13.295 49.235 13.645 49.405 ;
        RECT 13.865 49.215 14.815 49.495 ;
        RECT 14.985 49.045 15.175 49.485 ;
        RECT 15.345 49.425 15.515 49.655 ;
        RECT 15.685 49.595 15.925 49.995 ;
        RECT 16.095 49.955 17.010 50.255 ;
        RECT 16.095 49.780 16.420 49.955 ;
        RECT 16.095 49.425 16.415 49.780 ;
        RECT 17.180 49.755 17.390 50.405 ;
        RECT 15.345 49.255 16.415 49.425 ;
        RECT 16.660 49.045 16.965 49.505 ;
        RECT 17.135 49.225 17.390 49.755 ;
        RECT 18.485 49.045 18.775 49.770 ;
        RECT 19.005 49.045 19.215 49.865 ;
        RECT 19.385 49.845 19.635 50.445 ;
        RECT 19.805 50.035 20.135 50.285 ;
        RECT 19.385 49.215 19.715 49.845 ;
        RECT 19.885 49.045 20.115 49.865 ;
        RECT 20.325 49.795 20.845 50.335 ;
        RECT 21.015 49.965 21.535 50.505 ;
        RECT 21.705 50.455 22.045 51.425 ;
        RECT 22.215 50.455 22.385 51.595 ;
        RECT 22.655 50.795 22.905 51.595 ;
        RECT 23.550 50.625 23.880 51.425 ;
        RECT 24.180 50.795 24.510 51.595 ;
        RECT 24.680 50.625 25.010 51.425 ;
        RECT 22.575 50.455 25.010 50.625 ;
        RECT 25.425 50.455 25.655 51.595 ;
        RECT 21.705 49.845 21.880 50.455 ;
        RECT 22.575 50.205 22.745 50.455 ;
        RECT 22.050 50.035 22.745 50.205 ;
        RECT 22.920 50.035 23.340 50.235 ;
        RECT 23.510 50.035 23.840 50.235 ;
        RECT 24.010 50.035 24.340 50.235 ;
        RECT 20.325 49.045 21.535 49.795 ;
        RECT 21.705 49.215 22.045 49.845 ;
        RECT 22.215 49.045 22.465 49.845 ;
        RECT 22.655 49.695 23.880 49.865 ;
        RECT 22.655 49.215 22.985 49.695 ;
        RECT 23.155 49.045 23.380 49.505 ;
        RECT 23.550 49.215 23.880 49.695 ;
        RECT 24.510 49.825 24.680 50.455 ;
        RECT 25.825 50.445 26.155 51.425 ;
        RECT 26.325 50.455 26.535 51.595 ;
        RECT 26.765 51.160 32.110 51.595 ;
        RECT 24.865 50.035 25.215 50.285 ;
        RECT 25.405 50.035 25.735 50.285 ;
        RECT 24.510 49.215 25.010 49.825 ;
        RECT 25.425 49.045 25.655 49.865 ;
        RECT 25.905 49.845 26.155 50.445 ;
        RECT 25.825 49.215 26.155 49.845 ;
        RECT 26.325 49.045 26.535 49.865 ;
        RECT 28.350 49.590 28.690 50.420 ;
        RECT 30.170 49.910 30.520 51.160 ;
        RECT 33.210 50.925 33.465 51.425 ;
        RECT 33.635 51.095 33.965 51.595 ;
        RECT 33.210 50.755 33.960 50.925 ;
        RECT 33.210 49.935 33.560 50.585 ;
        RECT 33.730 49.765 33.960 50.755 ;
        RECT 33.210 49.595 33.960 49.765 ;
        RECT 26.765 49.045 32.110 49.590 ;
        RECT 33.210 49.305 33.465 49.595 ;
        RECT 33.635 49.045 33.965 49.425 ;
        RECT 34.135 49.305 34.305 51.425 ;
        RECT 34.475 50.625 34.800 51.410 ;
        RECT 34.970 51.135 35.220 51.595 ;
        RECT 35.390 51.095 35.640 51.425 ;
        RECT 35.855 51.095 36.535 51.425 ;
        RECT 35.390 50.965 35.560 51.095 ;
        RECT 35.165 50.795 35.560 50.965 ;
        RECT 34.535 49.575 34.995 50.625 ;
        RECT 35.165 49.435 35.335 50.795 ;
        RECT 35.730 50.535 36.195 50.925 ;
        RECT 35.505 49.725 35.855 50.345 ;
        RECT 36.025 49.945 36.195 50.535 ;
        RECT 36.365 50.315 36.535 51.095 ;
        RECT 36.705 50.995 36.875 51.335 ;
        RECT 37.110 51.165 37.440 51.595 ;
        RECT 37.610 50.995 37.780 51.335 ;
        RECT 38.075 51.135 38.445 51.595 ;
        RECT 36.705 50.825 37.780 50.995 ;
        RECT 38.615 50.965 38.785 51.425 ;
        RECT 39.020 51.085 39.890 51.425 ;
        RECT 40.060 51.135 40.310 51.595 ;
        RECT 38.225 50.795 38.785 50.965 ;
        RECT 38.225 50.655 38.395 50.795 ;
        RECT 36.895 50.485 38.395 50.655 ;
        RECT 39.090 50.625 39.550 50.915 ;
        RECT 36.365 50.145 38.055 50.315 ;
        RECT 36.025 49.725 36.380 49.945 ;
        RECT 36.550 49.435 36.720 50.145 ;
        RECT 36.925 49.725 37.715 49.975 ;
        RECT 37.885 49.965 38.055 50.145 ;
        RECT 38.225 49.795 38.395 50.485 ;
        RECT 34.665 49.045 34.995 49.405 ;
        RECT 35.165 49.265 35.660 49.435 ;
        RECT 35.865 49.265 36.720 49.435 ;
        RECT 37.595 49.045 37.925 49.505 ;
        RECT 38.135 49.405 38.395 49.795 ;
        RECT 38.585 50.615 39.550 50.625 ;
        RECT 39.720 50.705 39.890 51.085 ;
        RECT 40.480 51.045 40.650 51.335 ;
        RECT 40.830 51.215 41.160 51.595 ;
        RECT 40.480 50.875 41.280 51.045 ;
        RECT 38.585 50.455 39.260 50.615 ;
        RECT 39.720 50.535 40.940 50.705 ;
        RECT 38.585 49.665 38.795 50.455 ;
        RECT 39.720 50.445 39.890 50.535 ;
        RECT 38.965 49.665 39.315 50.285 ;
        RECT 39.485 50.275 39.890 50.445 ;
        RECT 39.485 49.495 39.655 50.275 ;
        RECT 39.825 49.825 40.045 50.105 ;
        RECT 40.225 49.995 40.765 50.365 ;
        RECT 41.110 50.285 41.280 50.875 ;
        RECT 41.500 50.455 41.805 51.595 ;
        RECT 41.975 50.405 42.230 51.285 ;
        RECT 42.465 50.455 42.675 51.595 ;
        RECT 41.110 50.255 41.850 50.285 ;
        RECT 39.825 49.655 40.355 49.825 ;
        RECT 38.135 49.235 38.485 49.405 ;
        RECT 38.705 49.215 39.655 49.495 ;
        RECT 39.825 49.045 40.015 49.485 ;
        RECT 40.185 49.425 40.355 49.655 ;
        RECT 40.525 49.595 40.765 49.995 ;
        RECT 40.935 49.955 41.850 50.255 ;
        RECT 40.935 49.780 41.260 49.955 ;
        RECT 40.935 49.425 41.255 49.780 ;
        RECT 42.020 49.755 42.230 50.405 ;
        RECT 42.845 50.445 43.175 51.425 ;
        RECT 43.345 50.455 43.575 51.595 ;
        RECT 40.185 49.255 41.255 49.425 ;
        RECT 41.500 49.045 41.805 49.505 ;
        RECT 41.975 49.225 42.230 49.755 ;
        RECT 42.465 49.045 42.675 49.865 ;
        RECT 42.845 49.845 43.095 50.445 ;
        RECT 44.245 50.430 44.535 51.595 ;
        RECT 44.705 50.455 45.090 51.425 ;
        RECT 45.260 51.135 45.585 51.595 ;
        RECT 46.105 50.965 46.385 51.425 ;
        RECT 45.260 50.745 46.385 50.965 ;
        RECT 43.265 50.035 43.595 50.285 ;
        RECT 42.845 49.215 43.175 49.845 ;
        RECT 43.345 49.045 43.575 49.865 ;
        RECT 44.705 49.785 44.985 50.455 ;
        RECT 45.260 50.285 45.710 50.745 ;
        RECT 46.575 50.575 46.975 51.425 ;
        RECT 47.375 51.135 47.645 51.595 ;
        RECT 47.815 50.965 48.100 51.425 ;
        RECT 45.155 49.955 45.710 50.285 ;
        RECT 45.880 50.015 46.975 50.575 ;
        RECT 45.260 49.845 45.710 49.955 ;
        RECT 44.245 49.045 44.535 49.770 ;
        RECT 44.705 49.215 45.090 49.785 ;
        RECT 45.260 49.675 46.385 49.845 ;
        RECT 45.260 49.045 45.585 49.505 ;
        RECT 46.105 49.215 46.385 49.675 ;
        RECT 46.575 49.215 46.975 50.015 ;
        RECT 47.145 50.745 48.100 50.965 ;
        RECT 47.145 49.845 47.355 50.745 ;
        RECT 47.525 50.015 48.215 50.575 ;
        RECT 48.535 50.445 48.865 51.595 ;
        RECT 49.035 50.575 49.205 51.425 ;
        RECT 49.375 50.795 49.705 51.595 ;
        RECT 49.875 50.575 50.045 51.425 ;
        RECT 50.225 50.795 50.465 51.595 ;
        RECT 50.635 50.615 50.965 51.425 ;
        RECT 51.145 51.160 56.490 51.595 ;
        RECT 56.665 51.160 62.010 51.595 ;
        RECT 62.185 51.160 67.530 51.595 ;
        RECT 49.035 50.405 50.045 50.575 ;
        RECT 50.250 50.445 50.965 50.615 ;
        RECT 49.035 49.895 49.530 50.405 ;
        RECT 50.250 50.205 50.420 50.445 ;
        RECT 49.920 50.035 50.420 50.205 ;
        RECT 50.590 50.035 50.970 50.275 ;
        RECT 49.035 49.865 49.535 49.895 ;
        RECT 50.250 49.865 50.420 50.035 ;
        RECT 47.145 49.675 48.100 49.845 ;
        RECT 47.375 49.045 47.645 49.505 ;
        RECT 47.815 49.215 48.100 49.675 ;
        RECT 48.535 49.045 48.865 49.845 ;
        RECT 49.035 49.695 50.045 49.865 ;
        RECT 50.250 49.695 50.885 49.865 ;
        RECT 49.035 49.215 49.205 49.695 ;
        RECT 49.375 49.045 49.705 49.525 ;
        RECT 49.875 49.215 50.045 49.695 ;
        RECT 50.295 49.045 50.535 49.525 ;
        RECT 50.715 49.215 50.885 49.695 ;
        RECT 52.730 49.590 53.070 50.420 ;
        RECT 54.550 49.910 54.900 51.160 ;
        RECT 58.250 49.590 58.590 50.420 ;
        RECT 60.070 49.910 60.420 51.160 ;
        RECT 63.770 49.590 64.110 50.420 ;
        RECT 65.590 49.910 65.940 51.160 ;
        RECT 67.705 50.505 69.375 51.595 ;
        RECT 67.705 49.815 68.455 50.335 ;
        RECT 68.625 49.985 69.375 50.505 ;
        RECT 70.005 50.430 70.295 51.595 ;
        RECT 70.465 50.520 70.735 51.425 ;
        RECT 70.905 50.835 71.235 51.595 ;
        RECT 71.415 50.665 71.585 51.425 ;
        RECT 51.145 49.045 56.490 49.590 ;
        RECT 56.665 49.045 62.010 49.590 ;
        RECT 62.185 49.045 67.530 49.590 ;
        RECT 67.705 49.045 69.375 49.815 ;
        RECT 70.005 49.045 70.295 49.770 ;
        RECT 70.465 49.720 70.635 50.520 ;
        RECT 70.920 50.495 71.585 50.665 ;
        RECT 70.920 50.350 71.090 50.495 ;
        RECT 71.885 50.455 72.115 51.595 ;
        RECT 72.285 50.445 72.615 51.425 ;
        RECT 72.785 50.455 72.995 51.595 ;
        RECT 73.225 50.505 76.735 51.595 ;
        RECT 76.905 50.505 78.115 51.595 ;
        RECT 70.805 50.020 71.090 50.350 ;
        RECT 70.920 49.765 71.090 50.020 ;
        RECT 71.325 49.945 71.655 50.315 ;
        RECT 71.865 50.035 72.195 50.285 ;
        RECT 70.465 49.215 70.725 49.720 ;
        RECT 70.920 49.595 71.585 49.765 ;
        RECT 70.905 49.045 71.235 49.425 ;
        RECT 71.415 49.215 71.585 49.595 ;
        RECT 71.885 49.045 72.115 49.865 ;
        RECT 72.365 49.845 72.615 50.445 ;
        RECT 72.285 49.215 72.615 49.845 ;
        RECT 72.785 49.045 72.995 49.865 ;
        RECT 73.225 49.815 74.875 50.335 ;
        RECT 75.045 49.985 76.735 50.505 ;
        RECT 73.225 49.045 76.735 49.815 ;
        RECT 76.905 49.795 77.425 50.335 ;
        RECT 77.595 49.965 78.115 50.505 ;
        RECT 78.490 50.625 78.820 51.425 ;
        RECT 78.990 50.795 79.320 51.595 ;
        RECT 79.620 50.625 79.950 51.425 ;
        RECT 80.595 50.795 80.845 51.595 ;
        RECT 78.490 50.455 80.925 50.625 ;
        RECT 81.115 50.455 81.285 51.595 ;
        RECT 81.455 50.455 81.795 51.425 ;
        RECT 82.170 50.625 82.500 51.425 ;
        RECT 82.670 50.795 83.000 51.595 ;
        RECT 83.300 50.625 83.630 51.425 ;
        RECT 84.275 50.795 84.525 51.595 ;
        RECT 82.170 50.455 84.605 50.625 ;
        RECT 84.795 50.455 84.965 51.595 ;
        RECT 85.135 50.455 85.475 51.425 ;
        RECT 85.850 50.625 86.180 51.425 ;
        RECT 86.350 50.795 86.680 51.595 ;
        RECT 86.980 50.625 87.310 51.425 ;
        RECT 87.955 50.795 88.205 51.595 ;
        RECT 85.850 50.455 88.285 50.625 ;
        RECT 88.475 50.455 88.645 51.595 ;
        RECT 88.815 50.455 89.155 51.425 ;
        RECT 90.335 50.665 90.505 51.425 ;
        RECT 90.685 50.835 91.015 51.595 ;
        RECT 90.335 50.495 91.000 50.665 ;
        RECT 91.185 50.520 91.455 51.425 ;
        RECT 78.285 50.035 78.635 50.285 ;
        RECT 78.820 49.825 78.990 50.455 ;
        RECT 79.160 50.035 79.490 50.235 ;
        RECT 79.660 50.035 79.990 50.235 ;
        RECT 80.160 50.035 80.580 50.235 ;
        RECT 80.755 50.205 80.925 50.455 ;
        RECT 80.755 50.035 81.450 50.205 ;
        RECT 76.905 49.045 78.115 49.795 ;
        RECT 78.490 49.215 78.990 49.825 ;
        RECT 79.620 49.695 80.845 49.865 ;
        RECT 81.620 49.845 81.795 50.455 ;
        RECT 81.965 50.035 82.315 50.285 ;
        RECT 79.620 49.215 79.950 49.695 ;
        RECT 80.120 49.045 80.345 49.505 ;
        RECT 80.515 49.215 80.845 49.695 ;
        RECT 81.035 49.045 81.285 49.845 ;
        RECT 81.455 49.215 81.795 49.845 ;
        RECT 82.500 49.825 82.670 50.455 ;
        RECT 82.840 50.035 83.170 50.235 ;
        RECT 83.340 50.035 83.670 50.235 ;
        RECT 83.840 50.035 84.260 50.235 ;
        RECT 84.435 50.205 84.605 50.455 ;
        RECT 84.435 50.035 85.130 50.205 ;
        RECT 82.170 49.215 82.670 49.825 ;
        RECT 83.300 49.695 84.525 49.865 ;
        RECT 85.300 49.845 85.475 50.455 ;
        RECT 85.645 50.035 85.995 50.285 ;
        RECT 83.300 49.215 83.630 49.695 ;
        RECT 83.800 49.045 84.025 49.505 ;
        RECT 84.195 49.215 84.525 49.695 ;
        RECT 84.715 49.045 84.965 49.845 ;
        RECT 85.135 49.215 85.475 49.845 ;
        RECT 86.180 49.825 86.350 50.455 ;
        RECT 86.520 50.035 86.850 50.235 ;
        RECT 87.020 50.035 87.350 50.235 ;
        RECT 87.520 50.035 87.940 50.235 ;
        RECT 88.115 50.205 88.285 50.455 ;
        RECT 88.115 50.035 88.810 50.205 ;
        RECT 85.850 49.215 86.350 49.825 ;
        RECT 86.980 49.695 88.205 49.865 ;
        RECT 88.980 49.845 89.155 50.455 ;
        RECT 90.830 50.350 91.000 50.495 ;
        RECT 90.265 49.945 90.595 50.315 ;
        RECT 90.830 50.020 91.115 50.350 ;
        RECT 86.980 49.215 87.310 49.695 ;
        RECT 87.480 49.045 87.705 49.505 ;
        RECT 87.875 49.215 88.205 49.695 ;
        RECT 88.395 49.045 88.645 49.845 ;
        RECT 88.815 49.215 89.155 49.845 ;
        RECT 90.830 49.765 91.000 50.020 ;
        RECT 90.335 49.595 91.000 49.765 ;
        RECT 91.285 49.720 91.455 50.520 ;
        RECT 92.290 50.625 92.620 51.425 ;
        RECT 92.790 50.795 93.120 51.595 ;
        RECT 93.420 50.625 93.750 51.425 ;
        RECT 94.395 50.795 94.645 51.595 ;
        RECT 92.290 50.455 94.725 50.625 ;
        RECT 94.915 50.455 95.085 51.595 ;
        RECT 95.255 50.455 95.595 51.425 ;
        RECT 92.085 50.035 92.435 50.285 ;
        RECT 92.620 49.825 92.790 50.455 ;
        RECT 92.960 50.035 93.290 50.235 ;
        RECT 93.460 50.035 93.790 50.235 ;
        RECT 93.960 50.035 94.380 50.235 ;
        RECT 94.555 50.205 94.725 50.455 ;
        RECT 94.555 50.035 95.250 50.205 ;
        RECT 90.335 49.215 90.505 49.595 ;
        RECT 90.685 49.045 91.015 49.425 ;
        RECT 91.195 49.215 91.455 49.720 ;
        RECT 92.290 49.215 92.790 49.825 ;
        RECT 93.420 49.695 94.645 49.865 ;
        RECT 95.420 49.845 95.595 50.455 ;
        RECT 95.765 50.430 96.055 51.595 ;
        RECT 96.225 51.160 101.570 51.595 ;
        RECT 101.745 51.160 107.090 51.595 ;
        RECT 107.265 51.160 112.610 51.595 ;
        RECT 93.420 49.215 93.750 49.695 ;
        RECT 93.920 49.045 94.145 49.505 ;
        RECT 94.315 49.215 94.645 49.695 ;
        RECT 94.835 49.045 95.085 49.845 ;
        RECT 95.255 49.215 95.595 49.845 ;
        RECT 95.765 49.045 96.055 49.770 ;
        RECT 97.810 49.590 98.150 50.420 ;
        RECT 99.630 49.910 99.980 51.160 ;
        RECT 103.330 49.590 103.670 50.420 ;
        RECT 105.150 49.910 105.500 51.160 ;
        RECT 108.850 49.590 109.190 50.420 ;
        RECT 110.670 49.910 111.020 51.160 ;
        RECT 112.785 50.505 116.295 51.595 ;
        RECT 112.785 49.815 114.435 50.335 ;
        RECT 114.605 49.985 116.295 50.505 ;
        RECT 117.385 50.505 118.595 51.595 ;
        RECT 117.385 49.965 117.905 50.505 ;
        RECT 96.225 49.045 101.570 49.590 ;
        RECT 101.745 49.045 107.090 49.590 ;
        RECT 107.265 49.045 112.610 49.590 ;
        RECT 112.785 49.045 116.295 49.815 ;
        RECT 118.075 49.795 118.595 50.335 ;
        RECT 117.385 49.045 118.595 49.795 ;
        RECT 5.520 48.875 118.680 49.045 ;
        RECT 5.605 48.125 6.815 48.875 ;
        RECT 6.985 48.330 12.330 48.875 ;
        RECT 5.605 47.585 6.125 48.125 ;
        RECT 6.295 47.415 6.815 47.955 ;
        RECT 8.570 47.500 8.910 48.330 ;
        RECT 12.505 48.125 13.715 48.875 ;
        RECT 5.605 46.325 6.815 47.415 ;
        RECT 10.390 46.760 10.740 48.010 ;
        RECT 12.505 47.585 13.025 48.125 ;
        RECT 13.945 48.055 14.155 48.875 ;
        RECT 14.325 48.075 14.655 48.705 ;
        RECT 13.195 47.415 13.715 47.955 ;
        RECT 14.325 47.475 14.575 48.075 ;
        RECT 14.825 48.055 15.055 48.875 ;
        RECT 15.265 48.330 20.610 48.875 ;
        RECT 14.745 47.635 15.075 47.885 ;
        RECT 16.850 47.500 17.190 48.330 ;
        RECT 20.785 48.125 21.995 48.875 ;
        RECT 6.985 46.325 12.330 46.760 ;
        RECT 12.505 46.325 13.715 47.415 ;
        RECT 13.945 46.325 14.155 47.465 ;
        RECT 14.325 46.495 14.655 47.475 ;
        RECT 14.825 46.325 15.055 47.465 ;
        RECT 18.670 46.760 19.020 48.010 ;
        RECT 20.785 47.585 21.305 48.125 ;
        RECT 22.370 48.095 22.870 48.705 ;
        RECT 21.475 47.415 21.995 47.955 ;
        RECT 22.165 47.635 22.515 47.885 ;
        RECT 22.700 47.465 22.870 48.095 ;
        RECT 23.500 48.225 23.830 48.705 ;
        RECT 24.000 48.415 24.225 48.875 ;
        RECT 24.395 48.225 24.725 48.705 ;
        RECT 23.500 48.055 24.725 48.225 ;
        RECT 24.915 48.075 25.165 48.875 ;
        RECT 25.335 48.075 25.675 48.705 ;
        RECT 25.445 48.025 25.675 48.075 ;
        RECT 23.040 47.685 23.370 47.885 ;
        RECT 23.540 47.685 23.870 47.885 ;
        RECT 24.040 47.685 24.460 47.885 ;
        RECT 24.635 47.715 25.330 47.885 ;
        RECT 24.635 47.465 24.805 47.715 ;
        RECT 25.500 47.465 25.675 48.025 ;
        RECT 15.265 46.325 20.610 46.760 ;
        RECT 20.785 46.325 21.995 47.415 ;
        RECT 22.370 47.295 24.805 47.465 ;
        RECT 22.370 46.495 22.700 47.295 ;
        RECT 22.870 46.325 23.200 47.125 ;
        RECT 23.500 46.495 23.830 47.295 ;
        RECT 24.475 46.325 24.725 47.125 ;
        RECT 24.995 46.325 25.165 47.465 ;
        RECT 25.335 46.495 25.675 47.465 ;
        RECT 25.845 48.075 26.185 48.705 ;
        RECT 26.355 48.075 26.605 48.875 ;
        RECT 26.795 48.225 27.125 48.705 ;
        RECT 27.295 48.415 27.520 48.875 ;
        RECT 27.690 48.225 28.020 48.705 ;
        RECT 25.845 47.465 26.020 48.075 ;
        RECT 26.795 48.055 28.020 48.225 ;
        RECT 28.650 48.095 29.150 48.705 ;
        RECT 29.525 48.105 31.195 48.875 ;
        RECT 31.365 48.150 31.655 48.875 ;
        RECT 31.825 48.330 37.170 48.875 ;
        RECT 37.345 48.330 42.690 48.875 ;
        RECT 42.865 48.330 48.210 48.875 ;
        RECT 26.190 47.715 26.885 47.885 ;
        RECT 26.715 47.465 26.885 47.715 ;
        RECT 27.060 47.685 27.480 47.885 ;
        RECT 27.650 47.685 27.980 47.885 ;
        RECT 28.150 47.685 28.480 47.885 ;
        RECT 28.650 47.465 28.820 48.095 ;
        RECT 29.005 47.635 29.355 47.885 ;
        RECT 29.525 47.585 30.275 48.105 ;
        RECT 25.845 46.495 26.185 47.465 ;
        RECT 26.355 46.325 26.525 47.465 ;
        RECT 26.715 47.295 29.150 47.465 ;
        RECT 30.445 47.415 31.195 47.935 ;
        RECT 33.410 47.500 33.750 48.330 ;
        RECT 26.795 46.325 27.045 47.125 ;
        RECT 27.690 46.495 28.020 47.295 ;
        RECT 28.320 46.325 28.650 47.125 ;
        RECT 28.820 46.495 29.150 47.295 ;
        RECT 29.525 46.325 31.195 47.415 ;
        RECT 31.365 46.325 31.655 47.490 ;
        RECT 35.230 46.760 35.580 48.010 ;
        RECT 38.930 47.500 39.270 48.330 ;
        RECT 40.750 46.760 41.100 48.010 ;
        RECT 44.450 47.500 44.790 48.330 ;
        RECT 49.050 48.095 49.550 48.705 ;
        RECT 46.270 46.760 46.620 48.010 ;
        RECT 48.845 47.635 49.195 47.885 ;
        RECT 49.380 47.465 49.550 48.095 ;
        RECT 50.180 48.225 50.510 48.705 ;
        RECT 50.680 48.415 50.905 48.875 ;
        RECT 51.075 48.225 51.405 48.705 ;
        RECT 50.180 48.055 51.405 48.225 ;
        RECT 51.595 48.075 51.845 48.875 ;
        RECT 52.015 48.075 52.355 48.705 ;
        RECT 52.125 48.025 52.355 48.075 ;
        RECT 49.720 47.685 50.050 47.885 ;
        RECT 50.220 47.685 50.550 47.885 ;
        RECT 50.720 47.685 51.140 47.885 ;
        RECT 51.315 47.715 52.010 47.885 ;
        RECT 51.315 47.465 51.485 47.715 ;
        RECT 52.180 47.465 52.355 48.025 ;
        RECT 52.525 48.105 56.035 48.875 ;
        RECT 57.125 48.150 57.415 48.875 ;
        RECT 57.585 48.105 60.175 48.875 ;
        RECT 60.435 48.325 60.605 48.705 ;
        RECT 60.820 48.495 61.150 48.875 ;
        RECT 60.435 48.155 61.150 48.325 ;
        RECT 52.525 47.585 54.175 48.105 ;
        RECT 49.050 47.295 51.485 47.465 ;
        RECT 31.825 46.325 37.170 46.760 ;
        RECT 37.345 46.325 42.690 46.760 ;
        RECT 42.865 46.325 48.210 46.760 ;
        RECT 49.050 46.495 49.380 47.295 ;
        RECT 49.550 46.325 49.880 47.125 ;
        RECT 50.180 46.495 50.510 47.295 ;
        RECT 51.155 46.325 51.405 47.125 ;
        RECT 51.675 46.325 51.845 47.465 ;
        RECT 52.015 46.495 52.355 47.465 ;
        RECT 54.345 47.415 56.035 47.935 ;
        RECT 57.585 47.585 58.795 48.105 ;
        RECT 52.525 46.325 56.035 47.415 ;
        RECT 57.125 46.325 57.415 47.490 ;
        RECT 58.965 47.415 60.175 47.935 ;
        RECT 60.345 47.605 60.700 47.975 ;
        RECT 60.980 47.965 61.150 48.155 ;
        RECT 61.320 48.130 61.575 48.705 ;
        RECT 60.980 47.635 61.235 47.965 ;
        RECT 60.980 47.425 61.150 47.635 ;
        RECT 57.585 46.325 60.175 47.415 ;
        RECT 60.435 47.255 61.150 47.425 ;
        RECT 61.405 47.400 61.575 48.130 ;
        RECT 61.750 48.035 62.010 48.875 ;
        RECT 62.335 48.075 62.665 48.875 ;
        RECT 62.835 48.225 63.005 48.705 ;
        RECT 63.175 48.395 63.505 48.875 ;
        RECT 63.675 48.225 63.845 48.705 ;
        RECT 64.095 48.395 64.335 48.875 ;
        RECT 64.515 48.225 64.685 48.705 ;
        RECT 62.835 48.055 63.845 48.225 ;
        RECT 64.050 48.055 64.685 48.225 ;
        RECT 64.945 48.105 66.615 48.875 ;
        RECT 66.790 48.325 67.045 48.615 ;
        RECT 67.215 48.495 67.545 48.875 ;
        RECT 66.790 48.155 67.540 48.325 ;
        RECT 62.835 47.515 63.330 48.055 ;
        RECT 64.050 47.885 64.220 48.055 ;
        RECT 63.720 47.715 64.220 47.885 ;
        RECT 60.435 46.495 60.605 47.255 ;
        RECT 60.820 46.325 61.150 47.085 ;
        RECT 61.320 46.495 61.575 47.400 ;
        RECT 61.750 46.325 62.010 47.475 ;
        RECT 62.335 46.325 62.665 47.475 ;
        RECT 62.835 47.345 63.845 47.515 ;
        RECT 62.835 46.495 63.005 47.345 ;
        RECT 63.175 46.325 63.505 47.125 ;
        RECT 63.675 46.495 63.845 47.345 ;
        RECT 64.050 47.475 64.220 47.715 ;
        RECT 64.390 47.645 64.770 47.885 ;
        RECT 64.945 47.585 65.695 48.105 ;
        RECT 64.050 47.305 64.765 47.475 ;
        RECT 65.865 47.415 66.615 47.935 ;
        RECT 64.025 46.325 64.265 47.125 ;
        RECT 64.435 46.495 64.765 47.305 ;
        RECT 64.945 46.325 66.615 47.415 ;
        RECT 66.790 47.335 67.140 47.985 ;
        RECT 67.310 47.165 67.540 48.155 ;
        RECT 66.790 46.995 67.540 47.165 ;
        RECT 66.790 46.495 67.045 46.995 ;
        RECT 67.215 46.325 67.545 46.825 ;
        RECT 67.715 46.495 67.885 48.615 ;
        RECT 68.245 48.515 68.575 48.875 ;
        RECT 68.745 48.485 69.240 48.655 ;
        RECT 69.445 48.485 70.300 48.655 ;
        RECT 68.115 47.295 68.575 48.345 ;
        RECT 68.055 46.510 68.380 47.295 ;
        RECT 68.745 47.125 68.915 48.485 ;
        RECT 69.085 47.575 69.435 48.195 ;
        RECT 69.605 47.975 69.960 48.195 ;
        RECT 69.605 47.385 69.775 47.975 ;
        RECT 70.130 47.775 70.300 48.485 ;
        RECT 71.175 48.415 71.505 48.875 ;
        RECT 71.715 48.515 72.065 48.685 ;
        RECT 70.505 47.945 71.295 48.195 ;
        RECT 71.715 48.125 71.975 48.515 ;
        RECT 72.285 48.425 73.235 48.705 ;
        RECT 73.405 48.435 73.595 48.875 ;
        RECT 73.765 48.495 74.835 48.665 ;
        RECT 71.465 47.775 71.635 47.955 ;
        RECT 68.745 46.955 69.140 47.125 ;
        RECT 69.310 46.995 69.775 47.385 ;
        RECT 69.945 47.605 71.635 47.775 ;
        RECT 68.970 46.825 69.140 46.955 ;
        RECT 69.945 46.825 70.115 47.605 ;
        RECT 71.805 47.435 71.975 48.125 ;
        RECT 70.475 47.265 71.975 47.435 ;
        RECT 72.165 47.465 72.375 48.255 ;
        RECT 72.545 47.635 72.895 48.255 ;
        RECT 73.065 47.645 73.235 48.425 ;
        RECT 73.765 48.265 73.935 48.495 ;
        RECT 73.405 48.095 73.935 48.265 ;
        RECT 73.405 47.815 73.625 48.095 ;
        RECT 74.105 47.925 74.345 48.325 ;
        RECT 73.065 47.475 73.470 47.645 ;
        RECT 73.805 47.555 74.345 47.925 ;
        RECT 74.515 48.140 74.835 48.495 ;
        RECT 75.080 48.415 75.385 48.875 ;
        RECT 75.555 48.165 75.810 48.695 ;
        RECT 74.515 47.965 74.840 48.140 ;
        RECT 74.515 47.665 75.430 47.965 ;
        RECT 74.690 47.635 75.430 47.665 ;
        RECT 72.165 47.305 72.840 47.465 ;
        RECT 73.300 47.385 73.470 47.475 ;
        RECT 72.165 47.295 73.130 47.305 ;
        RECT 71.805 47.125 71.975 47.265 ;
        RECT 68.550 46.325 68.800 46.785 ;
        RECT 68.970 46.495 69.220 46.825 ;
        RECT 69.435 46.495 70.115 46.825 ;
        RECT 70.285 46.925 71.360 47.095 ;
        RECT 71.805 46.955 72.365 47.125 ;
        RECT 72.670 47.005 73.130 47.295 ;
        RECT 73.300 47.215 74.520 47.385 ;
        RECT 70.285 46.585 70.455 46.925 ;
        RECT 70.690 46.325 71.020 46.755 ;
        RECT 71.190 46.585 71.360 46.925 ;
        RECT 71.655 46.325 72.025 46.785 ;
        RECT 72.195 46.495 72.365 46.955 ;
        RECT 73.300 46.835 73.470 47.215 ;
        RECT 74.690 47.045 74.860 47.635 ;
        RECT 75.600 47.515 75.810 48.165 ;
        RECT 72.600 46.495 73.470 46.835 ;
        RECT 74.060 46.875 74.860 47.045 ;
        RECT 73.640 46.325 73.890 46.785 ;
        RECT 74.060 46.585 74.230 46.875 ;
        RECT 74.410 46.325 74.740 46.705 ;
        RECT 75.080 46.325 75.385 47.465 ;
        RECT 75.555 46.635 75.810 47.515 ;
        RECT 75.990 48.135 76.245 48.705 ;
        RECT 76.415 48.475 76.745 48.875 ;
        RECT 77.170 48.340 77.700 48.705 ;
        RECT 77.170 48.305 77.345 48.340 ;
        RECT 76.415 48.135 77.345 48.305 ;
        RECT 75.990 47.465 76.160 48.135 ;
        RECT 76.415 47.965 76.585 48.135 ;
        RECT 76.330 47.635 76.585 47.965 ;
        RECT 76.810 47.635 77.005 47.965 ;
        RECT 75.990 46.495 76.325 47.465 ;
        RECT 76.495 46.325 76.665 47.465 ;
        RECT 76.835 46.665 77.005 47.635 ;
        RECT 77.175 47.005 77.345 48.135 ;
        RECT 77.515 47.345 77.685 48.145 ;
        RECT 77.890 47.855 78.165 48.705 ;
        RECT 77.885 47.685 78.165 47.855 ;
        RECT 77.890 47.545 78.165 47.685 ;
        RECT 78.335 47.345 78.525 48.705 ;
        RECT 78.705 48.340 79.215 48.875 ;
        RECT 79.435 48.065 79.680 48.670 ;
        RECT 80.125 48.105 82.715 48.875 ;
        RECT 82.885 48.150 83.175 48.875 ;
        RECT 83.345 48.135 83.730 48.705 ;
        RECT 83.900 48.415 84.225 48.875 ;
        RECT 84.745 48.245 85.025 48.705 ;
        RECT 78.725 47.895 79.955 48.065 ;
        RECT 77.515 47.175 78.525 47.345 ;
        RECT 78.695 47.330 79.445 47.520 ;
        RECT 77.175 46.835 78.300 47.005 ;
        RECT 78.695 46.665 78.865 47.330 ;
        RECT 79.615 47.085 79.955 47.895 ;
        RECT 80.125 47.585 81.335 48.105 ;
        RECT 81.505 47.415 82.715 47.935 ;
        RECT 76.835 46.495 78.865 46.665 ;
        RECT 79.035 46.325 79.205 47.085 ;
        RECT 79.440 46.675 79.955 47.085 ;
        RECT 80.125 46.325 82.715 47.415 ;
        RECT 82.885 46.325 83.175 47.490 ;
        RECT 83.345 47.465 83.625 48.135 ;
        RECT 83.900 48.075 85.025 48.245 ;
        RECT 83.900 47.965 84.350 48.075 ;
        RECT 83.795 47.635 84.350 47.965 ;
        RECT 85.215 47.905 85.615 48.705 ;
        RECT 86.015 48.415 86.285 48.875 ;
        RECT 86.455 48.245 86.740 48.705 ;
        RECT 83.345 46.495 83.730 47.465 ;
        RECT 83.900 47.175 84.350 47.635 ;
        RECT 84.520 47.345 85.615 47.905 ;
        RECT 83.900 46.955 85.025 47.175 ;
        RECT 83.900 46.325 84.225 46.785 ;
        RECT 84.745 46.495 85.025 46.955 ;
        RECT 85.215 46.495 85.615 47.345 ;
        RECT 85.785 48.075 86.740 48.245 ;
        RECT 87.025 48.075 87.365 48.705 ;
        RECT 87.535 48.075 87.785 48.875 ;
        RECT 87.975 48.225 88.305 48.705 ;
        RECT 88.475 48.415 88.700 48.875 ;
        RECT 88.870 48.225 89.200 48.705 ;
        RECT 85.785 47.175 85.995 48.075 ;
        RECT 87.025 48.025 87.255 48.075 ;
        RECT 87.975 48.055 89.200 48.225 ;
        RECT 89.830 48.095 90.330 48.705 ;
        RECT 90.910 48.095 91.410 48.705 ;
        RECT 86.165 47.345 86.855 47.905 ;
        RECT 87.025 47.465 87.200 48.025 ;
        RECT 87.370 47.715 88.065 47.885 ;
        RECT 87.895 47.465 88.065 47.715 ;
        RECT 88.240 47.685 88.660 47.885 ;
        RECT 88.830 47.685 89.160 47.885 ;
        RECT 89.330 47.685 89.660 47.885 ;
        RECT 89.830 47.465 90.000 48.095 ;
        RECT 90.185 47.635 90.535 47.885 ;
        RECT 90.705 47.635 91.055 47.885 ;
        RECT 91.240 47.465 91.410 48.095 ;
        RECT 92.040 48.225 92.370 48.705 ;
        RECT 92.540 48.415 92.765 48.875 ;
        RECT 92.935 48.225 93.265 48.705 ;
        RECT 92.040 48.055 93.265 48.225 ;
        RECT 93.455 48.075 93.705 48.875 ;
        RECT 93.875 48.075 94.215 48.705 ;
        RECT 91.580 47.685 91.910 47.885 ;
        RECT 92.080 47.685 92.410 47.885 ;
        RECT 92.580 47.685 93.000 47.885 ;
        RECT 93.175 47.715 93.870 47.885 ;
        RECT 93.175 47.465 93.345 47.715 ;
        RECT 94.040 47.465 94.215 48.075 ;
        RECT 85.785 46.955 86.740 47.175 ;
        RECT 86.015 46.325 86.285 46.785 ;
        RECT 86.455 46.495 86.740 46.955 ;
        RECT 87.025 46.495 87.365 47.465 ;
        RECT 87.535 46.325 87.705 47.465 ;
        RECT 87.895 47.295 90.330 47.465 ;
        RECT 87.975 46.325 88.225 47.125 ;
        RECT 88.870 46.495 89.200 47.295 ;
        RECT 89.500 46.325 89.830 47.125 ;
        RECT 90.000 46.495 90.330 47.295 ;
        RECT 90.910 47.295 93.345 47.465 ;
        RECT 90.910 46.495 91.240 47.295 ;
        RECT 91.410 46.325 91.740 47.125 ;
        RECT 92.040 46.495 92.370 47.295 ;
        RECT 93.015 46.325 93.265 47.125 ;
        RECT 93.535 46.325 93.705 47.465 ;
        RECT 93.875 46.495 94.215 47.465 ;
        RECT 94.385 48.075 94.725 48.705 ;
        RECT 94.895 48.075 95.145 48.875 ;
        RECT 95.335 48.225 95.665 48.705 ;
        RECT 95.835 48.415 96.060 48.875 ;
        RECT 96.230 48.225 96.560 48.705 ;
        RECT 94.385 48.025 94.615 48.075 ;
        RECT 95.335 48.055 96.560 48.225 ;
        RECT 97.190 48.095 97.690 48.705 ;
        RECT 94.385 47.465 94.560 48.025 ;
        RECT 94.730 47.715 95.425 47.885 ;
        RECT 95.255 47.465 95.425 47.715 ;
        RECT 95.600 47.685 96.020 47.885 ;
        RECT 96.190 47.685 96.520 47.885 ;
        RECT 96.690 47.685 97.020 47.885 ;
        RECT 97.190 47.465 97.360 48.095 ;
        RECT 98.800 48.065 99.045 48.670 ;
        RECT 99.265 48.340 99.775 48.875 ;
        RECT 98.525 47.895 99.755 48.065 ;
        RECT 97.545 47.635 97.895 47.885 ;
        RECT 94.385 46.495 94.725 47.465 ;
        RECT 94.895 46.325 95.065 47.465 ;
        RECT 95.255 47.295 97.690 47.465 ;
        RECT 95.335 46.325 95.585 47.125 ;
        RECT 96.230 46.495 96.560 47.295 ;
        RECT 96.860 46.325 97.190 47.125 ;
        RECT 97.360 46.495 97.690 47.295 ;
        RECT 98.525 47.085 98.865 47.895 ;
        RECT 99.035 47.330 99.785 47.520 ;
        RECT 98.525 46.675 99.040 47.085 ;
        RECT 99.275 46.325 99.445 47.085 ;
        RECT 99.615 46.665 99.785 47.330 ;
        RECT 99.955 47.345 100.145 48.705 ;
        RECT 100.315 47.855 100.590 48.705 ;
        RECT 100.780 48.340 101.310 48.705 ;
        RECT 101.735 48.475 102.065 48.875 ;
        RECT 101.135 48.305 101.310 48.340 ;
        RECT 100.315 47.685 100.595 47.855 ;
        RECT 100.315 47.545 100.590 47.685 ;
        RECT 100.795 47.345 100.965 48.145 ;
        RECT 99.955 47.175 100.965 47.345 ;
        RECT 101.135 48.135 102.065 48.305 ;
        RECT 102.235 48.135 102.490 48.705 ;
        RECT 101.135 47.005 101.305 48.135 ;
        RECT 101.895 47.965 102.065 48.135 ;
        RECT 100.180 46.835 101.305 47.005 ;
        RECT 101.475 47.635 101.670 47.965 ;
        RECT 101.895 47.635 102.150 47.965 ;
        RECT 101.475 46.665 101.645 47.635 ;
        RECT 102.320 47.465 102.490 48.135 ;
        RECT 99.615 46.495 101.645 46.665 ;
        RECT 101.815 46.325 101.985 47.465 ;
        RECT 102.155 46.495 102.490 47.465 ;
        RECT 102.665 48.135 103.050 48.705 ;
        RECT 103.220 48.415 103.545 48.875 ;
        RECT 104.065 48.245 104.345 48.705 ;
        RECT 102.665 47.465 102.945 48.135 ;
        RECT 103.220 48.075 104.345 48.245 ;
        RECT 103.220 47.965 103.670 48.075 ;
        RECT 103.115 47.635 103.670 47.965 ;
        RECT 104.535 47.905 104.935 48.705 ;
        RECT 105.335 48.415 105.605 48.875 ;
        RECT 105.775 48.245 106.060 48.705 ;
        RECT 102.665 46.495 103.050 47.465 ;
        RECT 103.220 47.175 103.670 47.635 ;
        RECT 103.840 47.345 104.935 47.905 ;
        RECT 103.220 46.955 104.345 47.175 ;
        RECT 103.220 46.325 103.545 46.785 ;
        RECT 104.065 46.495 104.345 46.955 ;
        RECT 104.535 46.495 104.935 47.345 ;
        RECT 105.105 48.075 106.060 48.245 ;
        RECT 106.435 48.325 106.605 48.705 ;
        RECT 106.785 48.495 107.115 48.875 ;
        RECT 106.435 48.155 107.100 48.325 ;
        RECT 107.295 48.200 107.555 48.705 ;
        RECT 105.105 47.175 105.315 48.075 ;
        RECT 105.485 47.345 106.175 47.905 ;
        RECT 106.365 47.605 106.695 47.975 ;
        RECT 106.930 47.900 107.100 48.155 ;
        RECT 106.930 47.570 107.215 47.900 ;
        RECT 106.930 47.425 107.100 47.570 ;
        RECT 106.435 47.255 107.100 47.425 ;
        RECT 107.385 47.400 107.555 48.200 ;
        RECT 108.645 48.150 108.935 48.875 ;
        RECT 109.105 48.330 114.450 48.875 ;
        RECT 110.690 47.500 111.030 48.330 ;
        RECT 114.625 48.105 117.215 48.875 ;
        RECT 117.385 48.125 118.595 48.875 ;
        RECT 105.105 46.955 106.060 47.175 ;
        RECT 105.335 46.325 105.605 46.785 ;
        RECT 105.775 46.495 106.060 46.955 ;
        RECT 106.435 46.495 106.605 47.255 ;
        RECT 106.785 46.325 107.115 47.085 ;
        RECT 107.285 46.495 107.555 47.400 ;
        RECT 108.645 46.325 108.935 47.490 ;
        RECT 112.510 46.760 112.860 48.010 ;
        RECT 114.625 47.585 115.835 48.105 ;
        RECT 116.005 47.415 117.215 47.935 ;
        RECT 109.105 46.325 114.450 46.760 ;
        RECT 114.625 46.325 117.215 47.415 ;
        RECT 117.385 47.415 117.905 47.955 ;
        RECT 118.075 47.585 118.595 48.125 ;
        RECT 117.385 46.325 118.595 47.415 ;
        RECT 5.520 46.155 118.680 46.325 ;
        RECT 5.605 45.065 6.815 46.155 ;
        RECT 6.985 45.720 12.330 46.155 ;
        RECT 5.605 44.355 6.125 44.895 ;
        RECT 6.295 44.525 6.815 45.065 ;
        RECT 5.605 43.605 6.815 44.355 ;
        RECT 8.570 44.150 8.910 44.980 ;
        RECT 10.390 44.470 10.740 45.720 ;
        RECT 12.505 45.065 15.095 46.155 ;
        RECT 12.505 44.375 13.715 44.895 ;
        RECT 13.885 44.545 15.095 45.065 ;
        RECT 15.265 45.080 15.535 45.985 ;
        RECT 15.705 45.395 16.035 46.155 ;
        RECT 16.215 45.225 16.385 45.985 ;
        RECT 6.985 43.605 12.330 44.150 ;
        RECT 12.505 43.605 15.095 44.375 ;
        RECT 15.265 44.280 15.435 45.080 ;
        RECT 15.720 45.055 16.385 45.225 ;
        RECT 16.645 45.065 18.315 46.155 ;
        RECT 15.720 44.910 15.890 45.055 ;
        RECT 15.605 44.580 15.890 44.910 ;
        RECT 15.720 44.325 15.890 44.580 ;
        RECT 16.125 44.505 16.455 44.875 ;
        RECT 16.645 44.375 17.395 44.895 ;
        RECT 17.565 44.545 18.315 45.065 ;
        RECT 18.485 44.990 18.775 46.155 ;
        RECT 18.950 45.015 19.285 45.985 ;
        RECT 19.455 45.015 19.625 46.155 ;
        RECT 19.795 45.815 21.825 45.985 ;
        RECT 15.265 43.775 15.525 44.280 ;
        RECT 15.720 44.155 16.385 44.325 ;
        RECT 15.705 43.605 16.035 43.985 ;
        RECT 16.215 43.775 16.385 44.155 ;
        RECT 16.645 43.605 18.315 44.375 ;
        RECT 18.950 44.345 19.120 45.015 ;
        RECT 19.795 44.845 19.965 45.815 ;
        RECT 19.290 44.515 19.545 44.845 ;
        RECT 19.770 44.515 19.965 44.845 ;
        RECT 20.135 45.475 21.260 45.645 ;
        RECT 19.375 44.345 19.545 44.515 ;
        RECT 20.135 44.345 20.305 45.475 ;
        RECT 18.485 43.605 18.775 44.330 ;
        RECT 18.950 43.775 19.205 44.345 ;
        RECT 19.375 44.175 20.305 44.345 ;
        RECT 20.475 45.135 21.485 45.305 ;
        RECT 20.475 44.335 20.645 45.135 ;
        RECT 20.130 44.140 20.305 44.175 ;
        RECT 19.375 43.605 19.705 44.005 ;
        RECT 20.130 43.775 20.660 44.140 ;
        RECT 20.850 44.115 21.125 44.935 ;
        RECT 20.845 43.945 21.125 44.115 ;
        RECT 20.850 43.775 21.125 43.945 ;
        RECT 21.295 43.775 21.485 45.135 ;
        RECT 21.655 45.150 21.825 45.815 ;
        RECT 21.995 45.395 22.165 46.155 ;
        RECT 22.400 45.395 22.915 45.805 ;
        RECT 21.655 44.960 22.405 45.150 ;
        RECT 22.575 44.585 22.915 45.395 ;
        RECT 23.085 45.065 24.755 46.155 ;
        RECT 21.685 44.415 22.915 44.585 ;
        RECT 21.665 43.605 22.175 44.140 ;
        RECT 22.395 43.810 22.640 44.415 ;
        RECT 23.085 44.375 23.835 44.895 ;
        RECT 24.005 44.545 24.755 45.065 ;
        RECT 25.130 45.185 25.460 45.985 ;
        RECT 25.630 45.355 25.960 46.155 ;
        RECT 26.260 45.185 26.590 45.985 ;
        RECT 27.235 45.355 27.485 46.155 ;
        RECT 25.130 45.015 27.565 45.185 ;
        RECT 27.755 45.015 27.925 46.155 ;
        RECT 28.095 45.015 28.435 45.985 ;
        RECT 28.605 45.065 29.815 46.155 ;
        RECT 24.925 44.595 25.275 44.845 ;
        RECT 25.460 44.385 25.630 45.015 ;
        RECT 25.800 44.595 26.130 44.795 ;
        RECT 26.300 44.595 26.630 44.795 ;
        RECT 26.800 44.595 27.220 44.795 ;
        RECT 27.395 44.765 27.565 45.015 ;
        RECT 27.395 44.595 28.090 44.765 ;
        RECT 23.085 43.605 24.755 44.375 ;
        RECT 25.130 43.775 25.630 44.385 ;
        RECT 26.260 44.255 27.485 44.425 ;
        RECT 28.260 44.405 28.435 45.015 ;
        RECT 26.260 43.775 26.590 44.255 ;
        RECT 26.760 43.605 26.985 44.065 ;
        RECT 27.155 43.775 27.485 44.255 ;
        RECT 27.675 43.605 27.925 44.405 ;
        RECT 28.095 43.775 28.435 44.405 ;
        RECT 28.605 44.355 29.125 44.895 ;
        RECT 29.295 44.525 29.815 45.065 ;
        RECT 30.075 45.225 30.245 45.985 ;
        RECT 30.425 45.395 30.755 46.155 ;
        RECT 30.075 45.055 30.740 45.225 ;
        RECT 30.925 45.080 31.195 45.985 ;
        RECT 30.570 44.910 30.740 45.055 ;
        RECT 30.005 44.505 30.335 44.875 ;
        RECT 30.570 44.580 30.855 44.910 ;
        RECT 28.605 43.605 29.815 44.355 ;
        RECT 30.570 44.325 30.740 44.580 ;
        RECT 30.075 44.155 30.740 44.325 ;
        RECT 31.025 44.280 31.195 45.080 ;
        RECT 30.075 43.775 30.245 44.155 ;
        RECT 30.425 43.605 30.755 43.985 ;
        RECT 30.935 43.775 31.195 44.280 ;
        RECT 31.365 45.015 31.705 45.985 ;
        RECT 31.875 45.015 32.045 46.155 ;
        RECT 32.315 45.355 32.565 46.155 ;
        RECT 33.210 45.185 33.540 45.985 ;
        RECT 33.840 45.355 34.170 46.155 ;
        RECT 34.340 45.185 34.670 45.985 ;
        RECT 35.045 45.720 40.390 46.155 ;
        RECT 32.235 45.015 34.670 45.185 ;
        RECT 31.365 44.405 31.540 45.015 ;
        RECT 32.235 44.765 32.405 45.015 ;
        RECT 31.710 44.595 32.405 44.765 ;
        RECT 32.580 44.595 33.000 44.795 ;
        RECT 33.170 44.595 33.500 44.795 ;
        RECT 33.670 44.595 34.000 44.795 ;
        RECT 31.365 43.775 31.705 44.405 ;
        RECT 31.875 43.605 32.125 44.405 ;
        RECT 32.315 44.255 33.540 44.425 ;
        RECT 32.315 43.775 32.645 44.255 ;
        RECT 32.815 43.605 33.040 44.065 ;
        RECT 33.210 43.775 33.540 44.255 ;
        RECT 34.170 44.385 34.340 45.015 ;
        RECT 34.525 44.595 34.875 44.845 ;
        RECT 34.170 43.775 34.670 44.385 ;
        RECT 36.630 44.150 36.970 44.980 ;
        RECT 38.450 44.470 38.800 45.720 ;
        RECT 40.565 45.065 44.075 46.155 ;
        RECT 40.565 44.375 42.215 44.895 ;
        RECT 42.385 44.545 44.075 45.065 ;
        RECT 44.245 44.990 44.535 46.155 ;
        RECT 44.705 45.015 45.090 45.985 ;
        RECT 45.260 45.695 45.585 46.155 ;
        RECT 46.105 45.525 46.385 45.985 ;
        RECT 45.260 45.305 46.385 45.525 ;
        RECT 35.045 43.605 40.390 44.150 ;
        RECT 40.565 43.605 44.075 44.375 ;
        RECT 44.705 44.345 44.985 45.015 ;
        RECT 45.260 44.845 45.710 45.305 ;
        RECT 46.575 45.135 46.975 45.985 ;
        RECT 47.375 45.695 47.645 46.155 ;
        RECT 47.815 45.525 48.100 45.985 ;
        RECT 45.155 44.515 45.710 44.845 ;
        RECT 45.880 44.575 46.975 45.135 ;
        RECT 45.260 44.405 45.710 44.515 ;
        RECT 44.245 43.605 44.535 44.330 ;
        RECT 44.705 43.775 45.090 44.345 ;
        RECT 45.260 44.235 46.385 44.405 ;
        RECT 45.260 43.605 45.585 44.065 ;
        RECT 46.105 43.775 46.385 44.235 ;
        RECT 46.575 43.775 46.975 44.575 ;
        RECT 47.145 45.305 48.100 45.525 ;
        RECT 47.145 44.405 47.355 45.305 ;
        RECT 47.525 44.575 48.215 45.135 ;
        RECT 48.385 45.065 49.595 46.155 ;
        RECT 47.145 44.235 48.100 44.405 ;
        RECT 47.375 43.605 47.645 44.065 ;
        RECT 47.815 43.775 48.100 44.235 ;
        RECT 48.385 44.355 48.905 44.895 ;
        RECT 49.075 44.525 49.595 45.065 ;
        RECT 49.970 45.185 50.300 45.985 ;
        RECT 50.470 45.355 50.800 46.155 ;
        RECT 51.100 45.185 51.430 45.985 ;
        RECT 52.075 45.355 52.325 46.155 ;
        RECT 49.970 45.015 52.405 45.185 ;
        RECT 52.595 45.015 52.765 46.155 ;
        RECT 52.935 45.015 53.275 45.985 ;
        RECT 49.765 44.595 50.115 44.845 ;
        RECT 50.300 44.385 50.470 45.015 ;
        RECT 50.640 44.595 50.970 44.795 ;
        RECT 51.140 44.595 51.470 44.795 ;
        RECT 51.640 44.595 52.060 44.795 ;
        RECT 52.235 44.765 52.405 45.015 ;
        RECT 52.235 44.595 52.930 44.765 ;
        RECT 53.100 44.455 53.275 45.015 ;
        RECT 48.385 43.605 49.595 44.355 ;
        RECT 49.970 43.775 50.470 44.385 ;
        RECT 51.100 44.255 52.325 44.425 ;
        RECT 53.045 44.405 53.275 44.455 ;
        RECT 51.100 43.775 51.430 44.255 ;
        RECT 51.600 43.605 51.825 44.065 ;
        RECT 51.995 43.775 52.325 44.255 ;
        RECT 52.515 43.605 52.765 44.405 ;
        RECT 52.935 43.775 53.275 44.405 ;
        RECT 53.445 45.015 53.785 45.985 ;
        RECT 53.955 45.015 54.125 46.155 ;
        RECT 54.395 45.355 54.645 46.155 ;
        RECT 55.290 45.185 55.620 45.985 ;
        RECT 55.920 45.355 56.250 46.155 ;
        RECT 56.420 45.185 56.750 45.985 ;
        RECT 54.315 45.015 56.750 45.185 ;
        RECT 57.595 45.095 57.925 46.155 ;
        RECT 53.445 44.965 53.675 45.015 ;
        RECT 53.445 44.405 53.620 44.965 ;
        RECT 54.315 44.765 54.485 45.015 ;
        RECT 53.790 44.595 54.485 44.765 ;
        RECT 54.660 44.595 55.080 44.795 ;
        RECT 55.250 44.595 55.580 44.795 ;
        RECT 55.750 44.595 56.080 44.795 ;
        RECT 53.445 43.775 53.785 44.405 ;
        RECT 53.955 43.605 54.205 44.405 ;
        RECT 54.395 44.255 55.620 44.425 ;
        RECT 54.395 43.775 54.725 44.255 ;
        RECT 54.895 43.605 55.120 44.065 ;
        RECT 55.290 43.775 55.620 44.255 ;
        RECT 56.250 44.385 56.420 45.015 ;
        RECT 58.105 44.845 58.275 45.770 ;
        RECT 58.445 45.565 58.775 45.965 ;
        RECT 58.945 45.795 59.275 46.155 ;
        RECT 59.475 45.565 60.175 45.985 ;
        RECT 58.445 45.335 60.175 45.565 ;
        RECT 58.445 45.115 58.775 45.335 ;
        RECT 58.970 44.845 59.295 45.135 ;
        RECT 56.605 44.595 56.955 44.845 ;
        RECT 57.585 44.515 57.895 44.845 ;
        RECT 58.105 44.515 58.480 44.845 ;
        RECT 58.800 44.515 59.295 44.845 ;
        RECT 59.470 44.595 59.800 45.135 ;
        RECT 56.250 43.775 56.750 44.385 ;
        RECT 59.970 44.365 60.175 45.335 ;
        RECT 60.350 45.005 60.610 46.155 ;
        RECT 60.785 45.080 61.040 45.985 ;
        RECT 61.210 45.395 61.540 46.155 ;
        RECT 61.755 45.225 61.925 45.985 ;
        RECT 57.595 44.135 58.955 44.345 ;
        RECT 57.595 43.775 57.925 44.135 ;
        RECT 58.095 43.605 58.425 43.965 ;
        RECT 58.625 43.775 58.955 44.135 ;
        RECT 59.465 43.775 60.175 44.365 ;
        RECT 60.350 43.605 60.610 44.445 ;
        RECT 60.785 44.350 60.955 45.080 ;
        RECT 61.210 45.055 61.925 45.225 ;
        RECT 61.210 44.845 61.380 45.055 ;
        RECT 62.190 45.005 62.450 46.155 ;
        RECT 62.625 45.080 62.880 45.985 ;
        RECT 63.050 45.395 63.380 46.155 ;
        RECT 63.595 45.225 63.765 45.985 ;
        RECT 61.125 44.515 61.380 44.845 ;
        RECT 60.785 43.775 61.040 44.350 ;
        RECT 61.210 44.325 61.380 44.515 ;
        RECT 61.660 44.505 62.015 44.875 ;
        RECT 61.210 44.155 61.925 44.325 ;
        RECT 61.210 43.605 61.540 43.985 ;
        RECT 61.755 43.775 61.925 44.155 ;
        RECT 62.190 43.605 62.450 44.445 ;
        RECT 62.625 44.350 62.795 45.080 ;
        RECT 63.050 45.055 63.765 45.225 ;
        RECT 64.115 45.225 64.285 45.985 ;
        RECT 64.500 45.395 64.830 46.155 ;
        RECT 64.115 45.055 64.830 45.225 ;
        RECT 65.000 45.080 65.255 45.985 ;
        RECT 63.050 44.845 63.220 45.055 ;
        RECT 62.965 44.515 63.220 44.845 ;
        RECT 62.625 43.775 62.880 44.350 ;
        RECT 63.050 44.325 63.220 44.515 ;
        RECT 63.500 44.505 63.855 44.875 ;
        RECT 64.025 44.505 64.380 44.875 ;
        RECT 64.660 44.845 64.830 45.055 ;
        RECT 64.660 44.515 64.915 44.845 ;
        RECT 64.660 44.325 64.830 44.515 ;
        RECT 65.085 44.350 65.255 45.080 ;
        RECT 65.430 45.005 65.690 46.155 ;
        RECT 65.865 45.065 68.455 46.155 ;
        RECT 63.050 44.155 63.765 44.325 ;
        RECT 63.050 43.605 63.380 43.985 ;
        RECT 63.595 43.775 63.765 44.155 ;
        RECT 64.115 44.155 64.830 44.325 ;
        RECT 64.115 43.775 64.285 44.155 ;
        RECT 64.500 43.605 64.830 43.985 ;
        RECT 65.000 43.775 65.255 44.350 ;
        RECT 65.430 43.605 65.690 44.445 ;
        RECT 65.865 44.375 67.075 44.895 ;
        RECT 67.245 44.545 68.455 45.065 ;
        RECT 68.715 45.225 68.885 45.985 ;
        RECT 69.065 45.395 69.395 46.155 ;
        RECT 68.715 45.055 69.380 45.225 ;
        RECT 69.565 45.080 69.835 45.985 ;
        RECT 69.210 44.910 69.380 45.055 ;
        RECT 68.645 44.505 68.975 44.875 ;
        RECT 69.210 44.580 69.495 44.910 ;
        RECT 65.865 43.605 68.455 44.375 ;
        RECT 69.210 44.325 69.380 44.580 ;
        RECT 68.715 44.155 69.380 44.325 ;
        RECT 69.665 44.280 69.835 45.080 ;
        RECT 70.005 44.990 70.295 46.155 ;
        RECT 70.470 45.485 70.725 45.985 ;
        RECT 70.895 45.655 71.225 46.155 ;
        RECT 70.470 45.315 71.220 45.485 ;
        RECT 70.470 44.495 70.820 45.145 ;
        RECT 68.715 43.775 68.885 44.155 ;
        RECT 69.065 43.605 69.395 43.985 ;
        RECT 69.575 43.775 69.835 44.280 ;
        RECT 70.005 43.605 70.295 44.330 ;
        RECT 70.990 44.325 71.220 45.315 ;
        RECT 70.470 44.155 71.220 44.325 ;
        RECT 70.470 43.865 70.725 44.155 ;
        RECT 70.895 43.605 71.225 43.985 ;
        RECT 71.395 43.865 71.565 45.985 ;
        RECT 71.735 45.185 72.060 45.970 ;
        RECT 72.230 45.695 72.480 46.155 ;
        RECT 72.650 45.655 72.900 45.985 ;
        RECT 73.115 45.655 73.795 45.985 ;
        RECT 72.650 45.525 72.820 45.655 ;
        RECT 72.425 45.355 72.820 45.525 ;
        RECT 71.795 44.135 72.255 45.185 ;
        RECT 72.425 43.995 72.595 45.355 ;
        RECT 72.990 45.095 73.455 45.485 ;
        RECT 72.765 44.285 73.115 44.905 ;
        RECT 73.285 44.505 73.455 45.095 ;
        RECT 73.625 44.875 73.795 45.655 ;
        RECT 73.965 45.555 74.135 45.895 ;
        RECT 74.370 45.725 74.700 46.155 ;
        RECT 74.870 45.555 75.040 45.895 ;
        RECT 75.335 45.695 75.705 46.155 ;
        RECT 73.965 45.385 75.040 45.555 ;
        RECT 75.875 45.525 76.045 45.985 ;
        RECT 76.280 45.645 77.150 45.985 ;
        RECT 77.320 45.695 77.570 46.155 ;
        RECT 75.485 45.355 76.045 45.525 ;
        RECT 75.485 45.215 75.655 45.355 ;
        RECT 74.155 45.045 75.655 45.215 ;
        RECT 76.350 45.185 76.810 45.475 ;
        RECT 73.625 44.705 75.315 44.875 ;
        RECT 73.285 44.285 73.640 44.505 ;
        RECT 73.810 43.995 73.980 44.705 ;
        RECT 74.185 44.285 74.975 44.535 ;
        RECT 75.145 44.525 75.315 44.705 ;
        RECT 75.485 44.355 75.655 45.045 ;
        RECT 71.925 43.605 72.255 43.965 ;
        RECT 72.425 43.825 72.920 43.995 ;
        RECT 73.125 43.825 73.980 43.995 ;
        RECT 74.855 43.605 75.185 44.065 ;
        RECT 75.395 43.965 75.655 44.355 ;
        RECT 75.845 45.175 76.810 45.185 ;
        RECT 76.980 45.265 77.150 45.645 ;
        RECT 77.740 45.605 77.910 45.895 ;
        RECT 78.090 45.775 78.420 46.155 ;
        RECT 77.740 45.435 78.540 45.605 ;
        RECT 75.845 45.015 76.520 45.175 ;
        RECT 76.980 45.095 78.200 45.265 ;
        RECT 75.845 44.225 76.055 45.015 ;
        RECT 76.980 45.005 77.150 45.095 ;
        RECT 76.225 44.225 76.575 44.845 ;
        RECT 76.745 44.835 77.150 45.005 ;
        RECT 76.745 44.055 76.915 44.835 ;
        RECT 77.085 44.385 77.305 44.665 ;
        RECT 77.485 44.555 78.025 44.925 ;
        RECT 78.370 44.845 78.540 45.435 ;
        RECT 78.760 45.015 79.065 46.155 ;
        RECT 79.235 44.965 79.490 45.845 ;
        RECT 78.370 44.815 79.110 44.845 ;
        RECT 77.085 44.215 77.615 44.385 ;
        RECT 75.395 43.795 75.745 43.965 ;
        RECT 75.965 43.775 76.915 44.055 ;
        RECT 77.085 43.605 77.275 44.045 ;
        RECT 77.445 43.985 77.615 44.215 ;
        RECT 77.785 44.155 78.025 44.555 ;
        RECT 78.195 44.515 79.110 44.815 ;
        RECT 78.195 44.340 78.520 44.515 ;
        RECT 78.195 43.985 78.515 44.340 ;
        RECT 79.280 44.315 79.490 44.965 ;
        RECT 77.445 43.815 78.515 43.985 ;
        RECT 78.760 43.605 79.065 44.065 ;
        RECT 79.235 43.785 79.490 44.315 ;
        RECT 79.665 45.015 80.050 45.985 ;
        RECT 80.220 45.695 80.545 46.155 ;
        RECT 81.065 45.525 81.345 45.985 ;
        RECT 80.220 45.305 81.345 45.525 ;
        RECT 79.665 44.345 79.945 45.015 ;
        RECT 80.220 44.845 80.670 45.305 ;
        RECT 81.535 45.135 81.935 45.985 ;
        RECT 82.335 45.695 82.605 46.155 ;
        RECT 82.775 45.525 83.060 45.985 ;
        RECT 80.115 44.515 80.670 44.845 ;
        RECT 80.840 44.575 81.935 45.135 ;
        RECT 80.220 44.405 80.670 44.515 ;
        RECT 79.665 43.775 80.050 44.345 ;
        RECT 80.220 44.235 81.345 44.405 ;
        RECT 80.220 43.605 80.545 44.065 ;
        RECT 81.065 43.775 81.345 44.235 ;
        RECT 81.535 43.775 81.935 44.575 ;
        RECT 82.105 45.305 83.060 45.525 ;
        RECT 82.105 44.405 82.315 45.305 ;
        RECT 82.485 44.575 83.175 45.135 ;
        RECT 83.345 45.015 83.685 45.985 ;
        RECT 83.855 45.015 84.025 46.155 ;
        RECT 84.295 45.355 84.545 46.155 ;
        RECT 85.190 45.185 85.520 45.985 ;
        RECT 85.820 45.355 86.150 46.155 ;
        RECT 86.320 45.185 86.650 45.985 ;
        RECT 84.215 45.015 86.650 45.185 ;
        RECT 87.025 45.015 87.410 45.985 ;
        RECT 87.580 45.695 87.905 46.155 ;
        RECT 88.425 45.525 88.705 45.985 ;
        RECT 87.580 45.305 88.705 45.525 ;
        RECT 83.345 44.405 83.520 45.015 ;
        RECT 84.215 44.765 84.385 45.015 ;
        RECT 83.690 44.595 84.385 44.765 ;
        RECT 84.560 44.595 84.980 44.795 ;
        RECT 85.150 44.595 85.480 44.795 ;
        RECT 85.650 44.595 85.980 44.795 ;
        RECT 82.105 44.235 83.060 44.405 ;
        RECT 82.335 43.605 82.605 44.065 ;
        RECT 82.775 43.775 83.060 44.235 ;
        RECT 83.345 43.775 83.685 44.405 ;
        RECT 83.855 43.605 84.105 44.405 ;
        RECT 84.295 44.255 85.520 44.425 ;
        RECT 84.295 43.775 84.625 44.255 ;
        RECT 84.795 43.605 85.020 44.065 ;
        RECT 85.190 43.775 85.520 44.255 ;
        RECT 86.150 44.385 86.320 45.015 ;
        RECT 86.505 44.595 86.855 44.845 ;
        RECT 86.150 43.775 86.650 44.385 ;
        RECT 87.025 44.345 87.305 45.015 ;
        RECT 87.580 44.845 88.030 45.305 ;
        RECT 88.895 45.135 89.295 45.985 ;
        RECT 89.695 45.695 89.965 46.155 ;
        RECT 90.135 45.525 90.420 45.985 ;
        RECT 87.475 44.515 88.030 44.845 ;
        RECT 88.200 44.575 89.295 45.135 ;
        RECT 87.580 44.405 88.030 44.515 ;
        RECT 87.025 43.775 87.410 44.345 ;
        RECT 87.580 44.235 88.705 44.405 ;
        RECT 87.580 43.605 87.905 44.065 ;
        RECT 88.425 43.775 88.705 44.235 ;
        RECT 88.895 43.775 89.295 44.575 ;
        RECT 89.465 45.305 90.420 45.525 ;
        RECT 89.465 44.405 89.675 45.305 ;
        RECT 89.845 44.575 90.535 45.135 ;
        RECT 91.630 45.015 91.965 45.985 ;
        RECT 92.135 45.015 92.305 46.155 ;
        RECT 92.475 45.815 94.505 45.985 ;
        RECT 89.465 44.235 90.420 44.405 ;
        RECT 89.695 43.605 89.965 44.065 ;
        RECT 90.135 43.775 90.420 44.235 ;
        RECT 91.630 44.345 91.800 45.015 ;
        RECT 92.475 44.845 92.645 45.815 ;
        RECT 91.970 44.515 92.225 44.845 ;
        RECT 92.450 44.515 92.645 44.845 ;
        RECT 92.815 45.475 93.940 45.645 ;
        RECT 92.055 44.345 92.225 44.515 ;
        RECT 92.815 44.345 92.985 45.475 ;
        RECT 91.630 43.775 91.885 44.345 ;
        RECT 92.055 44.175 92.985 44.345 ;
        RECT 93.155 45.135 94.165 45.305 ;
        RECT 93.155 44.335 93.325 45.135 ;
        RECT 92.810 44.140 92.985 44.175 ;
        RECT 92.055 43.605 92.385 44.005 ;
        RECT 92.810 43.775 93.340 44.140 ;
        RECT 93.530 44.115 93.805 44.935 ;
        RECT 93.525 43.945 93.805 44.115 ;
        RECT 93.530 43.775 93.805 43.945 ;
        RECT 93.975 43.775 94.165 45.135 ;
        RECT 94.335 45.150 94.505 45.815 ;
        RECT 94.675 45.395 94.845 46.155 ;
        RECT 95.080 45.395 95.595 45.805 ;
        RECT 94.335 44.960 95.085 45.150 ;
        RECT 95.255 44.585 95.595 45.395 ;
        RECT 95.765 44.990 96.055 46.155 ;
        RECT 96.230 45.485 96.485 45.985 ;
        RECT 96.655 45.655 96.985 46.155 ;
        RECT 96.230 45.315 96.980 45.485 ;
        RECT 94.365 44.415 95.595 44.585 ;
        RECT 96.230 44.495 96.580 45.145 ;
        RECT 94.345 43.605 94.855 44.140 ;
        RECT 95.075 43.810 95.320 44.415 ;
        RECT 95.765 43.605 96.055 44.330 ;
        RECT 96.750 44.325 96.980 45.315 ;
        RECT 96.230 44.155 96.980 44.325 ;
        RECT 96.230 43.865 96.485 44.155 ;
        RECT 96.655 43.605 96.985 43.985 ;
        RECT 97.155 43.865 97.325 45.985 ;
        RECT 97.495 45.185 97.820 45.970 ;
        RECT 97.990 45.695 98.240 46.155 ;
        RECT 98.410 45.655 98.660 45.985 ;
        RECT 98.875 45.655 99.555 45.985 ;
        RECT 98.410 45.525 98.580 45.655 ;
        RECT 98.185 45.355 98.580 45.525 ;
        RECT 97.555 44.135 98.015 45.185 ;
        RECT 98.185 43.995 98.355 45.355 ;
        RECT 98.750 45.095 99.215 45.485 ;
        RECT 98.525 44.285 98.875 44.905 ;
        RECT 99.045 44.505 99.215 45.095 ;
        RECT 99.385 44.875 99.555 45.655 ;
        RECT 99.725 45.555 99.895 45.895 ;
        RECT 100.130 45.725 100.460 46.155 ;
        RECT 100.630 45.555 100.800 45.895 ;
        RECT 101.095 45.695 101.465 46.155 ;
        RECT 99.725 45.385 100.800 45.555 ;
        RECT 101.635 45.525 101.805 45.985 ;
        RECT 102.040 45.645 102.910 45.985 ;
        RECT 103.080 45.695 103.330 46.155 ;
        RECT 101.245 45.355 101.805 45.525 ;
        RECT 101.245 45.215 101.415 45.355 ;
        RECT 99.915 45.045 101.415 45.215 ;
        RECT 102.110 45.185 102.570 45.475 ;
        RECT 99.385 44.705 101.075 44.875 ;
        RECT 99.045 44.285 99.400 44.505 ;
        RECT 99.570 43.995 99.740 44.705 ;
        RECT 99.945 44.285 100.735 44.535 ;
        RECT 100.905 44.525 101.075 44.705 ;
        RECT 101.245 44.355 101.415 45.045 ;
        RECT 97.685 43.605 98.015 43.965 ;
        RECT 98.185 43.825 98.680 43.995 ;
        RECT 98.885 43.825 99.740 43.995 ;
        RECT 100.615 43.605 100.945 44.065 ;
        RECT 101.155 43.965 101.415 44.355 ;
        RECT 101.605 45.175 102.570 45.185 ;
        RECT 102.740 45.265 102.910 45.645 ;
        RECT 103.500 45.605 103.670 45.895 ;
        RECT 103.850 45.775 104.180 46.155 ;
        RECT 103.500 45.435 104.300 45.605 ;
        RECT 101.605 45.015 102.280 45.175 ;
        RECT 102.740 45.095 103.960 45.265 ;
        RECT 101.605 44.225 101.815 45.015 ;
        RECT 102.740 45.005 102.910 45.095 ;
        RECT 101.985 44.225 102.335 44.845 ;
        RECT 102.505 44.835 102.910 45.005 ;
        RECT 102.505 44.055 102.675 44.835 ;
        RECT 102.845 44.385 103.065 44.665 ;
        RECT 103.245 44.555 103.785 44.925 ;
        RECT 104.130 44.845 104.300 45.435 ;
        RECT 104.520 45.015 104.825 46.155 ;
        RECT 104.995 44.965 105.250 45.845 ;
        RECT 105.485 45.015 105.695 46.155 ;
        RECT 104.130 44.815 104.870 44.845 ;
        RECT 102.845 44.215 103.375 44.385 ;
        RECT 101.155 43.795 101.505 43.965 ;
        RECT 101.725 43.775 102.675 44.055 ;
        RECT 102.845 43.605 103.035 44.045 ;
        RECT 103.205 43.985 103.375 44.215 ;
        RECT 103.545 44.155 103.785 44.555 ;
        RECT 103.955 44.515 104.870 44.815 ;
        RECT 103.955 44.340 104.280 44.515 ;
        RECT 103.955 43.985 104.275 44.340 ;
        RECT 105.040 44.315 105.250 44.965 ;
        RECT 105.865 45.005 106.195 45.985 ;
        RECT 106.365 45.015 106.595 46.155 ;
        RECT 106.845 45.015 107.075 46.155 ;
        RECT 107.245 45.005 107.575 45.985 ;
        RECT 107.745 45.015 107.955 46.155 ;
        RECT 108.185 45.720 113.530 46.155 ;
        RECT 103.205 43.815 104.275 43.985 ;
        RECT 104.520 43.605 104.825 44.065 ;
        RECT 104.995 43.785 105.250 44.315 ;
        RECT 105.485 43.605 105.695 44.425 ;
        RECT 105.865 44.405 106.115 45.005 ;
        RECT 106.285 44.595 106.615 44.845 ;
        RECT 106.825 44.595 107.155 44.845 ;
        RECT 105.865 43.775 106.195 44.405 ;
        RECT 106.365 43.605 106.595 44.425 ;
        RECT 106.845 43.605 107.075 44.425 ;
        RECT 107.325 44.405 107.575 45.005 ;
        RECT 107.245 43.775 107.575 44.405 ;
        RECT 107.745 43.605 107.955 44.425 ;
        RECT 109.770 44.150 110.110 44.980 ;
        RECT 111.590 44.470 111.940 45.720 ;
        RECT 113.705 45.065 117.215 46.155 ;
        RECT 113.705 44.375 115.355 44.895 ;
        RECT 115.525 44.545 117.215 45.065 ;
        RECT 117.385 45.065 118.595 46.155 ;
        RECT 117.385 44.525 117.905 45.065 ;
        RECT 108.185 43.605 113.530 44.150 ;
        RECT 113.705 43.605 117.215 44.375 ;
        RECT 118.075 44.355 118.595 44.895 ;
        RECT 117.385 43.605 118.595 44.355 ;
        RECT 5.520 43.435 118.680 43.605 ;
        RECT 5.605 42.685 6.815 43.435 ;
        RECT 5.605 42.145 6.125 42.685 ;
        RECT 6.985 42.665 9.575 43.435 ;
        RECT 10.205 42.760 10.465 43.265 ;
        RECT 10.645 43.055 10.975 43.435 ;
        RECT 11.155 42.885 11.325 43.265 ;
        RECT 6.295 41.975 6.815 42.515 ;
        RECT 6.985 42.145 8.195 42.665 ;
        RECT 8.365 41.975 9.575 42.495 ;
        RECT 5.605 40.885 6.815 41.975 ;
        RECT 6.985 40.885 9.575 41.975 ;
        RECT 10.205 41.960 10.375 42.760 ;
        RECT 10.660 42.715 11.325 42.885 ;
        RECT 10.660 42.460 10.830 42.715 ;
        RECT 11.645 42.615 11.855 43.435 ;
        RECT 12.025 42.635 12.355 43.265 ;
        RECT 10.545 42.130 10.830 42.460 ;
        RECT 11.065 42.165 11.395 42.535 ;
        RECT 10.660 41.985 10.830 42.130 ;
        RECT 12.025 42.035 12.275 42.635 ;
        RECT 12.525 42.615 12.755 43.435 ;
        RECT 12.970 42.885 13.225 43.175 ;
        RECT 13.395 43.055 13.725 43.435 ;
        RECT 12.970 42.715 13.720 42.885 ;
        RECT 12.445 42.195 12.775 42.445 ;
        RECT 10.205 41.055 10.475 41.960 ;
        RECT 10.660 41.815 11.325 41.985 ;
        RECT 10.645 40.885 10.975 41.645 ;
        RECT 11.155 41.055 11.325 41.815 ;
        RECT 11.645 40.885 11.855 42.025 ;
        RECT 12.025 41.055 12.355 42.035 ;
        RECT 12.525 40.885 12.755 42.025 ;
        RECT 12.970 41.895 13.320 42.545 ;
        RECT 13.490 41.725 13.720 42.715 ;
        RECT 12.970 41.555 13.720 41.725 ;
        RECT 12.970 41.055 13.225 41.555 ;
        RECT 13.395 40.885 13.725 41.385 ;
        RECT 13.895 41.055 14.065 43.175 ;
        RECT 14.425 43.075 14.755 43.435 ;
        RECT 14.925 43.045 15.420 43.215 ;
        RECT 15.625 43.045 16.480 43.215 ;
        RECT 14.295 41.855 14.755 42.905 ;
        RECT 14.235 41.070 14.560 41.855 ;
        RECT 14.925 41.685 15.095 43.045 ;
        RECT 15.265 42.135 15.615 42.755 ;
        RECT 15.785 42.535 16.140 42.755 ;
        RECT 15.785 41.945 15.955 42.535 ;
        RECT 16.310 42.335 16.480 43.045 ;
        RECT 17.355 42.975 17.685 43.435 ;
        RECT 17.895 43.075 18.245 43.245 ;
        RECT 16.685 42.505 17.475 42.755 ;
        RECT 17.895 42.685 18.155 43.075 ;
        RECT 18.465 42.985 19.415 43.265 ;
        RECT 19.585 42.995 19.775 43.435 ;
        RECT 19.945 43.055 21.015 43.225 ;
        RECT 17.645 42.335 17.815 42.515 ;
        RECT 14.925 41.515 15.320 41.685 ;
        RECT 15.490 41.555 15.955 41.945 ;
        RECT 16.125 42.165 17.815 42.335 ;
        RECT 15.150 41.385 15.320 41.515 ;
        RECT 16.125 41.385 16.295 42.165 ;
        RECT 17.985 41.995 18.155 42.685 ;
        RECT 16.655 41.825 18.155 41.995 ;
        RECT 18.345 42.025 18.555 42.815 ;
        RECT 18.725 42.195 19.075 42.815 ;
        RECT 19.245 42.205 19.415 42.985 ;
        RECT 19.945 42.825 20.115 43.055 ;
        RECT 19.585 42.655 20.115 42.825 ;
        RECT 19.585 42.375 19.805 42.655 ;
        RECT 20.285 42.485 20.525 42.885 ;
        RECT 19.245 42.035 19.650 42.205 ;
        RECT 19.985 42.115 20.525 42.485 ;
        RECT 20.695 42.700 21.015 43.055 ;
        RECT 21.260 42.975 21.565 43.435 ;
        RECT 21.735 42.725 21.990 43.255 ;
        RECT 20.695 42.525 21.020 42.700 ;
        RECT 20.695 42.225 21.610 42.525 ;
        RECT 20.870 42.195 21.610 42.225 ;
        RECT 18.345 41.865 19.020 42.025 ;
        RECT 19.480 41.945 19.650 42.035 ;
        RECT 18.345 41.855 19.310 41.865 ;
        RECT 17.985 41.685 18.155 41.825 ;
        RECT 14.730 40.885 14.980 41.345 ;
        RECT 15.150 41.055 15.400 41.385 ;
        RECT 15.615 41.055 16.295 41.385 ;
        RECT 16.465 41.485 17.540 41.655 ;
        RECT 17.985 41.515 18.545 41.685 ;
        RECT 18.850 41.565 19.310 41.855 ;
        RECT 19.480 41.775 20.700 41.945 ;
        RECT 16.465 41.145 16.635 41.485 ;
        RECT 16.870 40.885 17.200 41.315 ;
        RECT 17.370 41.145 17.540 41.485 ;
        RECT 17.835 40.885 18.205 41.345 ;
        RECT 18.375 41.055 18.545 41.515 ;
        RECT 19.480 41.395 19.650 41.775 ;
        RECT 20.870 41.605 21.040 42.195 ;
        RECT 21.780 42.075 21.990 42.725 ;
        RECT 22.225 42.615 22.435 43.435 ;
        RECT 22.605 42.635 22.935 43.265 ;
        RECT 18.780 41.055 19.650 41.395 ;
        RECT 20.240 41.435 21.040 41.605 ;
        RECT 19.820 40.885 20.070 41.345 ;
        RECT 20.240 41.145 20.410 41.435 ;
        RECT 20.590 40.885 20.920 41.265 ;
        RECT 21.260 40.885 21.565 42.025 ;
        RECT 21.735 41.195 21.990 42.075 ;
        RECT 22.605 42.035 22.855 42.635 ;
        RECT 23.105 42.615 23.335 43.435 ;
        RECT 24.120 42.805 24.405 43.265 ;
        RECT 24.575 42.975 24.845 43.435 ;
        RECT 24.120 42.635 25.075 42.805 ;
        RECT 23.025 42.195 23.355 42.445 ;
        RECT 22.225 40.885 22.435 42.025 ;
        RECT 22.605 41.055 22.935 42.035 ;
        RECT 23.105 40.885 23.335 42.025 ;
        RECT 24.005 41.905 24.695 42.465 ;
        RECT 24.865 41.735 25.075 42.635 ;
        RECT 24.120 41.515 25.075 41.735 ;
        RECT 25.245 42.465 25.645 43.265 ;
        RECT 25.835 42.805 26.115 43.265 ;
        RECT 26.635 42.975 26.960 43.435 ;
        RECT 25.835 42.635 26.960 42.805 ;
        RECT 27.130 42.695 27.515 43.265 ;
        RECT 26.510 42.525 26.960 42.635 ;
        RECT 25.245 41.905 26.340 42.465 ;
        RECT 26.510 42.195 27.065 42.525 ;
        RECT 24.120 41.055 24.405 41.515 ;
        RECT 24.575 40.885 24.845 41.345 ;
        RECT 25.245 41.055 25.645 41.905 ;
        RECT 26.510 41.735 26.960 42.195 ;
        RECT 27.235 42.025 27.515 42.695 ;
        RECT 27.800 42.805 28.085 43.265 ;
        RECT 28.255 42.975 28.525 43.435 ;
        RECT 27.800 42.635 28.755 42.805 ;
        RECT 25.835 41.515 26.960 41.735 ;
        RECT 25.835 41.055 26.115 41.515 ;
        RECT 26.635 40.885 26.960 41.345 ;
        RECT 27.130 41.055 27.515 42.025 ;
        RECT 27.685 41.905 28.375 42.465 ;
        RECT 28.545 41.735 28.755 42.635 ;
        RECT 27.800 41.515 28.755 41.735 ;
        RECT 28.925 42.465 29.325 43.265 ;
        RECT 29.515 42.805 29.795 43.265 ;
        RECT 30.315 42.975 30.640 43.435 ;
        RECT 29.515 42.635 30.640 42.805 ;
        RECT 30.810 42.695 31.195 43.265 ;
        RECT 31.365 42.710 31.655 43.435 ;
        RECT 31.830 42.885 32.085 43.175 ;
        RECT 32.255 43.055 32.585 43.435 ;
        RECT 31.830 42.715 32.580 42.885 ;
        RECT 30.190 42.525 30.640 42.635 ;
        RECT 28.925 41.905 30.020 42.465 ;
        RECT 30.190 42.195 30.745 42.525 ;
        RECT 27.800 41.055 28.085 41.515 ;
        RECT 28.255 40.885 28.525 41.345 ;
        RECT 28.925 41.055 29.325 41.905 ;
        RECT 30.190 41.735 30.640 42.195 ;
        RECT 30.915 42.025 31.195 42.695 ;
        RECT 29.515 41.515 30.640 41.735 ;
        RECT 29.515 41.055 29.795 41.515 ;
        RECT 30.315 40.885 30.640 41.345 ;
        RECT 30.810 41.055 31.195 42.025 ;
        RECT 31.365 40.885 31.655 42.050 ;
        RECT 31.830 41.895 32.180 42.545 ;
        RECT 32.350 41.725 32.580 42.715 ;
        RECT 31.830 41.555 32.580 41.725 ;
        RECT 31.830 41.055 32.085 41.555 ;
        RECT 32.255 40.885 32.585 41.385 ;
        RECT 32.755 41.055 32.925 43.175 ;
        RECT 33.285 43.075 33.615 43.435 ;
        RECT 33.785 43.045 34.280 43.215 ;
        RECT 34.485 43.045 35.340 43.215 ;
        RECT 33.155 41.855 33.615 42.905 ;
        RECT 33.095 41.070 33.420 41.855 ;
        RECT 33.785 41.685 33.955 43.045 ;
        RECT 34.125 42.135 34.475 42.755 ;
        RECT 34.645 42.535 35.000 42.755 ;
        RECT 34.645 41.945 34.815 42.535 ;
        RECT 35.170 42.335 35.340 43.045 ;
        RECT 36.215 42.975 36.545 43.435 ;
        RECT 36.755 43.075 37.105 43.245 ;
        RECT 35.545 42.505 36.335 42.755 ;
        RECT 36.755 42.685 37.015 43.075 ;
        RECT 37.325 42.985 38.275 43.265 ;
        RECT 38.445 42.995 38.635 43.435 ;
        RECT 38.805 43.055 39.875 43.225 ;
        RECT 36.505 42.335 36.675 42.515 ;
        RECT 33.785 41.515 34.180 41.685 ;
        RECT 34.350 41.555 34.815 41.945 ;
        RECT 34.985 42.165 36.675 42.335 ;
        RECT 34.010 41.385 34.180 41.515 ;
        RECT 34.985 41.385 35.155 42.165 ;
        RECT 36.845 41.995 37.015 42.685 ;
        RECT 35.515 41.825 37.015 41.995 ;
        RECT 37.205 42.025 37.415 42.815 ;
        RECT 37.585 42.195 37.935 42.815 ;
        RECT 38.105 42.205 38.275 42.985 ;
        RECT 38.805 42.825 38.975 43.055 ;
        RECT 38.445 42.655 38.975 42.825 ;
        RECT 38.445 42.375 38.665 42.655 ;
        RECT 39.145 42.485 39.385 42.885 ;
        RECT 38.105 42.035 38.510 42.205 ;
        RECT 38.845 42.115 39.385 42.485 ;
        RECT 39.555 42.700 39.875 43.055 ;
        RECT 40.120 42.975 40.425 43.435 ;
        RECT 40.595 42.725 40.850 43.255 ;
        RECT 39.555 42.525 39.880 42.700 ;
        RECT 39.555 42.225 40.470 42.525 ;
        RECT 39.730 42.195 40.470 42.225 ;
        RECT 37.205 41.865 37.880 42.025 ;
        RECT 38.340 41.945 38.510 42.035 ;
        RECT 37.205 41.855 38.170 41.865 ;
        RECT 36.845 41.685 37.015 41.825 ;
        RECT 33.590 40.885 33.840 41.345 ;
        RECT 34.010 41.055 34.260 41.385 ;
        RECT 34.475 41.055 35.155 41.385 ;
        RECT 35.325 41.485 36.400 41.655 ;
        RECT 36.845 41.515 37.405 41.685 ;
        RECT 37.710 41.565 38.170 41.855 ;
        RECT 38.340 41.775 39.560 41.945 ;
        RECT 35.325 41.145 35.495 41.485 ;
        RECT 35.730 40.885 36.060 41.315 ;
        RECT 36.230 41.145 36.400 41.485 ;
        RECT 36.695 40.885 37.065 41.345 ;
        RECT 37.235 41.055 37.405 41.515 ;
        RECT 38.340 41.395 38.510 41.775 ;
        RECT 39.730 41.605 39.900 42.195 ;
        RECT 40.640 42.075 40.850 42.725 ;
        RECT 41.085 42.615 41.295 43.435 ;
        RECT 41.465 42.635 41.795 43.265 ;
        RECT 37.640 41.055 38.510 41.395 ;
        RECT 39.100 41.435 39.900 41.605 ;
        RECT 38.680 40.885 38.930 41.345 ;
        RECT 39.100 41.145 39.270 41.435 ;
        RECT 39.450 40.885 39.780 41.265 ;
        RECT 40.120 40.885 40.425 42.025 ;
        RECT 40.595 41.195 40.850 42.075 ;
        RECT 41.465 42.035 41.715 42.635 ;
        RECT 41.965 42.615 42.195 43.435 ;
        RECT 42.495 42.885 42.665 43.265 ;
        RECT 42.845 43.055 43.175 43.435 ;
        RECT 42.495 42.715 43.160 42.885 ;
        RECT 43.355 42.760 43.615 43.265 ;
        RECT 41.885 42.195 42.215 42.445 ;
        RECT 42.425 42.165 42.755 42.535 ;
        RECT 42.990 42.460 43.160 42.715 ;
        RECT 42.990 42.130 43.275 42.460 ;
        RECT 41.085 40.885 41.295 42.025 ;
        RECT 41.465 41.055 41.795 42.035 ;
        RECT 41.965 40.885 42.195 42.025 ;
        RECT 42.990 41.985 43.160 42.130 ;
        RECT 42.495 41.815 43.160 41.985 ;
        RECT 43.445 41.960 43.615 42.760 ;
        RECT 42.495 41.055 42.665 41.815 ;
        RECT 42.845 40.885 43.175 41.645 ;
        RECT 43.345 41.055 43.615 41.960 ;
        RECT 43.790 42.695 44.045 43.265 ;
        RECT 44.215 43.035 44.545 43.435 ;
        RECT 44.970 42.900 45.500 43.265 ;
        RECT 45.690 43.095 45.965 43.265 ;
        RECT 45.685 42.925 45.965 43.095 ;
        RECT 44.970 42.865 45.145 42.900 ;
        RECT 44.215 42.695 45.145 42.865 ;
        RECT 43.790 42.025 43.960 42.695 ;
        RECT 44.215 42.525 44.385 42.695 ;
        RECT 44.130 42.195 44.385 42.525 ;
        RECT 44.610 42.195 44.805 42.525 ;
        RECT 43.790 41.055 44.125 42.025 ;
        RECT 44.295 40.885 44.465 42.025 ;
        RECT 44.635 41.225 44.805 42.195 ;
        RECT 44.975 41.565 45.145 42.695 ;
        RECT 45.315 41.905 45.485 42.705 ;
        RECT 45.690 42.105 45.965 42.925 ;
        RECT 46.135 41.905 46.325 43.265 ;
        RECT 46.505 42.900 47.015 43.435 ;
        RECT 47.235 42.625 47.480 43.230 ;
        RECT 47.925 42.665 49.595 43.435 ;
        RECT 46.525 42.455 47.755 42.625 ;
        RECT 45.315 41.735 46.325 41.905 ;
        RECT 46.495 41.890 47.245 42.080 ;
        RECT 44.975 41.395 46.100 41.565 ;
        RECT 46.495 41.225 46.665 41.890 ;
        RECT 47.415 41.645 47.755 42.455 ;
        RECT 47.925 42.145 48.675 42.665 ;
        RECT 49.765 42.635 50.105 43.265 ;
        RECT 50.275 42.635 50.525 43.435 ;
        RECT 50.715 42.785 51.045 43.265 ;
        RECT 51.215 42.975 51.440 43.435 ;
        RECT 51.610 42.785 51.940 43.265 ;
        RECT 48.845 41.975 49.595 42.495 ;
        RECT 44.635 41.055 46.665 41.225 ;
        RECT 46.835 40.885 47.005 41.645 ;
        RECT 47.240 41.235 47.755 41.645 ;
        RECT 47.925 40.885 49.595 41.975 ;
        RECT 49.765 42.025 49.940 42.635 ;
        RECT 50.715 42.615 51.940 42.785 ;
        RECT 52.570 42.655 53.070 43.265 ;
        RECT 53.445 42.695 53.830 43.265 ;
        RECT 54.000 42.975 54.325 43.435 ;
        RECT 54.845 42.805 55.125 43.265 ;
        RECT 50.110 42.275 50.805 42.445 ;
        RECT 50.635 42.025 50.805 42.275 ;
        RECT 50.980 42.245 51.400 42.445 ;
        RECT 51.570 42.245 51.900 42.445 ;
        RECT 52.070 42.245 52.400 42.445 ;
        RECT 52.570 42.025 52.740 42.655 ;
        RECT 52.925 42.195 53.275 42.445 ;
        RECT 53.445 42.025 53.725 42.695 ;
        RECT 54.000 42.635 55.125 42.805 ;
        RECT 54.000 42.525 54.450 42.635 ;
        RECT 53.895 42.195 54.450 42.525 ;
        RECT 55.315 42.465 55.715 43.265 ;
        RECT 56.115 42.975 56.385 43.435 ;
        RECT 56.555 42.805 56.840 43.265 ;
        RECT 49.765 41.055 50.105 42.025 ;
        RECT 50.275 40.885 50.445 42.025 ;
        RECT 50.635 41.855 53.070 42.025 ;
        RECT 50.715 40.885 50.965 41.685 ;
        RECT 51.610 41.055 51.940 41.855 ;
        RECT 52.240 40.885 52.570 41.685 ;
        RECT 52.740 41.055 53.070 41.855 ;
        RECT 53.445 41.055 53.830 42.025 ;
        RECT 54.000 41.735 54.450 42.195 ;
        RECT 54.620 41.905 55.715 42.465 ;
        RECT 54.000 41.515 55.125 41.735 ;
        RECT 54.000 40.885 54.325 41.345 ;
        RECT 54.845 41.055 55.125 41.515 ;
        RECT 55.315 41.055 55.715 41.905 ;
        RECT 55.885 42.635 56.840 42.805 ;
        RECT 57.125 42.710 57.415 43.435 ;
        RECT 58.810 42.865 58.980 43.115 ;
        RECT 58.505 42.695 58.980 42.865 ;
        RECT 59.215 42.695 59.545 43.435 ;
        RECT 59.715 42.865 59.915 43.210 ;
        RECT 60.085 43.035 60.415 43.435 ;
        RECT 60.585 42.865 60.785 43.220 ;
        RECT 60.955 43.040 61.285 43.435 ;
        RECT 61.785 42.955 62.065 43.435 ;
        RECT 59.715 42.695 61.555 42.865 ;
        RECT 62.235 42.785 62.495 43.175 ;
        RECT 62.670 42.955 62.925 43.435 ;
        RECT 63.095 42.785 63.390 43.175 ;
        RECT 63.570 42.955 63.845 43.435 ;
        RECT 64.015 42.935 64.315 43.265 ;
        RECT 55.885 41.735 56.095 42.635 ;
        RECT 56.265 41.905 56.955 42.465 ;
        RECT 55.885 41.515 56.840 41.735 ;
        RECT 56.115 40.885 56.385 41.345 ;
        RECT 56.555 41.055 56.840 41.515 ;
        RECT 57.125 40.885 57.415 42.050 ;
        RECT 58.505 41.725 58.675 42.695 ;
        RECT 58.845 41.905 59.195 42.525 ;
        RECT 59.365 41.905 59.685 42.525 ;
        RECT 59.855 41.905 60.185 42.525 ;
        RECT 60.355 41.905 60.655 42.525 ;
        RECT 60.895 41.725 61.115 42.525 ;
        RECT 58.505 41.515 61.115 41.725 ;
        RECT 59.215 40.885 59.545 41.335 ;
        RECT 61.295 41.070 61.555 42.695 ;
        RECT 61.740 42.615 63.390 42.785 ;
        RECT 61.740 42.105 62.145 42.615 ;
        RECT 62.315 42.275 63.455 42.445 ;
        RECT 61.740 41.935 62.495 42.105 ;
        RECT 61.780 40.885 62.065 41.755 ;
        RECT 62.235 41.685 62.495 41.935 ;
        RECT 63.285 42.025 63.455 42.275 ;
        RECT 63.625 42.195 63.975 42.765 ;
        RECT 64.145 42.025 64.315 42.935 ;
        RECT 64.575 42.885 64.745 43.265 ;
        RECT 64.960 43.055 65.290 43.435 ;
        RECT 64.575 42.715 65.290 42.885 ;
        RECT 64.485 42.165 64.840 42.535 ;
        RECT 65.120 42.525 65.290 42.715 ;
        RECT 65.460 42.690 65.715 43.265 ;
        RECT 65.120 42.195 65.375 42.525 ;
        RECT 63.285 41.855 64.315 42.025 ;
        RECT 65.120 41.985 65.290 42.195 ;
        RECT 62.235 41.515 63.355 41.685 ;
        RECT 62.235 41.055 62.495 41.515 ;
        RECT 62.670 40.885 62.925 41.345 ;
        RECT 63.095 41.055 63.355 41.515 ;
        RECT 63.525 40.885 63.835 41.685 ;
        RECT 64.005 41.055 64.315 41.855 ;
        RECT 64.575 41.815 65.290 41.985 ;
        RECT 65.545 41.960 65.715 42.690 ;
        RECT 65.890 42.595 66.150 43.435 ;
        RECT 66.385 42.615 66.595 43.435 ;
        RECT 66.765 42.635 67.095 43.265 ;
        RECT 66.765 42.035 67.015 42.635 ;
        RECT 67.265 42.615 67.495 43.435 ;
        RECT 67.705 42.665 70.295 43.435 ;
        RECT 70.465 42.935 70.765 43.265 ;
        RECT 70.935 42.955 71.210 43.435 ;
        RECT 67.185 42.195 67.515 42.445 ;
        RECT 67.705 42.145 68.915 42.665 ;
        RECT 64.575 41.055 64.745 41.815 ;
        RECT 64.960 40.885 65.290 41.645 ;
        RECT 65.460 41.055 65.715 41.960 ;
        RECT 65.890 40.885 66.150 42.035 ;
        RECT 66.385 40.885 66.595 42.025 ;
        RECT 66.765 41.055 67.095 42.035 ;
        RECT 67.265 40.885 67.495 42.025 ;
        RECT 69.085 41.975 70.295 42.495 ;
        RECT 67.705 40.885 70.295 41.975 ;
        RECT 70.465 42.025 70.635 42.935 ;
        RECT 71.390 42.785 71.685 43.175 ;
        RECT 71.855 42.955 72.110 43.435 ;
        RECT 72.285 42.785 72.545 43.175 ;
        RECT 72.715 42.955 72.995 43.435 ;
        RECT 70.805 42.195 71.155 42.765 ;
        RECT 71.390 42.615 73.040 42.785 ;
        RECT 73.500 42.625 73.745 43.230 ;
        RECT 73.965 42.900 74.475 43.435 ;
        RECT 71.325 42.275 72.465 42.445 ;
        RECT 71.325 42.025 71.495 42.275 ;
        RECT 72.635 42.105 73.040 42.615 ;
        RECT 70.465 41.855 71.495 42.025 ;
        RECT 72.285 41.935 73.040 42.105 ;
        RECT 73.225 42.455 74.455 42.625 ;
        RECT 70.465 41.055 70.775 41.855 ;
        RECT 72.285 41.685 72.545 41.935 ;
        RECT 70.945 40.885 71.255 41.685 ;
        RECT 71.425 41.515 72.545 41.685 ;
        RECT 71.425 41.055 71.685 41.515 ;
        RECT 71.855 40.885 72.110 41.345 ;
        RECT 72.285 41.055 72.545 41.515 ;
        RECT 72.715 40.885 73.000 41.755 ;
        RECT 73.225 41.645 73.565 42.455 ;
        RECT 73.735 41.890 74.485 42.080 ;
        RECT 73.225 41.235 73.740 41.645 ;
        RECT 73.975 40.885 74.145 41.645 ;
        RECT 74.315 41.225 74.485 41.890 ;
        RECT 74.655 41.905 74.845 43.265 ;
        RECT 75.015 43.095 75.290 43.265 ;
        RECT 75.015 42.925 75.295 43.095 ;
        RECT 75.015 42.105 75.290 42.925 ;
        RECT 75.480 42.900 76.010 43.265 ;
        RECT 76.435 43.035 76.765 43.435 ;
        RECT 75.835 42.865 76.010 42.900 ;
        RECT 75.495 41.905 75.665 42.705 ;
        RECT 74.655 41.735 75.665 41.905 ;
        RECT 75.835 42.695 76.765 42.865 ;
        RECT 76.935 42.695 77.190 43.265 ;
        RECT 75.835 41.565 76.005 42.695 ;
        RECT 76.595 42.525 76.765 42.695 ;
        RECT 74.880 41.395 76.005 41.565 ;
        RECT 76.175 42.195 76.370 42.525 ;
        RECT 76.595 42.195 76.850 42.525 ;
        RECT 76.175 41.225 76.345 42.195 ;
        RECT 77.020 42.025 77.190 42.695 ;
        RECT 77.365 42.665 79.035 43.435 ;
        RECT 79.205 42.695 79.590 43.265 ;
        RECT 79.760 42.975 80.085 43.435 ;
        RECT 80.605 42.805 80.885 43.265 ;
        RECT 77.365 42.145 78.115 42.665 ;
        RECT 74.315 41.055 76.345 41.225 ;
        RECT 76.515 40.885 76.685 42.025 ;
        RECT 76.855 41.055 77.190 42.025 ;
        RECT 78.285 41.975 79.035 42.495 ;
        RECT 77.365 40.885 79.035 41.975 ;
        RECT 79.205 42.025 79.485 42.695 ;
        RECT 79.760 42.635 80.885 42.805 ;
        RECT 79.760 42.525 80.210 42.635 ;
        RECT 79.655 42.195 80.210 42.525 ;
        RECT 81.075 42.465 81.475 43.265 ;
        RECT 81.875 42.975 82.145 43.435 ;
        RECT 82.315 42.805 82.600 43.265 ;
        RECT 79.205 41.055 79.590 42.025 ;
        RECT 79.760 41.735 80.210 42.195 ;
        RECT 80.380 41.905 81.475 42.465 ;
        RECT 79.760 41.515 80.885 41.735 ;
        RECT 79.760 40.885 80.085 41.345 ;
        RECT 80.605 41.055 80.885 41.515 ;
        RECT 81.075 41.055 81.475 41.905 ;
        RECT 81.645 42.635 82.600 42.805 ;
        RECT 82.885 42.710 83.175 43.435 ;
        RECT 83.350 42.695 83.605 43.265 ;
        RECT 83.775 43.035 84.105 43.435 ;
        RECT 84.530 42.900 85.060 43.265 ;
        RECT 85.250 43.095 85.525 43.265 ;
        RECT 85.245 42.925 85.525 43.095 ;
        RECT 84.530 42.865 84.705 42.900 ;
        RECT 83.775 42.695 84.705 42.865 ;
        RECT 81.645 41.735 81.855 42.635 ;
        RECT 82.025 41.905 82.715 42.465 ;
        RECT 81.645 41.515 82.600 41.735 ;
        RECT 81.875 40.885 82.145 41.345 ;
        RECT 82.315 41.055 82.600 41.515 ;
        RECT 82.885 40.885 83.175 42.050 ;
        RECT 83.350 42.025 83.520 42.695 ;
        RECT 83.775 42.525 83.945 42.695 ;
        RECT 83.690 42.195 83.945 42.525 ;
        RECT 84.170 42.195 84.365 42.525 ;
        RECT 83.350 41.055 83.685 42.025 ;
        RECT 83.855 40.885 84.025 42.025 ;
        RECT 84.195 41.225 84.365 42.195 ;
        RECT 84.535 41.565 84.705 42.695 ;
        RECT 84.875 41.905 85.045 42.705 ;
        RECT 85.250 42.105 85.525 42.925 ;
        RECT 85.695 41.905 85.885 43.265 ;
        RECT 86.065 42.900 86.575 43.435 ;
        RECT 86.795 42.625 87.040 43.230 ;
        RECT 87.690 42.655 88.190 43.265 ;
        RECT 86.085 42.455 87.315 42.625 ;
        RECT 84.875 41.735 85.885 41.905 ;
        RECT 86.055 41.890 86.805 42.080 ;
        RECT 84.535 41.395 85.660 41.565 ;
        RECT 86.055 41.225 86.225 41.890 ;
        RECT 86.975 41.645 87.315 42.455 ;
        RECT 87.485 42.195 87.835 42.445 ;
        RECT 88.020 42.025 88.190 42.655 ;
        RECT 88.820 42.785 89.150 43.265 ;
        RECT 89.320 42.975 89.545 43.435 ;
        RECT 89.715 42.785 90.045 43.265 ;
        RECT 88.820 42.615 90.045 42.785 ;
        RECT 90.235 42.635 90.485 43.435 ;
        RECT 90.655 42.635 90.995 43.265 ;
        RECT 91.830 42.655 92.330 43.265 ;
        RECT 88.360 42.245 88.690 42.445 ;
        RECT 88.860 42.245 89.190 42.445 ;
        RECT 89.360 42.245 89.780 42.445 ;
        RECT 89.955 42.275 90.650 42.445 ;
        RECT 89.955 42.025 90.125 42.275 ;
        RECT 90.820 42.025 90.995 42.635 ;
        RECT 91.625 42.195 91.975 42.445 ;
        RECT 92.160 42.025 92.330 42.655 ;
        RECT 92.960 42.785 93.290 43.265 ;
        RECT 93.460 42.975 93.685 43.435 ;
        RECT 93.855 42.785 94.185 43.265 ;
        RECT 92.960 42.615 94.185 42.785 ;
        RECT 94.375 42.635 94.625 43.435 ;
        RECT 94.795 42.635 95.135 43.265 ;
        RECT 95.880 42.805 96.165 43.265 ;
        RECT 96.335 42.975 96.605 43.435 ;
        RECT 95.880 42.635 96.835 42.805 ;
        RECT 94.905 42.585 95.135 42.635 ;
        RECT 92.500 42.245 92.830 42.445 ;
        RECT 93.000 42.245 93.330 42.445 ;
        RECT 93.500 42.245 93.920 42.445 ;
        RECT 94.095 42.275 94.790 42.445 ;
        RECT 94.095 42.025 94.265 42.275 ;
        RECT 94.960 42.025 95.135 42.585 ;
        RECT 84.195 41.055 86.225 41.225 ;
        RECT 86.395 40.885 86.565 41.645 ;
        RECT 86.800 41.235 87.315 41.645 ;
        RECT 87.690 41.855 90.125 42.025 ;
        RECT 87.690 41.055 88.020 41.855 ;
        RECT 88.190 40.885 88.520 41.685 ;
        RECT 88.820 41.055 89.150 41.855 ;
        RECT 89.795 40.885 90.045 41.685 ;
        RECT 90.315 40.885 90.485 42.025 ;
        RECT 90.655 41.055 90.995 42.025 ;
        RECT 91.830 41.855 94.265 42.025 ;
        RECT 91.830 41.055 92.160 41.855 ;
        RECT 92.330 40.885 92.660 41.685 ;
        RECT 92.960 41.055 93.290 41.855 ;
        RECT 93.935 40.885 94.185 41.685 ;
        RECT 94.455 40.885 94.625 42.025 ;
        RECT 94.795 41.055 95.135 42.025 ;
        RECT 95.765 41.905 96.455 42.465 ;
        RECT 96.625 41.735 96.835 42.635 ;
        RECT 95.880 41.515 96.835 41.735 ;
        RECT 97.005 42.465 97.405 43.265 ;
        RECT 97.595 42.805 97.875 43.265 ;
        RECT 98.395 42.975 98.720 43.435 ;
        RECT 97.595 42.635 98.720 42.805 ;
        RECT 98.890 42.695 99.275 43.265 ;
        RECT 98.270 42.525 98.720 42.635 ;
        RECT 97.005 41.905 98.100 42.465 ;
        RECT 98.270 42.195 98.825 42.525 ;
        RECT 95.880 41.055 96.165 41.515 ;
        RECT 96.335 40.885 96.605 41.345 ;
        RECT 97.005 41.055 97.405 41.905 ;
        RECT 98.270 41.735 98.720 42.195 ;
        RECT 98.995 42.025 99.275 42.695 ;
        RECT 97.595 41.515 98.720 41.735 ;
        RECT 97.595 41.055 97.875 41.515 ;
        RECT 98.395 40.885 98.720 41.345 ;
        RECT 98.890 41.055 99.275 42.025 ;
        RECT 99.450 42.725 99.705 43.255 ;
        RECT 99.875 42.975 100.180 43.435 ;
        RECT 100.425 43.055 101.495 43.225 ;
        RECT 99.450 42.075 99.660 42.725 ;
        RECT 100.425 42.700 100.745 43.055 ;
        RECT 100.420 42.525 100.745 42.700 ;
        RECT 99.830 42.225 100.745 42.525 ;
        RECT 100.915 42.485 101.155 42.885 ;
        RECT 101.325 42.825 101.495 43.055 ;
        RECT 101.665 42.995 101.855 43.435 ;
        RECT 102.025 42.985 102.975 43.265 ;
        RECT 103.195 43.075 103.545 43.245 ;
        RECT 101.325 42.655 101.855 42.825 ;
        RECT 99.830 42.195 100.570 42.225 ;
        RECT 99.450 41.195 99.705 42.075 ;
        RECT 99.875 40.885 100.180 42.025 ;
        RECT 100.400 41.605 100.570 42.195 ;
        RECT 100.915 42.115 101.455 42.485 ;
        RECT 101.635 42.375 101.855 42.655 ;
        RECT 102.025 42.205 102.195 42.985 ;
        RECT 101.790 42.035 102.195 42.205 ;
        RECT 102.365 42.195 102.715 42.815 ;
        RECT 101.790 41.945 101.960 42.035 ;
        RECT 102.885 42.025 103.095 42.815 ;
        RECT 100.740 41.775 101.960 41.945 ;
        RECT 102.420 41.865 103.095 42.025 ;
        RECT 100.400 41.435 101.200 41.605 ;
        RECT 100.520 40.885 100.850 41.265 ;
        RECT 101.030 41.145 101.200 41.435 ;
        RECT 101.790 41.395 101.960 41.775 ;
        RECT 102.130 41.855 103.095 41.865 ;
        RECT 103.285 42.685 103.545 43.075 ;
        RECT 103.755 42.975 104.085 43.435 ;
        RECT 104.960 43.045 105.815 43.215 ;
        RECT 106.020 43.045 106.515 43.215 ;
        RECT 106.685 43.075 107.015 43.435 ;
        RECT 103.285 41.995 103.455 42.685 ;
        RECT 103.625 42.335 103.795 42.515 ;
        RECT 103.965 42.505 104.755 42.755 ;
        RECT 104.960 42.335 105.130 43.045 ;
        RECT 105.300 42.535 105.655 42.755 ;
        RECT 103.625 42.165 105.315 42.335 ;
        RECT 102.130 41.565 102.590 41.855 ;
        RECT 103.285 41.825 104.785 41.995 ;
        RECT 103.285 41.685 103.455 41.825 ;
        RECT 102.895 41.515 103.455 41.685 ;
        RECT 101.370 40.885 101.620 41.345 ;
        RECT 101.790 41.055 102.660 41.395 ;
        RECT 102.895 41.055 103.065 41.515 ;
        RECT 103.900 41.485 104.975 41.655 ;
        RECT 103.235 40.885 103.605 41.345 ;
        RECT 103.900 41.145 104.070 41.485 ;
        RECT 104.240 40.885 104.570 41.315 ;
        RECT 104.805 41.145 104.975 41.485 ;
        RECT 105.145 41.385 105.315 42.165 ;
        RECT 105.485 41.945 105.655 42.535 ;
        RECT 105.825 42.135 106.175 42.755 ;
        RECT 105.485 41.555 105.950 41.945 ;
        RECT 106.345 41.685 106.515 43.045 ;
        RECT 106.685 41.855 107.145 42.905 ;
        RECT 106.120 41.515 106.515 41.685 ;
        RECT 106.120 41.385 106.290 41.515 ;
        RECT 105.145 41.055 105.825 41.385 ;
        RECT 106.040 41.055 106.290 41.385 ;
        RECT 106.460 40.885 106.710 41.345 ;
        RECT 106.880 41.070 107.205 41.855 ;
        RECT 107.375 41.055 107.545 43.175 ;
        RECT 107.715 43.055 108.045 43.435 ;
        RECT 108.215 42.885 108.470 43.175 ;
        RECT 107.720 42.715 108.470 42.885 ;
        RECT 107.720 41.725 107.950 42.715 ;
        RECT 108.645 42.710 108.935 43.435 ;
        RECT 109.105 42.890 114.450 43.435 ;
        RECT 108.120 41.895 108.470 42.545 ;
        RECT 110.690 42.060 111.030 42.890 ;
        RECT 114.625 42.665 117.215 43.435 ;
        RECT 117.385 42.685 118.595 43.435 ;
        RECT 107.720 41.555 108.470 41.725 ;
        RECT 107.715 40.885 108.045 41.385 ;
        RECT 108.215 41.055 108.470 41.555 ;
        RECT 108.645 40.885 108.935 42.050 ;
        RECT 112.510 41.320 112.860 42.570 ;
        RECT 114.625 42.145 115.835 42.665 ;
        RECT 116.005 41.975 117.215 42.495 ;
        RECT 109.105 40.885 114.450 41.320 ;
        RECT 114.625 40.885 117.215 41.975 ;
        RECT 117.385 41.975 117.905 42.515 ;
        RECT 118.075 42.145 118.595 42.685 ;
        RECT 117.385 40.885 118.595 41.975 ;
        RECT 5.520 40.715 118.680 40.885 ;
        RECT 5.605 39.625 6.815 40.715 ;
        RECT 6.985 39.625 8.195 40.715 ;
        RECT 8.370 40.045 8.625 40.545 ;
        RECT 8.795 40.215 9.125 40.715 ;
        RECT 8.370 39.875 9.120 40.045 ;
        RECT 5.605 38.915 6.125 39.455 ;
        RECT 6.295 39.085 6.815 39.625 ;
        RECT 6.985 38.915 7.505 39.455 ;
        RECT 7.675 39.085 8.195 39.625 ;
        RECT 8.370 39.055 8.720 39.705 ;
        RECT 5.605 38.165 6.815 38.915 ;
        RECT 6.985 38.165 8.195 38.915 ;
        RECT 8.890 38.885 9.120 39.875 ;
        RECT 8.370 38.715 9.120 38.885 ;
        RECT 8.370 38.425 8.625 38.715 ;
        RECT 8.795 38.165 9.125 38.545 ;
        RECT 9.295 38.425 9.465 40.545 ;
        RECT 9.635 39.745 9.960 40.530 ;
        RECT 10.130 40.255 10.380 40.715 ;
        RECT 10.550 40.215 10.800 40.545 ;
        RECT 11.015 40.215 11.695 40.545 ;
        RECT 10.550 40.085 10.720 40.215 ;
        RECT 10.325 39.915 10.720 40.085 ;
        RECT 9.695 38.695 10.155 39.745 ;
        RECT 10.325 38.555 10.495 39.915 ;
        RECT 10.890 39.655 11.355 40.045 ;
        RECT 10.665 38.845 11.015 39.465 ;
        RECT 11.185 39.065 11.355 39.655 ;
        RECT 11.525 39.435 11.695 40.215 ;
        RECT 11.865 40.115 12.035 40.455 ;
        RECT 12.270 40.285 12.600 40.715 ;
        RECT 12.770 40.115 12.940 40.455 ;
        RECT 13.235 40.255 13.605 40.715 ;
        RECT 11.865 39.945 12.940 40.115 ;
        RECT 13.775 40.085 13.945 40.545 ;
        RECT 14.180 40.205 15.050 40.545 ;
        RECT 15.220 40.255 15.470 40.715 ;
        RECT 13.385 39.915 13.945 40.085 ;
        RECT 13.385 39.775 13.555 39.915 ;
        RECT 12.055 39.605 13.555 39.775 ;
        RECT 14.250 39.745 14.710 40.035 ;
        RECT 11.525 39.265 13.215 39.435 ;
        RECT 11.185 38.845 11.540 39.065 ;
        RECT 11.710 38.555 11.880 39.265 ;
        RECT 12.085 38.845 12.875 39.095 ;
        RECT 13.045 39.085 13.215 39.265 ;
        RECT 13.385 38.915 13.555 39.605 ;
        RECT 9.825 38.165 10.155 38.525 ;
        RECT 10.325 38.385 10.820 38.555 ;
        RECT 11.025 38.385 11.880 38.555 ;
        RECT 12.755 38.165 13.085 38.625 ;
        RECT 13.295 38.525 13.555 38.915 ;
        RECT 13.745 39.735 14.710 39.745 ;
        RECT 14.880 39.825 15.050 40.205 ;
        RECT 15.640 40.165 15.810 40.455 ;
        RECT 15.990 40.335 16.320 40.715 ;
        RECT 15.640 39.995 16.440 40.165 ;
        RECT 13.745 39.575 14.420 39.735 ;
        RECT 14.880 39.655 16.100 39.825 ;
        RECT 13.745 38.785 13.955 39.575 ;
        RECT 14.880 39.565 15.050 39.655 ;
        RECT 14.125 38.785 14.475 39.405 ;
        RECT 14.645 39.395 15.050 39.565 ;
        RECT 14.645 38.615 14.815 39.395 ;
        RECT 14.985 38.945 15.205 39.225 ;
        RECT 15.385 39.115 15.925 39.485 ;
        RECT 16.270 39.405 16.440 39.995 ;
        RECT 16.660 39.575 16.965 40.715 ;
        RECT 17.135 39.525 17.390 40.405 ;
        RECT 18.485 39.550 18.775 40.715 ;
        RECT 18.950 39.575 19.285 40.545 ;
        RECT 19.455 39.575 19.625 40.715 ;
        RECT 19.795 40.375 21.825 40.545 ;
        RECT 16.270 39.375 17.010 39.405 ;
        RECT 14.985 38.775 15.515 38.945 ;
        RECT 13.295 38.355 13.645 38.525 ;
        RECT 13.865 38.335 14.815 38.615 ;
        RECT 14.985 38.165 15.175 38.605 ;
        RECT 15.345 38.545 15.515 38.775 ;
        RECT 15.685 38.715 15.925 39.115 ;
        RECT 16.095 39.075 17.010 39.375 ;
        RECT 16.095 38.900 16.420 39.075 ;
        RECT 16.095 38.545 16.415 38.900 ;
        RECT 17.180 38.875 17.390 39.525 ;
        RECT 18.950 38.905 19.120 39.575 ;
        RECT 19.795 39.405 19.965 40.375 ;
        RECT 19.290 39.075 19.545 39.405 ;
        RECT 19.770 39.075 19.965 39.405 ;
        RECT 20.135 40.035 21.260 40.205 ;
        RECT 19.375 38.905 19.545 39.075 ;
        RECT 20.135 38.905 20.305 40.035 ;
        RECT 15.345 38.375 16.415 38.545 ;
        RECT 16.660 38.165 16.965 38.625 ;
        RECT 17.135 38.345 17.390 38.875 ;
        RECT 18.485 38.165 18.775 38.890 ;
        RECT 18.950 38.335 19.205 38.905 ;
        RECT 19.375 38.735 20.305 38.905 ;
        RECT 20.475 39.695 21.485 39.865 ;
        RECT 20.475 38.895 20.645 39.695 ;
        RECT 20.850 39.355 21.125 39.495 ;
        RECT 20.845 39.185 21.125 39.355 ;
        RECT 20.130 38.700 20.305 38.735 ;
        RECT 19.375 38.165 19.705 38.565 ;
        RECT 20.130 38.335 20.660 38.700 ;
        RECT 20.850 38.335 21.125 39.185 ;
        RECT 21.295 38.335 21.485 39.695 ;
        RECT 21.655 39.710 21.825 40.375 ;
        RECT 21.995 39.955 22.165 40.715 ;
        RECT 22.400 39.955 22.915 40.365 ;
        RECT 21.655 39.520 22.405 39.710 ;
        RECT 22.575 39.145 22.915 39.955 ;
        RECT 23.290 39.745 23.620 40.545 ;
        RECT 23.790 39.915 24.120 40.715 ;
        RECT 24.420 39.745 24.750 40.545 ;
        RECT 25.395 39.915 25.645 40.715 ;
        RECT 23.290 39.575 25.725 39.745 ;
        RECT 25.915 39.575 26.085 40.715 ;
        RECT 26.255 39.575 26.595 40.545 ;
        RECT 23.085 39.155 23.435 39.405 ;
        RECT 21.685 38.975 22.915 39.145 ;
        RECT 21.665 38.165 22.175 38.700 ;
        RECT 22.395 38.370 22.640 38.975 ;
        RECT 23.620 38.945 23.790 39.575 ;
        RECT 23.960 39.155 24.290 39.355 ;
        RECT 24.460 39.155 24.790 39.355 ;
        RECT 24.960 39.155 25.380 39.355 ;
        RECT 25.555 39.325 25.725 39.575 ;
        RECT 26.365 39.525 26.595 39.575 ;
        RECT 25.555 39.155 26.250 39.325 ;
        RECT 23.290 38.335 23.790 38.945 ;
        RECT 24.420 38.815 25.645 38.985 ;
        RECT 26.420 38.965 26.595 39.525 ;
        RECT 24.420 38.335 24.750 38.815 ;
        RECT 24.920 38.165 25.145 38.625 ;
        RECT 25.315 38.335 25.645 38.815 ;
        RECT 25.835 38.165 26.085 38.965 ;
        RECT 26.255 38.335 26.595 38.965 ;
        RECT 26.770 39.575 27.105 40.545 ;
        RECT 27.275 39.575 27.445 40.715 ;
        RECT 27.615 40.375 29.645 40.545 ;
        RECT 26.770 38.905 26.940 39.575 ;
        RECT 27.615 39.405 27.785 40.375 ;
        RECT 27.110 39.075 27.365 39.405 ;
        RECT 27.590 39.075 27.785 39.405 ;
        RECT 27.955 40.035 29.080 40.205 ;
        RECT 27.195 38.905 27.365 39.075 ;
        RECT 27.955 38.905 28.125 40.035 ;
        RECT 26.770 38.335 27.025 38.905 ;
        RECT 27.195 38.735 28.125 38.905 ;
        RECT 28.295 39.695 29.305 39.865 ;
        RECT 28.295 38.895 28.465 39.695 ;
        RECT 28.670 39.015 28.945 39.495 ;
        RECT 28.665 38.845 28.945 39.015 ;
        RECT 27.950 38.700 28.125 38.735 ;
        RECT 27.195 38.165 27.525 38.565 ;
        RECT 27.950 38.335 28.480 38.700 ;
        RECT 28.670 38.335 28.945 38.845 ;
        RECT 29.115 38.335 29.305 39.695 ;
        RECT 29.475 39.710 29.645 40.375 ;
        RECT 29.815 39.955 29.985 40.715 ;
        RECT 30.220 39.955 30.735 40.365 ;
        RECT 29.475 39.520 30.225 39.710 ;
        RECT 30.395 39.145 30.735 39.955 ;
        RECT 30.905 39.625 33.495 40.715 ;
        RECT 29.505 38.975 30.735 39.145 ;
        RECT 29.485 38.165 29.995 38.700 ;
        RECT 30.215 38.370 30.460 38.975 ;
        RECT 30.905 38.935 32.115 39.455 ;
        RECT 32.285 39.105 33.495 39.625 ;
        RECT 33.670 39.575 34.005 40.545 ;
        RECT 34.175 39.575 34.345 40.715 ;
        RECT 34.515 40.375 36.545 40.545 ;
        RECT 30.905 38.165 33.495 38.935 ;
        RECT 33.670 38.905 33.840 39.575 ;
        RECT 34.515 39.405 34.685 40.375 ;
        RECT 34.010 39.075 34.265 39.405 ;
        RECT 34.490 39.075 34.685 39.405 ;
        RECT 34.855 40.035 35.980 40.205 ;
        RECT 34.095 38.905 34.265 39.075 ;
        RECT 34.855 38.905 35.025 40.035 ;
        RECT 33.670 38.335 33.925 38.905 ;
        RECT 34.095 38.735 35.025 38.905 ;
        RECT 35.195 39.695 36.205 39.865 ;
        RECT 35.195 38.895 35.365 39.695 ;
        RECT 34.850 38.700 35.025 38.735 ;
        RECT 34.095 38.165 34.425 38.565 ;
        RECT 34.850 38.335 35.380 38.700 ;
        RECT 35.570 38.675 35.845 39.495 ;
        RECT 35.565 38.505 35.845 38.675 ;
        RECT 35.570 38.335 35.845 38.505 ;
        RECT 36.015 38.335 36.205 39.695 ;
        RECT 36.375 39.710 36.545 40.375 ;
        RECT 36.715 39.955 36.885 40.715 ;
        RECT 37.120 39.955 37.635 40.365 ;
        RECT 36.375 39.520 37.125 39.710 ;
        RECT 37.295 39.145 37.635 39.955 ;
        RECT 37.805 39.625 41.315 40.715 ;
        RECT 41.485 39.625 42.695 40.715 ;
        RECT 36.405 38.975 37.635 39.145 ;
        RECT 36.385 38.165 36.895 38.700 ;
        RECT 37.115 38.370 37.360 38.975 ;
        RECT 37.805 38.935 39.455 39.455 ;
        RECT 39.625 39.105 41.315 39.625 ;
        RECT 37.805 38.165 41.315 38.935 ;
        RECT 41.485 38.915 42.005 39.455 ;
        RECT 42.175 39.085 42.695 39.625 ;
        RECT 42.905 39.575 43.135 40.715 ;
        RECT 43.305 39.565 43.635 40.545 ;
        RECT 43.805 39.575 44.015 40.715 ;
        RECT 42.885 39.155 43.215 39.405 ;
        RECT 41.485 38.165 42.695 38.915 ;
        RECT 42.905 38.165 43.135 38.985 ;
        RECT 43.385 38.965 43.635 39.565 ;
        RECT 44.245 39.550 44.535 40.715 ;
        RECT 44.710 40.045 44.965 40.545 ;
        RECT 45.135 40.215 45.465 40.715 ;
        RECT 44.710 39.875 45.460 40.045 ;
        RECT 44.710 39.055 45.060 39.705 ;
        RECT 43.305 38.335 43.635 38.965 ;
        RECT 43.805 38.165 44.015 38.985 ;
        RECT 44.245 38.165 44.535 38.890 ;
        RECT 45.230 38.885 45.460 39.875 ;
        RECT 44.710 38.715 45.460 38.885 ;
        RECT 44.710 38.425 44.965 38.715 ;
        RECT 45.135 38.165 45.465 38.545 ;
        RECT 45.635 38.425 45.805 40.545 ;
        RECT 45.975 39.745 46.300 40.530 ;
        RECT 46.470 40.255 46.720 40.715 ;
        RECT 46.890 40.215 47.140 40.545 ;
        RECT 47.355 40.215 48.035 40.545 ;
        RECT 46.890 40.085 47.060 40.215 ;
        RECT 46.665 39.915 47.060 40.085 ;
        RECT 46.035 38.695 46.495 39.745 ;
        RECT 46.665 38.555 46.835 39.915 ;
        RECT 47.230 39.655 47.695 40.045 ;
        RECT 47.005 38.845 47.355 39.465 ;
        RECT 47.525 39.065 47.695 39.655 ;
        RECT 47.865 39.435 48.035 40.215 ;
        RECT 48.205 40.115 48.375 40.455 ;
        RECT 48.610 40.285 48.940 40.715 ;
        RECT 49.110 40.115 49.280 40.455 ;
        RECT 49.575 40.255 49.945 40.715 ;
        RECT 48.205 39.945 49.280 40.115 ;
        RECT 50.115 40.085 50.285 40.545 ;
        RECT 50.520 40.205 51.390 40.545 ;
        RECT 51.560 40.255 51.810 40.715 ;
        RECT 49.725 39.915 50.285 40.085 ;
        RECT 49.725 39.775 49.895 39.915 ;
        RECT 48.395 39.605 49.895 39.775 ;
        RECT 50.590 39.745 51.050 40.035 ;
        RECT 47.865 39.265 49.555 39.435 ;
        RECT 47.525 38.845 47.880 39.065 ;
        RECT 48.050 38.555 48.220 39.265 ;
        RECT 48.425 38.845 49.215 39.095 ;
        RECT 49.385 39.085 49.555 39.265 ;
        RECT 49.725 38.915 49.895 39.605 ;
        RECT 46.165 38.165 46.495 38.525 ;
        RECT 46.665 38.385 47.160 38.555 ;
        RECT 47.365 38.385 48.220 38.555 ;
        RECT 49.095 38.165 49.425 38.625 ;
        RECT 49.635 38.525 49.895 38.915 ;
        RECT 50.085 39.735 51.050 39.745 ;
        RECT 51.220 39.825 51.390 40.205 ;
        RECT 51.980 40.165 52.150 40.455 ;
        RECT 52.330 40.335 52.660 40.715 ;
        RECT 51.980 39.995 52.780 40.165 ;
        RECT 50.085 39.575 50.760 39.735 ;
        RECT 51.220 39.655 52.440 39.825 ;
        RECT 50.085 38.785 50.295 39.575 ;
        RECT 51.220 39.565 51.390 39.655 ;
        RECT 50.465 38.785 50.815 39.405 ;
        RECT 50.985 39.395 51.390 39.565 ;
        RECT 50.985 38.615 51.155 39.395 ;
        RECT 51.325 38.945 51.545 39.225 ;
        RECT 51.725 39.115 52.265 39.485 ;
        RECT 52.610 39.405 52.780 39.995 ;
        RECT 53.000 39.575 53.305 40.715 ;
        RECT 53.475 39.525 53.730 40.405 ;
        RECT 52.610 39.375 53.350 39.405 ;
        RECT 51.325 38.775 51.855 38.945 ;
        RECT 49.635 38.355 49.985 38.525 ;
        RECT 50.205 38.335 51.155 38.615 ;
        RECT 51.325 38.165 51.515 38.605 ;
        RECT 51.685 38.545 51.855 38.775 ;
        RECT 52.025 38.715 52.265 39.115 ;
        RECT 52.435 39.075 53.350 39.375 ;
        RECT 52.435 38.900 52.760 39.075 ;
        RECT 52.435 38.545 52.755 38.900 ;
        RECT 53.520 38.875 53.730 39.525 ;
        RECT 51.685 38.375 52.755 38.545 ;
        RECT 53.000 38.165 53.305 38.625 ;
        RECT 53.475 38.345 53.730 38.875 ;
        RECT 54.825 38.905 55.085 40.530 ;
        RECT 56.835 40.265 57.165 40.715 ;
        RECT 58.240 40.215 58.490 40.715 ;
        RECT 58.660 40.115 59.015 40.530 ;
        RECT 55.265 39.875 57.875 40.085 ;
        RECT 55.265 39.075 55.485 39.875 ;
        RECT 55.725 39.075 56.025 39.695 ;
        RECT 56.195 39.075 56.525 39.695 ;
        RECT 56.695 39.075 57.015 39.695 ;
        RECT 57.185 39.075 57.535 39.695 ;
        RECT 57.705 38.905 57.875 39.875 ;
        RECT 58.045 39.365 58.295 40.035 ;
        RECT 58.045 39.155 58.675 39.365 ;
        RECT 58.845 39.325 59.015 40.115 ;
        RECT 59.185 40.375 60.270 40.545 ;
        RECT 59.185 39.875 59.430 40.375 ;
        RECT 59.600 39.705 59.850 40.205 ;
        RECT 59.445 39.535 59.850 39.705 ;
        RECT 60.020 39.705 60.270 40.375 ;
        RECT 60.440 40.375 62.085 40.545 ;
        RECT 60.440 39.875 60.650 40.375 ;
        RECT 60.820 39.705 61.205 40.205 ;
        RECT 60.020 39.535 61.205 39.705 ;
        RECT 61.375 39.705 61.705 40.205 ;
        RECT 61.875 39.875 62.085 40.375 ;
        RECT 62.255 39.705 62.505 40.545 ;
        RECT 62.675 39.875 62.885 40.715 ;
        RECT 63.055 39.705 63.395 40.545 ;
        RECT 64.275 40.265 64.605 40.715 ;
        RECT 61.375 39.535 63.395 39.705 ;
        RECT 63.565 39.875 66.175 40.085 ;
        RECT 58.845 39.155 59.160 39.325 ;
        RECT 59.445 39.155 59.765 39.535 ;
        RECT 59.945 39.155 60.665 39.365 ;
        RECT 60.845 39.155 62.060 39.365 ;
        RECT 62.240 39.155 63.380 39.365 ;
        RECT 58.845 38.985 59.015 39.155 ;
        RECT 54.825 38.735 56.665 38.905 ;
        RECT 55.095 38.165 55.425 38.560 ;
        RECT 55.595 38.380 55.795 38.735 ;
        RECT 55.965 38.165 56.295 38.565 ;
        RECT 56.465 38.390 56.665 38.735 ;
        RECT 56.835 38.165 57.165 38.905 ;
        RECT 57.400 38.735 57.875 38.905 ;
        RECT 57.400 38.485 57.570 38.735 ;
        RECT 58.240 38.165 58.490 38.905 ;
        RECT 58.660 38.460 59.015 38.985 ;
        RECT 59.560 38.985 59.765 39.155 ;
        RECT 59.185 38.165 59.390 38.975 ;
        RECT 59.560 38.805 62.965 38.985 ;
        RECT 59.560 38.335 59.890 38.805 ;
        RECT 60.060 38.165 60.230 38.635 ;
        RECT 60.400 38.335 60.730 38.805 ;
        RECT 60.900 38.165 61.625 38.635 ;
        RECT 61.795 38.335 62.125 38.805 ;
        RECT 62.295 38.165 62.465 38.635 ;
        RECT 62.635 38.335 62.965 38.805 ;
        RECT 63.135 38.165 63.395 38.985 ;
        RECT 63.565 38.905 63.735 39.875 ;
        RECT 63.905 39.075 64.255 39.695 ;
        RECT 64.425 39.075 64.745 39.695 ;
        RECT 64.915 39.075 65.245 39.695 ;
        RECT 65.415 39.075 65.715 39.695 ;
        RECT 65.955 39.075 66.175 39.875 ;
        RECT 66.355 38.905 66.615 40.530 ;
        RECT 66.785 39.625 69.375 40.715 ;
        RECT 63.565 38.735 64.040 38.905 ;
        RECT 63.870 38.485 64.040 38.735 ;
        RECT 64.275 38.165 64.605 38.905 ;
        RECT 64.775 38.735 66.615 38.905 ;
        RECT 66.785 38.935 67.995 39.455 ;
        RECT 68.165 39.105 69.375 39.625 ;
        RECT 70.005 39.550 70.295 40.715 ;
        RECT 70.465 39.625 72.135 40.715 ;
        RECT 70.465 38.935 71.215 39.455 ;
        RECT 71.385 39.105 72.135 39.625 ;
        RECT 72.805 39.575 73.035 40.715 ;
        RECT 73.205 39.565 73.535 40.545 ;
        RECT 73.705 39.575 73.915 40.715 ;
        RECT 74.145 39.625 76.735 40.715 ;
        RECT 72.785 39.155 73.115 39.405 ;
        RECT 64.775 38.390 64.975 38.735 ;
        RECT 65.145 38.165 65.475 38.565 ;
        RECT 65.645 38.380 65.845 38.735 ;
        RECT 66.015 38.165 66.345 38.560 ;
        RECT 66.785 38.165 69.375 38.935 ;
        RECT 70.005 38.165 70.295 38.890 ;
        RECT 70.465 38.165 72.135 38.935 ;
        RECT 72.805 38.165 73.035 38.985 ;
        RECT 73.285 38.965 73.535 39.565 ;
        RECT 73.205 38.335 73.535 38.965 ;
        RECT 73.705 38.165 73.915 38.985 ;
        RECT 74.145 38.935 75.355 39.455 ;
        RECT 75.525 39.105 76.735 39.625 ;
        RECT 77.410 39.575 77.705 40.715 ;
        RECT 77.965 39.745 78.295 40.545 ;
        RECT 78.465 39.915 78.635 40.715 ;
        RECT 78.805 39.745 79.135 40.545 ;
        RECT 79.305 39.915 79.475 40.715 ;
        RECT 79.645 39.765 79.975 40.545 ;
        RECT 80.145 40.255 80.315 40.715 ;
        RECT 79.645 39.745 80.415 39.765 ;
        RECT 77.965 39.575 80.415 39.745 ;
        RECT 77.385 39.155 79.895 39.405 ;
        RECT 80.065 38.985 80.415 39.575 ;
        RECT 74.145 38.165 76.735 38.935 ;
        RECT 78.045 38.805 80.415 38.985 ;
        RECT 80.585 39.640 80.855 40.545 ;
        RECT 81.025 39.955 81.355 40.715 ;
        RECT 81.535 39.785 81.705 40.545 ;
        RECT 80.585 38.840 80.755 39.640 ;
        RECT 81.040 39.615 81.705 39.785 ;
        RECT 82.055 39.785 82.225 40.545 ;
        RECT 82.405 39.955 82.735 40.715 ;
        RECT 82.055 39.615 82.720 39.785 ;
        RECT 82.905 39.640 83.175 40.545 ;
        RECT 81.040 39.470 81.210 39.615 ;
        RECT 80.925 39.140 81.210 39.470 ;
        RECT 82.550 39.470 82.720 39.615 ;
        RECT 81.040 38.885 81.210 39.140 ;
        RECT 81.445 39.065 81.775 39.435 ;
        RECT 81.985 39.065 82.315 39.435 ;
        RECT 82.550 39.140 82.835 39.470 ;
        RECT 82.550 38.885 82.720 39.140 ;
        RECT 77.410 38.165 77.675 38.625 ;
        RECT 78.045 38.335 78.215 38.805 ;
        RECT 78.465 38.165 78.635 38.625 ;
        RECT 78.885 38.335 79.055 38.805 ;
        RECT 79.305 38.165 79.475 38.625 ;
        RECT 79.725 38.335 79.895 38.805 ;
        RECT 80.065 38.165 80.315 38.630 ;
        RECT 80.585 38.335 80.845 38.840 ;
        RECT 81.040 38.715 81.705 38.885 ;
        RECT 81.025 38.165 81.355 38.545 ;
        RECT 81.535 38.335 81.705 38.715 ;
        RECT 82.055 38.715 82.720 38.885 ;
        RECT 83.005 38.840 83.175 39.640 ;
        RECT 83.435 39.785 83.605 40.545 ;
        RECT 83.785 39.955 84.115 40.715 ;
        RECT 83.435 39.615 84.100 39.785 ;
        RECT 84.285 39.640 84.555 40.545 ;
        RECT 83.930 39.470 84.100 39.615 ;
        RECT 83.365 39.065 83.695 39.435 ;
        RECT 83.930 39.140 84.215 39.470 ;
        RECT 83.930 38.885 84.100 39.140 ;
        RECT 82.055 38.335 82.225 38.715 ;
        RECT 82.405 38.165 82.735 38.545 ;
        RECT 82.915 38.335 83.175 38.840 ;
        RECT 83.435 38.715 84.100 38.885 ;
        RECT 84.385 38.840 84.555 39.640 ;
        RECT 83.435 38.335 83.605 38.715 ;
        RECT 83.785 38.165 84.115 38.545 ;
        RECT 84.295 38.335 84.555 38.840 ;
        RECT 84.725 39.575 85.110 40.545 ;
        RECT 85.280 40.255 85.605 40.715 ;
        RECT 86.125 40.085 86.405 40.545 ;
        RECT 85.280 39.865 86.405 40.085 ;
        RECT 84.725 38.905 85.005 39.575 ;
        RECT 85.280 39.405 85.730 39.865 ;
        RECT 86.595 39.695 86.995 40.545 ;
        RECT 87.395 40.255 87.665 40.715 ;
        RECT 87.835 40.085 88.120 40.545 ;
        RECT 85.175 39.075 85.730 39.405 ;
        RECT 85.900 39.135 86.995 39.695 ;
        RECT 85.280 38.965 85.730 39.075 ;
        RECT 84.725 38.335 85.110 38.905 ;
        RECT 85.280 38.795 86.405 38.965 ;
        RECT 85.280 38.165 85.605 38.625 ;
        RECT 86.125 38.335 86.405 38.795 ;
        RECT 86.595 38.335 86.995 39.135 ;
        RECT 87.165 39.865 88.120 40.085 ;
        RECT 87.165 38.965 87.375 39.865 ;
        RECT 87.545 39.135 88.235 39.695 ;
        RECT 88.405 39.575 88.790 40.545 ;
        RECT 88.960 40.255 89.285 40.715 ;
        RECT 89.805 40.085 90.085 40.545 ;
        RECT 88.960 39.865 90.085 40.085 ;
        RECT 87.165 38.795 88.120 38.965 ;
        RECT 87.395 38.165 87.665 38.625 ;
        RECT 87.835 38.335 88.120 38.795 ;
        RECT 88.405 38.905 88.685 39.575 ;
        RECT 88.960 39.405 89.410 39.865 ;
        RECT 90.275 39.695 90.675 40.545 ;
        RECT 91.075 40.255 91.345 40.715 ;
        RECT 91.515 40.085 91.800 40.545 ;
        RECT 88.855 39.075 89.410 39.405 ;
        RECT 89.580 39.135 90.675 39.695 ;
        RECT 88.960 38.965 89.410 39.075 ;
        RECT 88.405 38.335 88.790 38.905 ;
        RECT 88.960 38.795 90.085 38.965 ;
        RECT 88.960 38.165 89.285 38.625 ;
        RECT 89.805 38.335 90.085 38.795 ;
        RECT 90.275 38.335 90.675 39.135 ;
        RECT 90.845 39.865 91.800 40.085 ;
        RECT 90.845 38.965 91.055 39.865 ;
        RECT 91.225 39.135 91.915 39.695 ;
        RECT 92.085 39.575 92.470 40.545 ;
        RECT 92.640 40.255 92.965 40.715 ;
        RECT 93.485 40.085 93.765 40.545 ;
        RECT 92.640 39.865 93.765 40.085 ;
        RECT 90.845 38.795 91.800 38.965 ;
        RECT 91.075 38.165 91.345 38.625 ;
        RECT 91.515 38.335 91.800 38.795 ;
        RECT 92.085 38.905 92.365 39.575 ;
        RECT 92.640 39.405 93.090 39.865 ;
        RECT 93.955 39.695 94.355 40.545 ;
        RECT 94.755 40.255 95.025 40.715 ;
        RECT 95.195 40.085 95.480 40.545 ;
        RECT 92.535 39.075 93.090 39.405 ;
        RECT 93.260 39.135 94.355 39.695 ;
        RECT 92.640 38.965 93.090 39.075 ;
        RECT 92.085 38.335 92.470 38.905 ;
        RECT 92.640 38.795 93.765 38.965 ;
        RECT 92.640 38.165 92.965 38.625 ;
        RECT 93.485 38.335 93.765 38.795 ;
        RECT 93.955 38.335 94.355 39.135 ;
        RECT 94.525 39.865 95.480 40.085 ;
        RECT 94.525 38.965 94.735 39.865 ;
        RECT 94.905 39.135 95.595 39.695 ;
        RECT 95.765 39.550 96.055 40.715 ;
        RECT 96.225 39.625 97.895 40.715 ;
        RECT 94.525 38.795 95.480 38.965 ;
        RECT 96.225 38.935 96.975 39.455 ;
        RECT 97.145 39.105 97.895 39.625 ;
        RECT 98.525 39.955 99.040 40.365 ;
        RECT 99.275 39.955 99.445 40.715 ;
        RECT 99.615 40.375 101.645 40.545 ;
        RECT 98.525 39.145 98.865 39.955 ;
        RECT 99.615 39.710 99.785 40.375 ;
        RECT 100.180 40.035 101.305 40.205 ;
        RECT 99.035 39.520 99.785 39.710 ;
        RECT 99.955 39.695 100.965 39.865 ;
        RECT 98.525 38.975 99.755 39.145 ;
        RECT 94.755 38.165 95.025 38.625 ;
        RECT 95.195 38.335 95.480 38.795 ;
        RECT 95.765 38.165 96.055 38.890 ;
        RECT 96.225 38.165 97.895 38.935 ;
        RECT 98.800 38.370 99.045 38.975 ;
        RECT 99.265 38.165 99.775 38.700 ;
        RECT 99.955 38.335 100.145 39.695 ;
        RECT 100.315 39.015 100.590 39.495 ;
        RECT 100.315 38.845 100.595 39.015 ;
        RECT 100.795 38.895 100.965 39.695 ;
        RECT 101.135 38.905 101.305 40.035 ;
        RECT 101.475 39.405 101.645 40.375 ;
        RECT 101.815 39.575 101.985 40.715 ;
        RECT 102.155 39.575 102.490 40.545 ;
        RECT 101.475 39.075 101.670 39.405 ;
        RECT 101.895 39.075 102.150 39.405 ;
        RECT 101.895 38.905 102.065 39.075 ;
        RECT 102.320 38.905 102.490 39.575 ;
        RECT 100.315 38.335 100.590 38.845 ;
        RECT 101.135 38.735 102.065 38.905 ;
        RECT 101.135 38.700 101.310 38.735 ;
        RECT 100.780 38.335 101.310 38.700 ;
        RECT 101.735 38.165 102.065 38.565 ;
        RECT 102.235 38.335 102.490 38.905 ;
        RECT 102.665 39.575 103.050 40.545 ;
        RECT 103.220 40.255 103.545 40.715 ;
        RECT 104.065 40.085 104.345 40.545 ;
        RECT 103.220 39.865 104.345 40.085 ;
        RECT 102.665 38.905 102.945 39.575 ;
        RECT 103.220 39.405 103.670 39.865 ;
        RECT 104.535 39.695 104.935 40.545 ;
        RECT 105.335 40.255 105.605 40.715 ;
        RECT 105.775 40.085 106.060 40.545 ;
        RECT 103.115 39.075 103.670 39.405 ;
        RECT 103.840 39.135 104.935 39.695 ;
        RECT 103.220 38.965 103.670 39.075 ;
        RECT 102.665 38.335 103.050 38.905 ;
        RECT 103.220 38.795 104.345 38.965 ;
        RECT 103.220 38.165 103.545 38.625 ;
        RECT 104.065 38.335 104.345 38.795 ;
        RECT 104.535 38.335 104.935 39.135 ;
        RECT 105.105 39.865 106.060 40.085 ;
        RECT 106.460 40.085 106.745 40.545 ;
        RECT 106.915 40.255 107.185 40.715 ;
        RECT 106.460 39.865 107.415 40.085 ;
        RECT 105.105 38.965 105.315 39.865 ;
        RECT 105.485 39.135 106.175 39.695 ;
        RECT 106.345 39.135 107.035 39.695 ;
        RECT 107.205 38.965 107.415 39.865 ;
        RECT 105.105 38.795 106.060 38.965 ;
        RECT 105.335 38.165 105.605 38.625 ;
        RECT 105.775 38.335 106.060 38.795 ;
        RECT 106.460 38.795 107.415 38.965 ;
        RECT 107.585 39.695 107.985 40.545 ;
        RECT 108.175 40.085 108.455 40.545 ;
        RECT 108.975 40.255 109.300 40.715 ;
        RECT 108.175 39.865 109.300 40.085 ;
        RECT 107.585 39.135 108.680 39.695 ;
        RECT 108.850 39.405 109.300 39.865 ;
        RECT 109.470 39.575 109.855 40.545 ;
        RECT 106.460 38.335 106.745 38.795 ;
        RECT 106.915 38.165 107.185 38.625 ;
        RECT 107.585 38.335 107.985 39.135 ;
        RECT 108.850 39.075 109.405 39.405 ;
        RECT 108.850 38.965 109.300 39.075 ;
        RECT 108.175 38.795 109.300 38.965 ;
        RECT 109.575 38.905 109.855 39.575 ;
        RECT 108.175 38.335 108.455 38.795 ;
        RECT 108.975 38.165 109.300 38.625 ;
        RECT 109.470 38.335 109.855 38.905 ;
        RECT 110.025 39.640 110.295 40.545 ;
        RECT 110.465 39.955 110.795 40.715 ;
        RECT 110.975 39.785 111.145 40.545 ;
        RECT 111.405 40.280 116.750 40.715 ;
        RECT 110.025 38.840 110.195 39.640 ;
        RECT 110.480 39.615 111.145 39.785 ;
        RECT 110.480 39.470 110.650 39.615 ;
        RECT 110.365 39.140 110.650 39.470 ;
        RECT 110.480 38.885 110.650 39.140 ;
        RECT 110.885 39.065 111.215 39.435 ;
        RECT 110.025 38.335 110.285 38.840 ;
        RECT 110.480 38.715 111.145 38.885 ;
        RECT 110.465 38.165 110.795 38.545 ;
        RECT 110.975 38.335 111.145 38.715 ;
        RECT 112.990 38.710 113.330 39.540 ;
        RECT 114.810 39.030 115.160 40.280 ;
        RECT 117.385 39.625 118.595 40.715 ;
        RECT 117.385 39.085 117.905 39.625 ;
        RECT 118.075 38.915 118.595 39.455 ;
        RECT 111.405 38.165 116.750 38.710 ;
        RECT 117.385 38.165 118.595 38.915 ;
        RECT 5.520 37.995 118.680 38.165 ;
        RECT 5.605 37.245 6.815 37.995 ;
        RECT 6.985 37.450 12.330 37.995 ;
        RECT 12.505 37.450 17.850 37.995 ;
        RECT 5.605 36.705 6.125 37.245 ;
        RECT 6.295 36.535 6.815 37.075 ;
        RECT 8.570 36.620 8.910 37.450 ;
        RECT 5.605 35.445 6.815 36.535 ;
        RECT 10.390 35.880 10.740 37.130 ;
        RECT 14.090 36.620 14.430 37.450 ;
        RECT 18.025 37.245 19.235 37.995 ;
        RECT 19.405 37.255 19.790 37.825 ;
        RECT 19.960 37.535 20.285 37.995 ;
        RECT 20.805 37.365 21.085 37.825 ;
        RECT 15.910 35.880 16.260 37.130 ;
        RECT 18.025 36.705 18.545 37.245 ;
        RECT 18.715 36.535 19.235 37.075 ;
        RECT 6.985 35.445 12.330 35.880 ;
        RECT 12.505 35.445 17.850 35.880 ;
        RECT 18.025 35.445 19.235 36.535 ;
        RECT 19.405 36.585 19.685 37.255 ;
        RECT 19.960 37.195 21.085 37.365 ;
        RECT 19.960 37.085 20.410 37.195 ;
        RECT 19.855 36.755 20.410 37.085 ;
        RECT 21.275 37.025 21.675 37.825 ;
        RECT 22.075 37.535 22.345 37.995 ;
        RECT 22.515 37.365 22.800 37.825 ;
        RECT 19.405 35.615 19.790 36.585 ;
        RECT 19.960 36.295 20.410 36.755 ;
        RECT 20.580 36.465 21.675 37.025 ;
        RECT 19.960 36.075 21.085 36.295 ;
        RECT 19.960 35.445 20.285 35.905 ;
        RECT 20.805 35.615 21.085 36.075 ;
        RECT 21.275 35.615 21.675 36.465 ;
        RECT 21.845 37.195 22.800 37.365 ;
        RECT 23.085 37.255 23.470 37.825 ;
        RECT 23.640 37.535 23.965 37.995 ;
        RECT 24.485 37.365 24.765 37.825 ;
        RECT 21.845 36.295 22.055 37.195 ;
        RECT 22.225 36.465 22.915 37.025 ;
        RECT 23.085 36.585 23.365 37.255 ;
        RECT 23.640 37.195 24.765 37.365 ;
        RECT 23.640 37.085 24.090 37.195 ;
        RECT 23.535 36.755 24.090 37.085 ;
        RECT 24.955 37.025 25.355 37.825 ;
        RECT 25.755 37.535 26.025 37.995 ;
        RECT 26.195 37.365 26.480 37.825 ;
        RECT 21.845 36.075 22.800 36.295 ;
        RECT 22.075 35.445 22.345 35.905 ;
        RECT 22.515 35.615 22.800 36.075 ;
        RECT 23.085 35.615 23.470 36.585 ;
        RECT 23.640 36.295 24.090 36.755 ;
        RECT 24.260 36.465 25.355 37.025 ;
        RECT 23.640 36.075 24.765 36.295 ;
        RECT 23.640 35.445 23.965 35.905 ;
        RECT 24.485 35.615 24.765 36.075 ;
        RECT 24.955 35.615 25.355 36.465 ;
        RECT 25.525 37.195 26.480 37.365 ;
        RECT 27.340 37.365 27.625 37.825 ;
        RECT 27.795 37.535 28.065 37.995 ;
        RECT 27.340 37.195 28.295 37.365 ;
        RECT 25.525 36.295 25.735 37.195 ;
        RECT 25.905 36.465 26.595 37.025 ;
        RECT 27.225 36.465 27.915 37.025 ;
        RECT 28.085 36.295 28.295 37.195 ;
        RECT 25.525 36.075 26.480 36.295 ;
        RECT 25.755 35.445 26.025 35.905 ;
        RECT 26.195 35.615 26.480 36.075 ;
        RECT 27.340 36.075 28.295 36.295 ;
        RECT 28.465 37.025 28.865 37.825 ;
        RECT 29.055 37.365 29.335 37.825 ;
        RECT 29.855 37.535 30.180 37.995 ;
        RECT 29.055 37.195 30.180 37.365 ;
        RECT 30.350 37.255 30.735 37.825 ;
        RECT 31.365 37.270 31.655 37.995 ;
        RECT 29.730 37.085 30.180 37.195 ;
        RECT 28.465 36.465 29.560 37.025 ;
        RECT 29.730 36.755 30.285 37.085 ;
        RECT 27.340 35.615 27.625 36.075 ;
        RECT 27.795 35.445 28.065 35.905 ;
        RECT 28.465 35.615 28.865 36.465 ;
        RECT 29.730 36.295 30.180 36.755 ;
        RECT 30.455 36.585 30.735 37.255 ;
        RECT 31.885 37.175 32.095 37.995 ;
        RECT 32.265 37.195 32.595 37.825 ;
        RECT 29.055 36.075 30.180 36.295 ;
        RECT 29.055 35.615 29.335 36.075 ;
        RECT 29.855 35.445 30.180 35.905 ;
        RECT 30.350 35.615 30.735 36.585 ;
        RECT 31.365 35.445 31.655 36.610 ;
        RECT 32.265 36.595 32.515 37.195 ;
        RECT 32.765 37.175 32.995 37.995 ;
        RECT 33.205 37.320 33.465 37.825 ;
        RECT 33.645 37.615 33.975 37.995 ;
        RECT 34.155 37.445 34.325 37.825 ;
        RECT 32.685 36.755 33.015 37.005 ;
        RECT 31.885 35.445 32.095 36.585 ;
        RECT 32.265 35.615 32.595 36.595 ;
        RECT 32.765 35.445 32.995 36.585 ;
        RECT 33.205 36.520 33.375 37.320 ;
        RECT 33.660 37.275 34.325 37.445 ;
        RECT 33.660 37.020 33.830 37.275 ;
        RECT 35.505 37.255 35.890 37.825 ;
        RECT 36.060 37.535 36.385 37.995 ;
        RECT 36.905 37.365 37.185 37.825 ;
        RECT 33.545 36.690 33.830 37.020 ;
        RECT 34.065 36.725 34.395 37.095 ;
        RECT 33.660 36.545 33.830 36.690 ;
        RECT 35.505 36.585 35.785 37.255 ;
        RECT 36.060 37.195 37.185 37.365 ;
        RECT 36.060 37.085 36.510 37.195 ;
        RECT 35.955 36.755 36.510 37.085 ;
        RECT 37.375 37.025 37.775 37.825 ;
        RECT 38.175 37.535 38.445 37.995 ;
        RECT 38.615 37.365 38.900 37.825 ;
        RECT 39.185 37.450 44.530 37.995 ;
        RECT 33.205 35.615 33.475 36.520 ;
        RECT 33.660 36.375 34.325 36.545 ;
        RECT 33.645 35.445 33.975 36.205 ;
        RECT 34.155 35.615 34.325 36.375 ;
        RECT 35.505 35.615 35.890 36.585 ;
        RECT 36.060 36.295 36.510 36.755 ;
        RECT 36.680 36.465 37.775 37.025 ;
        RECT 36.060 36.075 37.185 36.295 ;
        RECT 36.060 35.445 36.385 35.905 ;
        RECT 36.905 35.615 37.185 36.075 ;
        RECT 37.375 35.615 37.775 36.465 ;
        RECT 37.945 37.195 38.900 37.365 ;
        RECT 37.945 36.295 38.155 37.195 ;
        RECT 38.325 36.465 39.015 37.025 ;
        RECT 40.770 36.620 41.110 37.450 ;
        RECT 44.710 37.255 44.965 37.825 ;
        RECT 45.135 37.595 45.465 37.995 ;
        RECT 45.890 37.460 46.420 37.825 ;
        RECT 46.610 37.655 46.885 37.825 ;
        RECT 46.605 37.485 46.885 37.655 ;
        RECT 45.890 37.425 46.065 37.460 ;
        RECT 45.135 37.255 46.065 37.425 ;
        RECT 37.945 36.075 38.900 36.295 ;
        RECT 38.175 35.445 38.445 35.905 ;
        RECT 38.615 35.615 38.900 36.075 ;
        RECT 42.590 35.880 42.940 37.130 ;
        RECT 44.710 36.585 44.880 37.255 ;
        RECT 45.135 37.085 45.305 37.255 ;
        RECT 45.050 36.755 45.305 37.085 ;
        RECT 45.530 36.755 45.725 37.085 ;
        RECT 39.185 35.445 44.530 35.880 ;
        RECT 44.710 35.615 45.045 36.585 ;
        RECT 45.215 35.445 45.385 36.585 ;
        RECT 45.555 35.785 45.725 36.755 ;
        RECT 45.895 36.125 46.065 37.255 ;
        RECT 46.235 36.465 46.405 37.265 ;
        RECT 46.610 36.665 46.885 37.485 ;
        RECT 47.055 36.465 47.245 37.825 ;
        RECT 47.425 37.460 47.935 37.995 ;
        RECT 48.155 37.185 48.400 37.790 ;
        RECT 48.845 37.450 54.190 37.995 ;
        RECT 47.445 37.015 48.675 37.185 ;
        RECT 46.235 36.295 47.245 36.465 ;
        RECT 47.415 36.450 48.165 36.640 ;
        RECT 45.895 35.955 47.020 36.125 ;
        RECT 47.415 35.785 47.585 36.450 ;
        RECT 48.335 36.205 48.675 37.015 ;
        RECT 50.430 36.620 50.770 37.450 ;
        RECT 54.365 37.225 56.955 37.995 ;
        RECT 57.125 37.270 57.415 37.995 ;
        RECT 57.585 37.495 57.845 37.825 ;
        RECT 58.155 37.615 58.485 37.995 ;
        RECT 58.665 37.655 60.145 37.825 ;
        RECT 45.555 35.615 47.585 35.785 ;
        RECT 47.755 35.445 47.925 36.205 ;
        RECT 48.160 35.795 48.675 36.205 ;
        RECT 52.250 35.880 52.600 37.130 ;
        RECT 54.365 36.705 55.575 37.225 ;
        RECT 55.745 36.535 56.955 37.055 ;
        RECT 57.585 36.795 57.755 37.495 ;
        RECT 58.665 37.325 59.065 37.655 ;
        RECT 58.105 37.135 58.315 37.315 ;
        RECT 58.105 36.965 58.725 37.135 ;
        RECT 58.895 36.845 59.065 37.325 ;
        RECT 59.255 37.155 59.805 37.485 ;
        RECT 57.585 36.625 58.715 36.795 ;
        RECT 58.895 36.675 59.465 36.845 ;
        RECT 48.845 35.445 54.190 35.880 ;
        RECT 54.365 35.445 56.955 36.535 ;
        RECT 57.125 35.445 57.415 36.610 ;
        RECT 57.585 35.945 57.755 36.625 ;
        RECT 58.545 36.505 58.715 36.625 ;
        RECT 57.925 36.125 58.275 36.455 ;
        RECT 58.545 36.335 59.125 36.505 ;
        RECT 59.295 36.165 59.465 36.675 ;
        RECT 58.725 35.995 59.465 36.165 ;
        RECT 59.635 36.165 59.805 37.155 ;
        RECT 59.975 36.755 60.145 37.655 ;
        RECT 60.395 37.085 60.580 37.665 ;
        RECT 60.850 37.085 61.045 37.660 ;
        RECT 61.255 37.615 61.585 37.995 ;
        RECT 60.395 36.755 60.625 37.085 ;
        RECT 60.850 36.755 61.105 37.085 ;
        RECT 60.395 36.445 60.580 36.755 ;
        RECT 60.850 36.445 61.045 36.755 ;
        RECT 61.415 36.165 61.585 37.085 ;
        RECT 59.635 35.995 61.585 36.165 ;
        RECT 57.585 35.615 57.845 35.945 ;
        RECT 58.155 35.445 58.485 35.825 ;
        RECT 58.725 35.615 58.915 35.995 ;
        RECT 59.165 35.445 59.495 35.825 ;
        RECT 59.705 35.615 59.875 35.995 ;
        RECT 60.070 35.445 60.400 35.825 ;
        RECT 60.660 35.615 60.830 35.995 ;
        RECT 61.255 35.445 61.585 35.825 ;
        RECT 61.755 35.615 62.015 37.825 ;
        RECT 62.185 37.450 67.530 37.995 ;
        RECT 67.705 37.450 73.050 37.995 ;
        RECT 63.770 36.620 64.110 37.450 ;
        RECT 65.590 35.880 65.940 37.130 ;
        RECT 69.290 36.620 69.630 37.450 ;
        RECT 73.690 37.445 73.945 37.735 ;
        RECT 74.115 37.615 74.445 37.995 ;
        RECT 73.690 37.275 74.440 37.445 ;
        RECT 71.110 35.880 71.460 37.130 ;
        RECT 73.690 36.455 74.040 37.105 ;
        RECT 74.210 36.285 74.440 37.275 ;
        RECT 73.690 36.115 74.440 36.285 ;
        RECT 62.185 35.445 67.530 35.880 ;
        RECT 67.705 35.445 73.050 35.880 ;
        RECT 73.690 35.615 73.945 36.115 ;
        RECT 74.115 35.445 74.445 35.945 ;
        RECT 74.615 35.615 74.785 37.735 ;
        RECT 75.145 37.635 75.475 37.995 ;
        RECT 75.645 37.605 76.140 37.775 ;
        RECT 76.345 37.605 77.200 37.775 ;
        RECT 75.015 36.415 75.475 37.465 ;
        RECT 74.955 35.630 75.280 36.415 ;
        RECT 75.645 36.245 75.815 37.605 ;
        RECT 75.985 36.695 76.335 37.315 ;
        RECT 76.505 37.095 76.860 37.315 ;
        RECT 76.505 36.505 76.675 37.095 ;
        RECT 77.030 36.895 77.200 37.605 ;
        RECT 78.075 37.535 78.405 37.995 ;
        RECT 78.615 37.635 78.965 37.805 ;
        RECT 77.405 37.065 78.195 37.315 ;
        RECT 78.615 37.245 78.875 37.635 ;
        RECT 79.185 37.545 80.135 37.825 ;
        RECT 80.305 37.555 80.495 37.995 ;
        RECT 80.665 37.615 81.735 37.785 ;
        RECT 78.365 36.895 78.535 37.075 ;
        RECT 75.645 36.075 76.040 36.245 ;
        RECT 76.210 36.115 76.675 36.505 ;
        RECT 76.845 36.725 78.535 36.895 ;
        RECT 75.870 35.945 76.040 36.075 ;
        RECT 76.845 35.945 77.015 36.725 ;
        RECT 78.705 36.555 78.875 37.245 ;
        RECT 77.375 36.385 78.875 36.555 ;
        RECT 79.065 36.585 79.275 37.375 ;
        RECT 79.445 36.755 79.795 37.375 ;
        RECT 79.965 36.765 80.135 37.545 ;
        RECT 80.665 37.385 80.835 37.615 ;
        RECT 80.305 37.215 80.835 37.385 ;
        RECT 80.305 36.935 80.525 37.215 ;
        RECT 81.005 37.045 81.245 37.445 ;
        RECT 79.965 36.595 80.370 36.765 ;
        RECT 80.705 36.675 81.245 37.045 ;
        RECT 81.415 37.260 81.735 37.615 ;
        RECT 81.980 37.535 82.285 37.995 ;
        RECT 82.455 37.285 82.710 37.815 ;
        RECT 81.415 37.085 81.740 37.260 ;
        RECT 81.415 36.785 82.330 37.085 ;
        RECT 81.590 36.755 82.330 36.785 ;
        RECT 79.065 36.425 79.740 36.585 ;
        RECT 80.200 36.505 80.370 36.595 ;
        RECT 79.065 36.415 80.030 36.425 ;
        RECT 78.705 36.245 78.875 36.385 ;
        RECT 75.450 35.445 75.700 35.905 ;
        RECT 75.870 35.615 76.120 35.945 ;
        RECT 76.335 35.615 77.015 35.945 ;
        RECT 77.185 36.045 78.260 36.215 ;
        RECT 78.705 36.075 79.265 36.245 ;
        RECT 79.570 36.125 80.030 36.415 ;
        RECT 80.200 36.335 81.420 36.505 ;
        RECT 77.185 35.705 77.355 36.045 ;
        RECT 77.590 35.445 77.920 35.875 ;
        RECT 78.090 35.705 78.260 36.045 ;
        RECT 78.555 35.445 78.925 35.905 ;
        RECT 79.095 35.615 79.265 36.075 ;
        RECT 80.200 35.955 80.370 36.335 ;
        RECT 81.590 36.165 81.760 36.755 ;
        RECT 82.500 36.635 82.710 37.285 ;
        RECT 82.885 37.270 83.175 37.995 ;
        RECT 83.405 37.175 83.615 37.995 ;
        RECT 83.785 37.195 84.115 37.825 ;
        RECT 79.500 35.615 80.370 35.955 ;
        RECT 80.960 35.995 81.760 36.165 ;
        RECT 80.540 35.445 80.790 35.905 ;
        RECT 80.960 35.705 81.130 35.995 ;
        RECT 81.310 35.445 81.640 35.825 ;
        RECT 81.980 35.445 82.285 36.585 ;
        RECT 82.455 35.755 82.710 36.635 ;
        RECT 82.885 35.445 83.175 36.610 ;
        RECT 83.785 36.595 84.035 37.195 ;
        RECT 84.285 37.175 84.515 37.995 ;
        RECT 85.460 37.185 85.705 37.790 ;
        RECT 85.925 37.460 86.435 37.995 ;
        RECT 85.185 37.015 86.415 37.185 ;
        RECT 84.205 36.755 84.535 37.005 ;
        RECT 83.405 35.445 83.615 36.585 ;
        RECT 83.785 35.615 84.115 36.595 ;
        RECT 84.285 35.445 84.515 36.585 ;
        RECT 85.185 36.205 85.525 37.015 ;
        RECT 85.695 36.450 86.445 36.640 ;
        RECT 85.185 35.795 85.700 36.205 ;
        RECT 85.935 35.445 86.105 36.205 ;
        RECT 86.275 35.785 86.445 36.450 ;
        RECT 86.615 36.465 86.805 37.825 ;
        RECT 86.975 37.655 87.250 37.825 ;
        RECT 86.975 37.485 87.255 37.655 ;
        RECT 86.975 36.665 87.250 37.485 ;
        RECT 87.440 37.460 87.970 37.825 ;
        RECT 88.395 37.595 88.725 37.995 ;
        RECT 87.795 37.425 87.970 37.460 ;
        RECT 87.455 36.465 87.625 37.265 ;
        RECT 86.615 36.295 87.625 36.465 ;
        RECT 87.795 37.255 88.725 37.425 ;
        RECT 88.895 37.255 89.150 37.825 ;
        RECT 87.795 36.125 87.965 37.255 ;
        RECT 88.555 37.085 88.725 37.255 ;
        RECT 86.840 35.955 87.965 36.125 ;
        RECT 88.135 36.755 88.330 37.085 ;
        RECT 88.555 36.755 88.810 37.085 ;
        RECT 88.135 35.785 88.305 36.755 ;
        RECT 88.980 36.585 89.150 37.255 ;
        RECT 86.275 35.615 88.305 35.785 ;
        RECT 88.475 35.445 88.645 36.585 ;
        RECT 88.815 35.615 89.150 36.585 ;
        RECT 89.330 37.255 89.585 37.825 ;
        RECT 89.755 37.595 90.085 37.995 ;
        RECT 90.510 37.460 91.040 37.825 ;
        RECT 91.230 37.655 91.505 37.825 ;
        RECT 91.225 37.485 91.505 37.655 ;
        RECT 90.510 37.425 90.685 37.460 ;
        RECT 89.755 37.255 90.685 37.425 ;
        RECT 89.330 36.585 89.500 37.255 ;
        RECT 89.755 37.085 89.925 37.255 ;
        RECT 89.670 36.755 89.925 37.085 ;
        RECT 90.150 36.755 90.345 37.085 ;
        RECT 89.330 35.615 89.665 36.585 ;
        RECT 89.835 35.445 90.005 36.585 ;
        RECT 90.175 35.785 90.345 36.755 ;
        RECT 90.515 36.125 90.685 37.255 ;
        RECT 90.855 36.465 91.025 37.265 ;
        RECT 91.230 36.665 91.505 37.485 ;
        RECT 91.675 36.465 91.865 37.825 ;
        RECT 92.045 37.460 92.555 37.995 ;
        RECT 92.775 37.185 93.020 37.790 ;
        RECT 92.065 37.015 93.295 37.185 ;
        RECT 93.525 37.175 93.735 37.995 ;
        RECT 93.905 37.195 94.235 37.825 ;
        RECT 90.855 36.295 91.865 36.465 ;
        RECT 92.035 36.450 92.785 36.640 ;
        RECT 90.515 35.955 91.640 36.125 ;
        RECT 92.035 35.785 92.205 36.450 ;
        RECT 92.955 36.205 93.295 37.015 ;
        RECT 93.905 36.595 94.155 37.195 ;
        RECT 94.405 37.175 94.635 37.995 ;
        RECT 94.845 37.225 97.435 37.995 ;
        RECT 98.070 37.445 98.325 37.735 ;
        RECT 98.495 37.615 98.825 37.995 ;
        RECT 98.070 37.275 98.820 37.445 ;
        RECT 94.325 36.755 94.655 37.005 ;
        RECT 94.845 36.705 96.055 37.225 ;
        RECT 90.175 35.615 92.205 35.785 ;
        RECT 92.375 35.445 92.545 36.205 ;
        RECT 92.780 35.795 93.295 36.205 ;
        RECT 93.525 35.445 93.735 36.585 ;
        RECT 93.905 35.615 94.235 36.595 ;
        RECT 94.405 35.445 94.635 36.585 ;
        RECT 96.225 36.535 97.435 37.055 ;
        RECT 94.845 35.445 97.435 36.535 ;
        RECT 98.070 36.455 98.420 37.105 ;
        RECT 98.590 36.285 98.820 37.275 ;
        RECT 98.070 36.115 98.820 36.285 ;
        RECT 98.070 35.615 98.325 36.115 ;
        RECT 98.495 35.445 98.825 35.945 ;
        RECT 98.995 35.615 99.165 37.735 ;
        RECT 99.525 37.635 99.855 37.995 ;
        RECT 100.025 37.605 100.520 37.775 ;
        RECT 100.725 37.605 101.580 37.775 ;
        RECT 99.395 36.415 99.855 37.465 ;
        RECT 99.335 35.630 99.660 36.415 ;
        RECT 100.025 36.245 100.195 37.605 ;
        RECT 100.365 36.695 100.715 37.315 ;
        RECT 100.885 37.095 101.240 37.315 ;
        RECT 100.885 36.505 101.055 37.095 ;
        RECT 101.410 36.895 101.580 37.605 ;
        RECT 102.455 37.535 102.785 37.995 ;
        RECT 102.995 37.635 103.345 37.805 ;
        RECT 101.785 37.065 102.575 37.315 ;
        RECT 102.995 37.245 103.255 37.635 ;
        RECT 103.565 37.545 104.515 37.825 ;
        RECT 104.685 37.555 104.875 37.995 ;
        RECT 105.045 37.615 106.115 37.785 ;
        RECT 102.745 36.895 102.915 37.075 ;
        RECT 100.025 36.075 100.420 36.245 ;
        RECT 100.590 36.115 101.055 36.505 ;
        RECT 101.225 36.725 102.915 36.895 ;
        RECT 100.250 35.945 100.420 36.075 ;
        RECT 101.225 35.945 101.395 36.725 ;
        RECT 103.085 36.555 103.255 37.245 ;
        RECT 101.755 36.385 103.255 36.555 ;
        RECT 103.445 36.585 103.655 37.375 ;
        RECT 103.825 36.755 104.175 37.375 ;
        RECT 104.345 36.765 104.515 37.545 ;
        RECT 105.045 37.385 105.215 37.615 ;
        RECT 104.685 37.215 105.215 37.385 ;
        RECT 104.685 36.935 104.905 37.215 ;
        RECT 105.385 37.045 105.625 37.445 ;
        RECT 104.345 36.595 104.750 36.765 ;
        RECT 105.085 36.675 105.625 37.045 ;
        RECT 105.795 37.260 106.115 37.615 ;
        RECT 106.360 37.535 106.665 37.995 ;
        RECT 106.835 37.285 107.090 37.815 ;
        RECT 105.795 37.085 106.120 37.260 ;
        RECT 105.795 36.785 106.710 37.085 ;
        RECT 105.970 36.755 106.710 36.785 ;
        RECT 103.445 36.425 104.120 36.585 ;
        RECT 104.580 36.505 104.750 36.595 ;
        RECT 103.445 36.415 104.410 36.425 ;
        RECT 103.085 36.245 103.255 36.385 ;
        RECT 99.830 35.445 100.080 35.905 ;
        RECT 100.250 35.615 100.500 35.945 ;
        RECT 100.715 35.615 101.395 35.945 ;
        RECT 101.565 36.045 102.640 36.215 ;
        RECT 103.085 36.075 103.645 36.245 ;
        RECT 103.950 36.125 104.410 36.415 ;
        RECT 104.580 36.335 105.800 36.505 ;
        RECT 101.565 35.705 101.735 36.045 ;
        RECT 101.970 35.445 102.300 35.875 ;
        RECT 102.470 35.705 102.640 36.045 ;
        RECT 102.935 35.445 103.305 35.905 ;
        RECT 103.475 35.615 103.645 36.075 ;
        RECT 104.580 35.955 104.750 36.335 ;
        RECT 105.970 36.165 106.140 36.755 ;
        RECT 106.880 36.635 107.090 37.285 ;
        RECT 107.265 37.245 108.475 37.995 ;
        RECT 108.645 37.270 108.935 37.995 ;
        RECT 109.105 37.450 114.450 37.995 ;
        RECT 107.265 36.705 107.785 37.245 ;
        RECT 103.880 35.615 104.750 35.955 ;
        RECT 105.340 35.995 106.140 36.165 ;
        RECT 104.920 35.445 105.170 35.905 ;
        RECT 105.340 35.705 105.510 35.995 ;
        RECT 105.690 35.445 106.020 35.825 ;
        RECT 106.360 35.445 106.665 36.585 ;
        RECT 106.835 35.755 107.090 36.635 ;
        RECT 107.955 36.535 108.475 37.075 ;
        RECT 110.690 36.620 111.030 37.450 ;
        RECT 114.625 37.225 117.215 37.995 ;
        RECT 117.385 37.245 118.595 37.995 ;
        RECT 107.265 35.445 108.475 36.535 ;
        RECT 108.645 35.445 108.935 36.610 ;
        RECT 112.510 35.880 112.860 37.130 ;
        RECT 114.625 36.705 115.835 37.225 ;
        RECT 116.005 36.535 117.215 37.055 ;
        RECT 109.105 35.445 114.450 35.880 ;
        RECT 114.625 35.445 117.215 36.535 ;
        RECT 117.385 36.535 117.905 37.075 ;
        RECT 118.075 36.705 118.595 37.245 ;
        RECT 117.385 35.445 118.595 36.535 ;
        RECT 5.520 35.275 118.680 35.445 ;
        RECT 5.605 34.185 6.815 35.275 ;
        RECT 6.985 34.840 12.330 35.275 ;
        RECT 12.505 34.840 17.850 35.275 ;
        RECT 5.605 33.475 6.125 34.015 ;
        RECT 6.295 33.645 6.815 34.185 ;
        RECT 5.605 32.725 6.815 33.475 ;
        RECT 8.570 33.270 8.910 34.100 ;
        RECT 10.390 33.590 10.740 34.840 ;
        RECT 14.090 33.270 14.430 34.100 ;
        RECT 15.910 33.590 16.260 34.840 ;
        RECT 18.485 34.110 18.775 35.275 ;
        RECT 18.945 34.200 19.215 35.105 ;
        RECT 19.385 34.515 19.715 35.275 ;
        RECT 19.895 34.345 20.065 35.105 ;
        RECT 6.985 32.725 12.330 33.270 ;
        RECT 12.505 32.725 17.850 33.270 ;
        RECT 18.485 32.725 18.775 33.450 ;
        RECT 18.945 33.400 19.115 34.200 ;
        RECT 19.400 34.175 20.065 34.345 ;
        RECT 20.325 34.185 21.995 35.275 ;
        RECT 22.740 34.645 23.025 35.105 ;
        RECT 23.195 34.815 23.465 35.275 ;
        RECT 22.740 34.425 23.695 34.645 ;
        RECT 19.400 34.030 19.570 34.175 ;
        RECT 19.285 33.700 19.570 34.030 ;
        RECT 19.400 33.445 19.570 33.700 ;
        RECT 19.805 33.625 20.135 33.995 ;
        RECT 20.325 33.495 21.075 34.015 ;
        RECT 21.245 33.665 21.995 34.185 ;
        RECT 22.625 33.695 23.315 34.255 ;
        RECT 23.485 33.525 23.695 34.425 ;
        RECT 18.945 32.895 19.205 33.400 ;
        RECT 19.400 33.275 20.065 33.445 ;
        RECT 19.385 32.725 19.715 33.105 ;
        RECT 19.895 32.895 20.065 33.275 ;
        RECT 20.325 32.725 21.995 33.495 ;
        RECT 22.740 33.355 23.695 33.525 ;
        RECT 23.865 34.255 24.265 35.105 ;
        RECT 24.455 34.645 24.735 35.105 ;
        RECT 25.255 34.815 25.580 35.275 ;
        RECT 24.455 34.425 25.580 34.645 ;
        RECT 23.865 33.695 24.960 34.255 ;
        RECT 25.130 33.965 25.580 34.425 ;
        RECT 25.750 34.135 26.135 35.105 ;
        RECT 26.310 34.605 26.565 35.105 ;
        RECT 26.735 34.775 27.065 35.275 ;
        RECT 26.310 34.435 27.060 34.605 ;
        RECT 22.740 32.895 23.025 33.355 ;
        RECT 23.195 32.725 23.465 33.185 ;
        RECT 23.865 32.895 24.265 33.695 ;
        RECT 25.130 33.635 25.685 33.965 ;
        RECT 25.130 33.525 25.580 33.635 ;
        RECT 24.455 33.355 25.580 33.525 ;
        RECT 25.855 33.465 26.135 34.135 ;
        RECT 26.310 33.615 26.660 34.265 ;
        RECT 24.455 32.895 24.735 33.355 ;
        RECT 25.255 32.725 25.580 33.185 ;
        RECT 25.750 32.895 26.135 33.465 ;
        RECT 26.830 33.445 27.060 34.435 ;
        RECT 26.310 33.275 27.060 33.445 ;
        RECT 26.310 32.985 26.565 33.275 ;
        RECT 26.735 32.725 27.065 33.105 ;
        RECT 27.235 32.985 27.405 35.105 ;
        RECT 27.575 34.305 27.900 35.090 ;
        RECT 28.070 34.815 28.320 35.275 ;
        RECT 28.490 34.775 28.740 35.105 ;
        RECT 28.955 34.775 29.635 35.105 ;
        RECT 28.490 34.645 28.660 34.775 ;
        RECT 28.265 34.475 28.660 34.645 ;
        RECT 27.635 33.255 28.095 34.305 ;
        RECT 28.265 33.115 28.435 34.475 ;
        RECT 28.830 34.215 29.295 34.605 ;
        RECT 28.605 33.405 28.955 34.025 ;
        RECT 29.125 33.625 29.295 34.215 ;
        RECT 29.465 33.995 29.635 34.775 ;
        RECT 29.805 34.675 29.975 35.015 ;
        RECT 30.210 34.845 30.540 35.275 ;
        RECT 30.710 34.675 30.880 35.015 ;
        RECT 31.175 34.815 31.545 35.275 ;
        RECT 29.805 34.505 30.880 34.675 ;
        RECT 31.715 34.645 31.885 35.105 ;
        RECT 32.120 34.765 32.990 35.105 ;
        RECT 33.160 34.815 33.410 35.275 ;
        RECT 31.325 34.475 31.885 34.645 ;
        RECT 31.325 34.335 31.495 34.475 ;
        RECT 29.995 34.165 31.495 34.335 ;
        RECT 32.190 34.305 32.650 34.595 ;
        RECT 29.465 33.825 31.155 33.995 ;
        RECT 29.125 33.405 29.480 33.625 ;
        RECT 29.650 33.115 29.820 33.825 ;
        RECT 30.025 33.405 30.815 33.655 ;
        RECT 30.985 33.645 31.155 33.825 ;
        RECT 31.325 33.475 31.495 34.165 ;
        RECT 27.765 32.725 28.095 33.085 ;
        RECT 28.265 32.945 28.760 33.115 ;
        RECT 28.965 32.945 29.820 33.115 ;
        RECT 30.695 32.725 31.025 33.185 ;
        RECT 31.235 33.085 31.495 33.475 ;
        RECT 31.685 34.295 32.650 34.305 ;
        RECT 32.820 34.385 32.990 34.765 ;
        RECT 33.580 34.725 33.750 35.015 ;
        RECT 33.930 34.895 34.260 35.275 ;
        RECT 33.580 34.555 34.380 34.725 ;
        RECT 31.685 34.135 32.360 34.295 ;
        RECT 32.820 34.215 34.040 34.385 ;
        RECT 31.685 33.345 31.895 34.135 ;
        RECT 32.820 34.125 32.990 34.215 ;
        RECT 32.065 33.345 32.415 33.965 ;
        RECT 32.585 33.955 32.990 34.125 ;
        RECT 32.585 33.175 32.755 33.955 ;
        RECT 32.925 33.505 33.145 33.785 ;
        RECT 33.325 33.675 33.865 34.045 ;
        RECT 34.210 33.965 34.380 34.555 ;
        RECT 34.600 34.135 34.905 35.275 ;
        RECT 35.075 34.085 35.330 34.965 ;
        RECT 35.505 34.840 40.850 35.275 ;
        RECT 34.210 33.935 34.950 33.965 ;
        RECT 32.925 33.335 33.455 33.505 ;
        RECT 31.235 32.915 31.585 33.085 ;
        RECT 31.805 32.895 32.755 33.175 ;
        RECT 32.925 32.725 33.115 33.165 ;
        RECT 33.285 33.105 33.455 33.335 ;
        RECT 33.625 33.275 33.865 33.675 ;
        RECT 34.035 33.635 34.950 33.935 ;
        RECT 34.035 33.460 34.360 33.635 ;
        RECT 34.035 33.105 34.355 33.460 ;
        RECT 35.120 33.435 35.330 34.085 ;
        RECT 33.285 32.935 34.355 33.105 ;
        RECT 34.600 32.725 34.905 33.185 ;
        RECT 35.075 32.905 35.330 33.435 ;
        RECT 37.090 33.270 37.430 34.100 ;
        RECT 38.910 33.590 39.260 34.840 ;
        RECT 41.025 34.185 42.695 35.275 ;
        RECT 41.025 33.495 41.775 34.015 ;
        RECT 41.945 33.665 42.695 34.185 ;
        RECT 42.865 34.200 43.135 35.105 ;
        RECT 43.305 34.515 43.635 35.275 ;
        RECT 43.815 34.345 43.985 35.105 ;
        RECT 35.505 32.725 40.850 33.270 ;
        RECT 41.025 32.725 42.695 33.495 ;
        RECT 42.865 33.400 43.035 34.200 ;
        RECT 43.320 34.175 43.985 34.345 ;
        RECT 43.320 34.030 43.490 34.175 ;
        RECT 44.245 34.110 44.535 35.275 ;
        RECT 45.205 34.135 45.435 35.275 ;
        RECT 45.605 34.125 45.935 35.105 ;
        RECT 46.105 34.135 46.315 35.275 ;
        RECT 46.545 34.840 51.890 35.275 ;
        RECT 52.065 34.840 57.410 35.275 ;
        RECT 57.585 34.840 62.930 35.275 ;
        RECT 43.205 33.700 43.490 34.030 ;
        RECT 43.320 33.445 43.490 33.700 ;
        RECT 43.725 33.625 44.055 33.995 ;
        RECT 45.185 33.715 45.515 33.965 ;
        RECT 42.865 32.895 43.125 33.400 ;
        RECT 43.320 33.275 43.985 33.445 ;
        RECT 43.305 32.725 43.635 33.105 ;
        RECT 43.815 32.895 43.985 33.275 ;
        RECT 44.245 32.725 44.535 33.450 ;
        RECT 45.205 32.725 45.435 33.545 ;
        RECT 45.685 33.525 45.935 34.125 ;
        RECT 45.605 32.895 45.935 33.525 ;
        RECT 46.105 32.725 46.315 33.545 ;
        RECT 48.130 33.270 48.470 34.100 ;
        RECT 49.950 33.590 50.300 34.840 ;
        RECT 53.650 33.270 53.990 34.100 ;
        RECT 55.470 33.590 55.820 34.840 ;
        RECT 59.170 33.270 59.510 34.100 ;
        RECT 60.990 33.590 61.340 34.840 ;
        RECT 63.105 34.185 65.695 35.275 ;
        RECT 63.105 33.495 64.315 34.015 ;
        RECT 64.485 33.665 65.695 34.185 ;
        RECT 65.865 34.135 66.250 35.105 ;
        RECT 66.420 34.815 66.745 35.275 ;
        RECT 67.265 34.645 67.545 35.105 ;
        RECT 66.420 34.425 67.545 34.645 ;
        RECT 46.545 32.725 51.890 33.270 ;
        RECT 52.065 32.725 57.410 33.270 ;
        RECT 57.585 32.725 62.930 33.270 ;
        RECT 63.105 32.725 65.695 33.495 ;
        RECT 65.865 33.465 66.145 34.135 ;
        RECT 66.420 33.965 66.870 34.425 ;
        RECT 67.735 34.255 68.135 35.105 ;
        RECT 68.535 34.815 68.805 35.275 ;
        RECT 68.975 34.645 69.260 35.105 ;
        RECT 66.315 33.635 66.870 33.965 ;
        RECT 67.040 33.695 68.135 34.255 ;
        RECT 66.420 33.525 66.870 33.635 ;
        RECT 65.865 32.895 66.250 33.465 ;
        RECT 66.420 33.355 67.545 33.525 ;
        RECT 66.420 32.725 66.745 33.185 ;
        RECT 67.265 32.895 67.545 33.355 ;
        RECT 67.735 32.895 68.135 33.695 ;
        RECT 68.305 34.425 69.260 34.645 ;
        RECT 68.305 33.525 68.515 34.425 ;
        RECT 68.685 33.695 69.375 34.255 ;
        RECT 70.005 34.110 70.295 35.275 ;
        RECT 70.465 34.185 71.675 35.275 ;
        RECT 68.305 33.355 69.260 33.525 ;
        RECT 70.465 33.475 70.985 34.015 ;
        RECT 71.155 33.645 71.675 34.185 ;
        RECT 71.935 34.345 72.105 35.105 ;
        RECT 72.285 34.515 72.615 35.275 ;
        RECT 71.935 34.175 72.600 34.345 ;
        RECT 72.785 34.200 73.055 35.105 ;
        RECT 72.430 34.030 72.600 34.175 ;
        RECT 71.865 33.625 72.195 33.995 ;
        RECT 72.430 33.700 72.715 34.030 ;
        RECT 68.535 32.725 68.805 33.185 ;
        RECT 68.975 32.895 69.260 33.355 ;
        RECT 70.005 32.725 70.295 33.450 ;
        RECT 70.465 32.725 71.675 33.475 ;
        RECT 72.430 33.445 72.600 33.700 ;
        RECT 71.935 33.275 72.600 33.445 ;
        RECT 72.885 33.400 73.055 34.200 ;
        RECT 71.935 32.895 72.105 33.275 ;
        RECT 72.285 32.725 72.615 33.105 ;
        RECT 72.795 32.895 73.055 33.400 ;
        RECT 73.230 34.135 73.565 35.105 ;
        RECT 73.735 34.135 73.905 35.275 ;
        RECT 74.075 34.935 76.105 35.105 ;
        RECT 73.230 33.465 73.400 34.135 ;
        RECT 74.075 33.965 74.245 34.935 ;
        RECT 73.570 33.635 73.825 33.965 ;
        RECT 74.050 33.635 74.245 33.965 ;
        RECT 74.415 34.595 75.540 34.765 ;
        RECT 73.655 33.465 73.825 33.635 ;
        RECT 74.415 33.465 74.585 34.595 ;
        RECT 73.230 32.895 73.485 33.465 ;
        RECT 73.655 33.295 74.585 33.465 ;
        RECT 74.755 34.255 75.765 34.425 ;
        RECT 74.755 33.455 74.925 34.255 ;
        RECT 74.410 33.260 74.585 33.295 ;
        RECT 73.655 32.725 73.985 33.125 ;
        RECT 74.410 32.895 74.940 33.260 ;
        RECT 75.130 33.235 75.405 34.055 ;
        RECT 75.125 33.065 75.405 33.235 ;
        RECT 75.130 32.895 75.405 33.065 ;
        RECT 75.575 32.895 75.765 34.255 ;
        RECT 75.935 34.270 76.105 34.935 ;
        RECT 76.275 34.515 76.445 35.275 ;
        RECT 76.680 34.515 77.195 34.925 ;
        RECT 75.935 34.080 76.685 34.270 ;
        RECT 76.855 33.705 77.195 34.515 ;
        RECT 77.375 34.465 77.670 35.275 ;
        RECT 77.850 33.965 78.095 35.105 ;
        RECT 78.270 34.465 78.530 35.275 ;
        RECT 79.130 35.270 85.405 35.275 ;
        RECT 78.710 33.965 78.960 35.100 ;
        RECT 79.130 34.475 79.390 35.270 ;
        RECT 79.560 34.375 79.820 35.100 ;
        RECT 79.990 34.545 80.250 35.270 ;
        RECT 80.420 34.375 80.680 35.100 ;
        RECT 80.850 34.545 81.110 35.270 ;
        RECT 81.280 34.375 81.540 35.100 ;
        RECT 81.710 34.545 81.970 35.270 ;
        RECT 82.140 34.375 82.400 35.100 ;
        RECT 82.570 34.545 82.815 35.270 ;
        RECT 82.985 34.375 83.245 35.100 ;
        RECT 83.430 34.545 83.675 35.270 ;
        RECT 83.845 34.375 84.105 35.100 ;
        RECT 84.290 34.545 84.535 35.270 ;
        RECT 84.705 34.375 84.965 35.100 ;
        RECT 85.150 34.545 85.405 35.270 ;
        RECT 79.560 34.360 84.965 34.375 ;
        RECT 85.575 34.360 85.865 35.100 ;
        RECT 86.035 34.530 86.305 35.275 ;
        RECT 86.570 34.605 86.825 35.105 ;
        RECT 86.995 34.775 87.325 35.275 ;
        RECT 86.570 34.435 87.320 34.605 ;
        RECT 79.560 34.135 86.305 34.360 ;
        RECT 75.965 33.535 77.195 33.705 ;
        RECT 75.945 32.725 76.455 33.260 ;
        RECT 76.675 32.930 76.920 33.535 ;
        RECT 77.365 33.405 77.680 33.965 ;
        RECT 77.850 33.715 84.970 33.965 ;
        RECT 77.365 32.725 77.670 33.235 ;
        RECT 77.850 32.905 78.100 33.715 ;
        RECT 78.270 32.725 78.530 33.250 ;
        RECT 78.710 32.905 78.960 33.715 ;
        RECT 85.140 33.545 86.305 34.135 ;
        RECT 86.570 33.615 86.920 34.265 ;
        RECT 79.560 33.375 86.305 33.545 ;
        RECT 87.090 33.445 87.320 34.435 ;
        RECT 79.130 32.725 79.390 33.285 ;
        RECT 79.560 32.920 79.820 33.375 ;
        RECT 79.990 32.725 80.250 33.205 ;
        RECT 80.420 32.920 80.680 33.375 ;
        RECT 80.850 32.725 81.110 33.205 ;
        RECT 81.280 32.920 81.540 33.375 ;
        RECT 81.710 32.725 81.955 33.205 ;
        RECT 82.125 32.920 82.400 33.375 ;
        RECT 82.570 32.725 82.815 33.205 ;
        RECT 82.985 32.920 83.245 33.375 ;
        RECT 83.425 32.725 83.675 33.205 ;
        RECT 83.845 32.920 84.105 33.375 ;
        RECT 84.285 32.725 84.535 33.205 ;
        RECT 84.705 32.920 84.965 33.375 ;
        RECT 85.145 32.725 85.405 33.205 ;
        RECT 85.575 32.920 85.835 33.375 ;
        RECT 86.570 33.275 87.320 33.445 ;
        RECT 86.005 32.725 86.305 33.205 ;
        RECT 86.570 32.985 86.825 33.275 ;
        RECT 86.995 32.725 87.325 33.105 ;
        RECT 87.495 32.985 87.665 35.105 ;
        RECT 87.835 34.305 88.160 35.090 ;
        RECT 88.330 34.815 88.580 35.275 ;
        RECT 88.750 34.775 89.000 35.105 ;
        RECT 89.215 34.775 89.895 35.105 ;
        RECT 88.750 34.645 88.920 34.775 ;
        RECT 88.525 34.475 88.920 34.645 ;
        RECT 87.895 33.255 88.355 34.305 ;
        RECT 88.525 33.115 88.695 34.475 ;
        RECT 89.090 34.215 89.555 34.605 ;
        RECT 88.865 33.405 89.215 34.025 ;
        RECT 89.385 33.625 89.555 34.215 ;
        RECT 89.725 33.995 89.895 34.775 ;
        RECT 90.065 34.675 90.235 35.015 ;
        RECT 90.470 34.845 90.800 35.275 ;
        RECT 90.970 34.675 91.140 35.015 ;
        RECT 91.435 34.815 91.805 35.275 ;
        RECT 90.065 34.505 91.140 34.675 ;
        RECT 91.975 34.645 92.145 35.105 ;
        RECT 92.380 34.765 93.250 35.105 ;
        RECT 93.420 34.815 93.670 35.275 ;
        RECT 91.585 34.475 92.145 34.645 ;
        RECT 91.585 34.335 91.755 34.475 ;
        RECT 90.255 34.165 91.755 34.335 ;
        RECT 92.450 34.305 92.910 34.595 ;
        RECT 89.725 33.825 91.415 33.995 ;
        RECT 89.385 33.405 89.740 33.625 ;
        RECT 89.910 33.115 90.080 33.825 ;
        RECT 90.285 33.405 91.075 33.655 ;
        RECT 91.245 33.645 91.415 33.825 ;
        RECT 91.585 33.475 91.755 34.165 ;
        RECT 88.025 32.725 88.355 33.085 ;
        RECT 88.525 32.945 89.020 33.115 ;
        RECT 89.225 32.945 90.080 33.115 ;
        RECT 90.955 32.725 91.285 33.185 ;
        RECT 91.495 33.085 91.755 33.475 ;
        RECT 91.945 34.295 92.910 34.305 ;
        RECT 93.080 34.385 93.250 34.765 ;
        RECT 93.840 34.725 94.010 35.015 ;
        RECT 94.190 34.895 94.520 35.275 ;
        RECT 93.840 34.555 94.640 34.725 ;
        RECT 91.945 34.135 92.620 34.295 ;
        RECT 93.080 34.215 94.300 34.385 ;
        RECT 91.945 33.345 92.155 34.135 ;
        RECT 93.080 34.125 93.250 34.215 ;
        RECT 92.325 33.345 92.675 33.965 ;
        RECT 92.845 33.955 93.250 34.125 ;
        RECT 92.845 33.175 93.015 33.955 ;
        RECT 93.185 33.505 93.405 33.785 ;
        RECT 93.585 33.675 94.125 34.045 ;
        RECT 94.470 33.965 94.640 34.555 ;
        RECT 94.860 34.135 95.165 35.275 ;
        RECT 95.335 34.085 95.590 34.965 ;
        RECT 95.765 34.110 96.055 35.275 ;
        RECT 96.285 34.135 96.495 35.275 ;
        RECT 96.665 34.125 96.995 35.105 ;
        RECT 97.165 34.135 97.395 35.275 ;
        RECT 97.605 34.185 101.115 35.275 ;
        RECT 101.285 34.185 102.495 35.275 ;
        RECT 94.470 33.935 95.210 33.965 ;
        RECT 93.185 33.335 93.715 33.505 ;
        RECT 91.495 32.915 91.845 33.085 ;
        RECT 92.065 32.895 93.015 33.175 ;
        RECT 93.185 32.725 93.375 33.165 ;
        RECT 93.545 33.105 93.715 33.335 ;
        RECT 93.885 33.275 94.125 33.675 ;
        RECT 94.295 33.635 95.210 33.935 ;
        RECT 94.295 33.460 94.620 33.635 ;
        RECT 94.295 33.105 94.615 33.460 ;
        RECT 95.380 33.435 95.590 34.085 ;
        RECT 93.545 32.935 94.615 33.105 ;
        RECT 94.860 32.725 95.165 33.185 ;
        RECT 95.335 32.905 95.590 33.435 ;
        RECT 95.765 32.725 96.055 33.450 ;
        RECT 96.285 32.725 96.495 33.545 ;
        RECT 96.665 33.525 96.915 34.125 ;
        RECT 97.085 33.715 97.415 33.965 ;
        RECT 96.665 32.895 96.995 33.525 ;
        RECT 97.165 32.725 97.395 33.545 ;
        RECT 97.605 33.495 99.255 34.015 ;
        RECT 99.425 33.665 101.115 34.185 ;
        RECT 97.605 32.725 101.115 33.495 ;
        RECT 101.285 33.475 101.805 34.015 ;
        RECT 101.975 33.645 102.495 34.185 ;
        RECT 102.705 34.135 102.935 35.275 ;
        RECT 103.105 34.125 103.435 35.105 ;
        RECT 103.605 34.135 103.815 35.275 ;
        RECT 104.045 34.840 109.390 35.275 ;
        RECT 109.565 34.840 114.910 35.275 ;
        RECT 102.685 33.715 103.015 33.965 ;
        RECT 101.285 32.725 102.495 33.475 ;
        RECT 102.705 32.725 102.935 33.545 ;
        RECT 103.185 33.525 103.435 34.125 ;
        RECT 103.105 32.895 103.435 33.525 ;
        RECT 103.605 32.725 103.815 33.545 ;
        RECT 105.630 33.270 105.970 34.100 ;
        RECT 107.450 33.590 107.800 34.840 ;
        RECT 111.150 33.270 111.490 34.100 ;
        RECT 112.970 33.590 113.320 34.840 ;
        RECT 115.085 34.185 116.755 35.275 ;
        RECT 115.085 33.495 115.835 34.015 ;
        RECT 116.005 33.665 116.755 34.185 ;
        RECT 117.385 34.185 118.595 35.275 ;
        RECT 117.385 33.645 117.905 34.185 ;
        RECT 104.045 32.725 109.390 33.270 ;
        RECT 109.565 32.725 114.910 33.270 ;
        RECT 115.085 32.725 116.755 33.495 ;
        RECT 118.075 33.475 118.595 34.015 ;
        RECT 117.385 32.725 118.595 33.475 ;
        RECT 5.520 32.555 118.680 32.725 ;
        RECT 5.605 31.805 6.815 32.555 ;
        RECT 6.985 32.010 12.330 32.555 ;
        RECT 5.605 31.265 6.125 31.805 ;
        RECT 6.295 31.095 6.815 31.635 ;
        RECT 8.570 31.180 8.910 32.010 ;
        RECT 12.505 31.805 13.715 32.555 ;
        RECT 13.975 32.005 14.145 32.385 ;
        RECT 14.325 32.175 14.655 32.555 ;
        RECT 13.975 31.835 14.640 32.005 ;
        RECT 14.835 31.880 15.095 32.385 ;
        RECT 5.605 30.005 6.815 31.095 ;
        RECT 10.390 30.440 10.740 31.690 ;
        RECT 12.505 31.265 13.025 31.805 ;
        RECT 13.195 31.095 13.715 31.635 ;
        RECT 13.905 31.285 14.235 31.655 ;
        RECT 14.470 31.580 14.640 31.835 ;
        RECT 14.470 31.250 14.755 31.580 ;
        RECT 14.470 31.105 14.640 31.250 ;
        RECT 6.985 30.005 12.330 30.440 ;
        RECT 12.505 30.005 13.715 31.095 ;
        RECT 13.975 30.935 14.640 31.105 ;
        RECT 14.925 31.080 15.095 31.880 ;
        RECT 15.270 32.005 15.525 32.295 ;
        RECT 15.695 32.175 16.025 32.555 ;
        RECT 15.270 31.835 16.020 32.005 ;
        RECT 13.975 30.175 14.145 30.935 ;
        RECT 14.325 30.005 14.655 30.765 ;
        RECT 14.825 30.175 15.095 31.080 ;
        RECT 15.270 31.015 15.620 31.665 ;
        RECT 15.790 30.845 16.020 31.835 ;
        RECT 15.270 30.675 16.020 30.845 ;
        RECT 15.270 30.175 15.525 30.675 ;
        RECT 15.695 30.005 16.025 30.505 ;
        RECT 16.195 30.175 16.365 32.295 ;
        RECT 16.725 32.195 17.055 32.555 ;
        RECT 17.225 32.165 17.720 32.335 ;
        RECT 17.925 32.165 18.780 32.335 ;
        RECT 16.595 30.975 17.055 32.025 ;
        RECT 16.535 30.190 16.860 30.975 ;
        RECT 17.225 30.805 17.395 32.165 ;
        RECT 17.565 31.255 17.915 31.875 ;
        RECT 18.085 31.655 18.440 31.875 ;
        RECT 18.085 31.065 18.255 31.655 ;
        RECT 18.610 31.455 18.780 32.165 ;
        RECT 19.655 32.095 19.985 32.555 ;
        RECT 20.195 32.195 20.545 32.365 ;
        RECT 18.985 31.625 19.775 31.875 ;
        RECT 20.195 31.805 20.455 32.195 ;
        RECT 20.765 32.105 21.715 32.385 ;
        RECT 21.885 32.115 22.075 32.555 ;
        RECT 22.245 32.175 23.315 32.345 ;
        RECT 19.945 31.455 20.115 31.635 ;
        RECT 17.225 30.635 17.620 30.805 ;
        RECT 17.790 30.675 18.255 31.065 ;
        RECT 18.425 31.285 20.115 31.455 ;
        RECT 17.450 30.505 17.620 30.635 ;
        RECT 18.425 30.505 18.595 31.285 ;
        RECT 20.285 31.115 20.455 31.805 ;
        RECT 18.955 30.945 20.455 31.115 ;
        RECT 20.645 31.145 20.855 31.935 ;
        RECT 21.025 31.315 21.375 31.935 ;
        RECT 21.545 31.325 21.715 32.105 ;
        RECT 22.245 31.945 22.415 32.175 ;
        RECT 21.885 31.775 22.415 31.945 ;
        RECT 21.885 31.495 22.105 31.775 ;
        RECT 22.585 31.605 22.825 32.005 ;
        RECT 21.545 31.155 21.950 31.325 ;
        RECT 22.285 31.235 22.825 31.605 ;
        RECT 22.995 31.820 23.315 32.175 ;
        RECT 23.560 32.095 23.865 32.555 ;
        RECT 24.035 31.845 24.290 32.375 ;
        RECT 22.995 31.645 23.320 31.820 ;
        RECT 22.995 31.345 23.910 31.645 ;
        RECT 23.170 31.315 23.910 31.345 ;
        RECT 20.645 30.985 21.320 31.145 ;
        RECT 21.780 31.065 21.950 31.155 ;
        RECT 20.645 30.975 21.610 30.985 ;
        RECT 20.285 30.805 20.455 30.945 ;
        RECT 17.030 30.005 17.280 30.465 ;
        RECT 17.450 30.175 17.700 30.505 ;
        RECT 17.915 30.175 18.595 30.505 ;
        RECT 18.765 30.605 19.840 30.775 ;
        RECT 20.285 30.635 20.845 30.805 ;
        RECT 21.150 30.685 21.610 30.975 ;
        RECT 21.780 30.895 23.000 31.065 ;
        RECT 18.765 30.265 18.935 30.605 ;
        RECT 19.170 30.005 19.500 30.435 ;
        RECT 19.670 30.265 19.840 30.605 ;
        RECT 20.135 30.005 20.505 30.465 ;
        RECT 20.675 30.175 20.845 30.635 ;
        RECT 21.780 30.515 21.950 30.895 ;
        RECT 23.170 30.725 23.340 31.315 ;
        RECT 24.080 31.195 24.290 31.845 ;
        RECT 21.080 30.175 21.950 30.515 ;
        RECT 22.540 30.555 23.340 30.725 ;
        RECT 22.120 30.005 22.370 30.465 ;
        RECT 22.540 30.265 22.710 30.555 ;
        RECT 22.890 30.005 23.220 30.385 ;
        RECT 23.560 30.005 23.865 31.145 ;
        RECT 24.035 30.315 24.290 31.195 ;
        RECT 24.470 31.815 24.725 32.385 ;
        RECT 24.895 32.155 25.225 32.555 ;
        RECT 25.650 32.020 26.180 32.385 ;
        RECT 25.650 31.985 25.825 32.020 ;
        RECT 24.895 31.815 25.825 31.985 ;
        RECT 24.470 31.145 24.640 31.815 ;
        RECT 24.895 31.645 25.065 31.815 ;
        RECT 24.810 31.315 25.065 31.645 ;
        RECT 25.290 31.315 25.485 31.645 ;
        RECT 24.470 30.175 24.805 31.145 ;
        RECT 24.975 30.005 25.145 31.145 ;
        RECT 25.315 30.345 25.485 31.315 ;
        RECT 25.655 30.685 25.825 31.815 ;
        RECT 25.995 31.025 26.165 31.825 ;
        RECT 26.370 31.535 26.645 32.385 ;
        RECT 26.365 31.365 26.645 31.535 ;
        RECT 26.370 31.225 26.645 31.365 ;
        RECT 26.815 31.025 27.005 32.385 ;
        RECT 27.185 32.020 27.695 32.555 ;
        RECT 27.915 31.745 28.160 32.350 ;
        RECT 28.605 31.805 29.815 32.555 ;
        RECT 29.985 31.880 30.245 32.385 ;
        RECT 30.425 32.175 30.755 32.555 ;
        RECT 30.935 32.005 31.105 32.385 ;
        RECT 27.205 31.575 28.435 31.745 ;
        RECT 25.995 30.855 27.005 31.025 ;
        RECT 27.175 31.010 27.925 31.200 ;
        RECT 25.655 30.515 26.780 30.685 ;
        RECT 27.175 30.345 27.345 31.010 ;
        RECT 28.095 30.765 28.435 31.575 ;
        RECT 28.605 31.265 29.125 31.805 ;
        RECT 29.295 31.095 29.815 31.635 ;
        RECT 25.315 30.175 27.345 30.345 ;
        RECT 27.515 30.005 27.685 30.765 ;
        RECT 27.920 30.355 28.435 30.765 ;
        RECT 28.605 30.005 29.815 31.095 ;
        RECT 29.985 31.080 30.155 31.880 ;
        RECT 30.440 31.835 31.105 32.005 ;
        RECT 30.440 31.580 30.610 31.835 ;
        RECT 31.365 31.830 31.655 32.555 ;
        RECT 31.830 31.815 32.085 32.385 ;
        RECT 32.255 32.155 32.585 32.555 ;
        RECT 33.010 32.020 33.540 32.385 ;
        RECT 33.010 31.985 33.185 32.020 ;
        RECT 32.255 31.815 33.185 31.985 ;
        RECT 30.325 31.250 30.610 31.580 ;
        RECT 30.845 31.285 31.175 31.655 ;
        RECT 30.440 31.105 30.610 31.250 ;
        RECT 29.985 30.175 30.255 31.080 ;
        RECT 30.440 30.935 31.105 31.105 ;
        RECT 30.425 30.005 30.755 30.765 ;
        RECT 30.935 30.175 31.105 30.935 ;
        RECT 31.365 30.005 31.655 31.170 ;
        RECT 31.830 31.145 32.000 31.815 ;
        RECT 32.255 31.645 32.425 31.815 ;
        RECT 32.170 31.315 32.425 31.645 ;
        RECT 32.650 31.315 32.845 31.645 ;
        RECT 31.830 30.175 32.165 31.145 ;
        RECT 32.335 30.005 32.505 31.145 ;
        RECT 32.675 30.345 32.845 31.315 ;
        RECT 33.015 30.685 33.185 31.815 ;
        RECT 33.355 31.025 33.525 31.825 ;
        RECT 33.730 31.535 34.005 32.385 ;
        RECT 33.725 31.365 34.005 31.535 ;
        RECT 33.730 31.225 34.005 31.365 ;
        RECT 34.175 31.025 34.365 32.385 ;
        RECT 34.545 32.020 35.055 32.555 ;
        RECT 35.275 31.745 35.520 32.350 ;
        RECT 36.445 32.085 36.740 32.555 ;
        RECT 36.910 31.915 37.170 32.360 ;
        RECT 37.340 32.085 37.600 32.555 ;
        RECT 37.770 31.915 38.025 32.360 ;
        RECT 38.195 32.085 38.495 32.555 ;
        RECT 35.985 31.745 39.015 31.915 ;
        RECT 34.565 31.575 35.795 31.745 ;
        RECT 33.355 30.855 34.365 31.025 ;
        RECT 34.535 31.010 35.285 31.200 ;
        RECT 33.015 30.515 34.140 30.685 ;
        RECT 34.535 30.345 34.705 31.010 ;
        RECT 35.455 30.765 35.795 31.575 ;
        RECT 35.985 31.180 36.155 31.745 ;
        RECT 36.325 31.350 38.540 31.575 ;
        RECT 38.715 31.180 39.015 31.745 ;
        RECT 35.985 31.010 39.015 31.180 ;
        RECT 39.185 31.880 39.445 32.385 ;
        RECT 39.625 32.175 39.955 32.555 ;
        RECT 40.135 32.005 40.305 32.385 ;
        RECT 39.185 31.080 39.355 31.880 ;
        RECT 39.640 31.835 40.305 32.005 ;
        RECT 40.655 32.005 40.825 32.295 ;
        RECT 40.995 32.175 41.325 32.555 ;
        RECT 40.655 31.835 41.320 32.005 ;
        RECT 39.640 31.580 39.810 31.835 ;
        RECT 39.525 31.250 39.810 31.580 ;
        RECT 40.045 31.285 40.375 31.655 ;
        RECT 39.640 31.105 39.810 31.250 ;
        RECT 32.675 30.175 34.705 30.345 ;
        RECT 34.875 30.005 35.045 30.765 ;
        RECT 35.280 30.355 35.795 30.765 ;
        RECT 35.965 30.005 36.310 30.840 ;
        RECT 36.485 30.205 36.740 31.010 ;
        RECT 36.910 30.005 37.170 30.840 ;
        RECT 37.345 30.205 37.600 31.010 ;
        RECT 37.770 30.005 38.030 30.840 ;
        RECT 38.200 30.205 38.460 31.010 ;
        RECT 38.630 30.005 39.015 30.840 ;
        RECT 39.185 30.175 39.455 31.080 ;
        RECT 39.640 30.935 40.305 31.105 ;
        RECT 40.570 31.015 40.920 31.665 ;
        RECT 39.625 30.005 39.955 30.765 ;
        RECT 40.135 30.175 40.305 30.935 ;
        RECT 41.090 30.845 41.320 31.835 ;
        RECT 40.655 30.675 41.320 30.845 ;
        RECT 40.655 30.175 40.825 30.675 ;
        RECT 40.995 30.005 41.325 30.505 ;
        RECT 41.495 30.175 41.720 32.295 ;
        RECT 41.935 32.175 42.265 32.555 ;
        RECT 42.435 32.005 42.605 32.335 ;
        RECT 42.905 32.175 43.920 32.375 ;
        RECT 41.910 31.815 42.605 32.005 ;
        RECT 41.910 30.845 42.080 31.815 ;
        RECT 42.250 31.015 42.660 31.635 ;
        RECT 42.830 31.065 43.050 31.935 ;
        RECT 43.230 31.625 43.580 31.995 ;
        RECT 43.750 31.445 43.920 32.175 ;
        RECT 44.090 32.115 44.500 32.555 ;
        RECT 44.790 31.915 45.040 32.345 ;
        RECT 45.240 32.095 45.560 32.555 ;
        RECT 46.120 32.165 46.970 32.335 ;
        RECT 44.090 31.575 44.500 31.905 ;
        RECT 44.790 31.575 45.210 31.915 ;
        RECT 43.500 31.405 43.920 31.445 ;
        RECT 43.500 31.235 44.850 31.405 ;
        RECT 41.910 30.675 42.605 30.845 ;
        RECT 42.830 30.685 43.330 31.065 ;
        RECT 41.935 30.005 42.265 30.505 ;
        RECT 42.435 30.175 42.605 30.675 ;
        RECT 43.500 30.390 43.670 31.235 ;
        RECT 44.600 31.075 44.850 31.235 ;
        RECT 43.840 30.805 44.090 31.065 ;
        RECT 45.020 30.805 45.210 31.575 ;
        RECT 43.840 30.555 45.210 30.805 ;
        RECT 45.380 31.745 46.630 31.915 ;
        RECT 45.380 30.985 45.550 31.745 ;
        RECT 46.300 31.625 46.630 31.745 ;
        RECT 45.720 31.165 45.900 31.575 ;
        RECT 46.800 31.405 46.970 32.165 ;
        RECT 47.170 32.075 47.830 32.555 ;
        RECT 48.010 31.960 48.330 32.290 ;
        RECT 47.160 31.635 47.820 31.905 ;
        RECT 47.160 31.575 47.490 31.635 ;
        RECT 47.640 31.405 47.970 31.465 ;
        RECT 46.070 31.235 47.970 31.405 ;
        RECT 45.380 30.675 45.900 30.985 ;
        RECT 46.070 30.725 46.240 31.235 ;
        RECT 48.140 31.065 48.330 31.960 ;
        RECT 46.410 30.895 48.330 31.065 ;
        RECT 48.010 30.875 48.330 30.895 ;
        RECT 48.530 31.645 48.780 32.295 ;
        RECT 48.960 32.095 49.245 32.555 ;
        RECT 49.425 32.215 49.680 32.375 ;
        RECT 49.425 32.045 49.765 32.215 ;
        RECT 49.425 31.845 49.680 32.045 ;
        RECT 48.530 31.315 49.330 31.645 ;
        RECT 46.070 30.555 47.280 30.725 ;
        RECT 42.840 30.220 43.670 30.390 ;
        RECT 43.910 30.005 44.290 30.385 ;
        RECT 44.470 30.265 44.640 30.555 ;
        RECT 46.070 30.475 46.240 30.555 ;
        RECT 44.810 30.005 45.140 30.385 ;
        RECT 45.610 30.225 46.240 30.475 ;
        RECT 46.420 30.005 46.840 30.385 ;
        RECT 47.040 30.265 47.280 30.555 ;
        RECT 47.510 30.005 47.840 30.695 ;
        RECT 48.010 30.265 48.180 30.875 ;
        RECT 48.530 30.725 48.780 31.315 ;
        RECT 49.500 30.985 49.680 31.845 ;
        RECT 50.225 31.785 53.735 32.555 ;
        RECT 54.825 31.815 55.520 32.385 ;
        RECT 55.690 31.815 56.040 32.340 ;
        RECT 50.225 31.265 51.875 31.785 ;
        RECT 52.045 31.095 53.735 31.615 ;
        RECT 48.450 30.215 48.780 30.725 ;
        RECT 48.960 30.005 49.245 30.805 ;
        RECT 49.425 30.315 49.680 30.985 ;
        RECT 50.225 30.005 53.735 31.095 ;
        RECT 54.825 30.975 55.065 31.645 ;
        RECT 55.245 31.145 55.415 31.815 ;
        RECT 55.690 31.645 55.895 31.815 ;
        RECT 56.230 31.645 56.445 32.340 ;
        RECT 56.615 31.815 56.950 32.555 ;
        RECT 57.125 31.830 57.415 32.555 ;
        RECT 57.585 31.805 58.795 32.555 ;
        RECT 58.965 31.815 59.430 32.360 ;
        RECT 55.585 31.315 55.895 31.645 ;
        RECT 56.065 31.315 56.445 31.645 ;
        RECT 56.645 31.315 56.930 31.645 ;
        RECT 57.585 31.265 58.105 31.805 ;
        RECT 55.245 30.975 56.525 31.145 ;
        RECT 54.845 30.005 55.125 30.805 ;
        RECT 55.325 30.175 55.655 30.975 ;
        RECT 55.855 30.005 56.025 30.805 ;
        RECT 56.195 30.175 56.525 30.975 ;
        RECT 56.695 30.005 56.955 31.145 ;
        RECT 57.125 30.005 57.415 31.170 ;
        RECT 58.275 31.095 58.795 31.635 ;
        RECT 57.585 30.005 58.795 31.095 ;
        RECT 58.965 30.855 59.135 31.815 ;
        RECT 59.935 31.735 60.105 32.555 ;
        RECT 60.275 31.905 60.605 32.385 ;
        RECT 60.775 32.165 61.125 32.555 ;
        RECT 61.295 31.985 61.525 32.385 ;
        RECT 61.015 31.905 61.525 31.985 ;
        RECT 60.275 31.815 61.525 31.905 ;
        RECT 61.695 31.815 62.015 32.295 ;
        RECT 62.190 32.005 62.445 32.295 ;
        RECT 62.615 32.175 62.945 32.555 ;
        RECT 62.190 31.835 62.940 32.005 ;
        RECT 60.275 31.735 61.185 31.815 ;
        RECT 59.305 31.195 59.550 31.645 ;
        RECT 59.810 31.365 60.505 31.565 ;
        RECT 60.675 31.395 61.275 31.565 ;
        RECT 60.675 31.195 60.845 31.395 ;
        RECT 61.505 31.225 61.675 31.645 ;
        RECT 59.305 31.025 60.845 31.195 ;
        RECT 61.015 31.055 61.675 31.225 ;
        RECT 61.015 30.855 61.185 31.055 ;
        RECT 61.845 30.885 62.015 31.815 ;
        RECT 62.190 31.015 62.540 31.665 ;
        RECT 58.965 30.685 61.185 30.855 ;
        RECT 61.355 30.685 62.015 30.885 ;
        RECT 62.710 30.845 62.940 31.835 ;
        RECT 58.965 30.005 59.265 30.515 ;
        RECT 59.435 30.175 59.765 30.685 ;
        RECT 61.355 30.515 61.525 30.685 ;
        RECT 62.190 30.675 62.940 30.845 ;
        RECT 59.935 30.005 60.565 30.515 ;
        RECT 61.145 30.345 61.525 30.515 ;
        RECT 61.695 30.005 61.995 30.515 ;
        RECT 62.190 30.175 62.445 30.675 ;
        RECT 62.615 30.005 62.945 30.505 ;
        RECT 63.115 30.175 63.285 32.295 ;
        RECT 63.645 32.195 63.975 32.555 ;
        RECT 64.145 32.165 64.640 32.335 ;
        RECT 64.845 32.165 65.700 32.335 ;
        RECT 63.515 30.975 63.975 32.025 ;
        RECT 63.455 30.190 63.780 30.975 ;
        RECT 64.145 30.805 64.315 32.165 ;
        RECT 64.485 31.255 64.835 31.875 ;
        RECT 65.005 31.655 65.360 31.875 ;
        RECT 65.005 31.065 65.175 31.655 ;
        RECT 65.530 31.455 65.700 32.165 ;
        RECT 66.575 32.095 66.905 32.555 ;
        RECT 67.115 32.195 67.465 32.365 ;
        RECT 65.905 31.625 66.695 31.875 ;
        RECT 67.115 31.805 67.375 32.195 ;
        RECT 67.685 32.105 68.635 32.385 ;
        RECT 68.805 32.115 68.995 32.555 ;
        RECT 69.165 32.175 70.235 32.345 ;
        RECT 66.865 31.455 67.035 31.635 ;
        RECT 64.145 30.635 64.540 30.805 ;
        RECT 64.710 30.675 65.175 31.065 ;
        RECT 65.345 31.285 67.035 31.455 ;
        RECT 64.370 30.505 64.540 30.635 ;
        RECT 65.345 30.505 65.515 31.285 ;
        RECT 67.205 31.115 67.375 31.805 ;
        RECT 65.875 30.945 67.375 31.115 ;
        RECT 67.565 31.145 67.775 31.935 ;
        RECT 67.945 31.315 68.295 31.935 ;
        RECT 68.465 31.325 68.635 32.105 ;
        RECT 69.165 31.945 69.335 32.175 ;
        RECT 68.805 31.775 69.335 31.945 ;
        RECT 68.805 31.495 69.025 31.775 ;
        RECT 69.505 31.605 69.745 32.005 ;
        RECT 68.465 31.155 68.870 31.325 ;
        RECT 69.205 31.235 69.745 31.605 ;
        RECT 69.915 31.820 70.235 32.175 ;
        RECT 70.480 32.095 70.785 32.555 ;
        RECT 70.955 31.845 71.205 32.375 ;
        RECT 69.915 31.645 70.240 31.820 ;
        RECT 69.915 31.345 70.830 31.645 ;
        RECT 70.090 31.315 70.830 31.345 ;
        RECT 67.565 30.985 68.240 31.145 ;
        RECT 68.700 31.065 68.870 31.155 ;
        RECT 67.565 30.975 68.530 30.985 ;
        RECT 67.205 30.805 67.375 30.945 ;
        RECT 63.950 30.005 64.200 30.465 ;
        RECT 64.370 30.175 64.620 30.505 ;
        RECT 64.835 30.175 65.515 30.505 ;
        RECT 65.685 30.605 66.760 30.775 ;
        RECT 67.205 30.635 67.765 30.805 ;
        RECT 68.070 30.685 68.530 30.975 ;
        RECT 68.700 30.895 69.920 31.065 ;
        RECT 65.685 30.265 65.855 30.605 ;
        RECT 66.090 30.005 66.420 30.435 ;
        RECT 66.590 30.265 66.760 30.605 ;
        RECT 67.055 30.005 67.425 30.465 ;
        RECT 67.595 30.175 67.765 30.635 ;
        RECT 68.700 30.515 68.870 30.895 ;
        RECT 70.090 30.725 70.260 31.315 ;
        RECT 71.000 31.195 71.205 31.845 ;
        RECT 71.375 31.800 71.625 32.555 ;
        RECT 71.850 32.005 72.105 32.295 ;
        RECT 72.275 32.175 72.605 32.555 ;
        RECT 71.850 31.835 72.600 32.005 ;
        RECT 68.000 30.175 68.870 30.515 ;
        RECT 69.460 30.555 70.260 30.725 ;
        RECT 69.040 30.005 69.290 30.465 ;
        RECT 69.460 30.265 69.630 30.555 ;
        RECT 69.810 30.005 70.140 30.385 ;
        RECT 70.480 30.005 70.785 31.145 ;
        RECT 70.955 30.315 71.205 31.195 ;
        RECT 71.375 30.005 71.625 31.145 ;
        RECT 71.850 31.015 72.200 31.665 ;
        RECT 72.370 30.845 72.600 31.835 ;
        RECT 71.850 30.675 72.600 30.845 ;
        RECT 71.850 30.175 72.105 30.675 ;
        RECT 72.275 30.005 72.605 30.505 ;
        RECT 72.775 30.175 72.945 32.295 ;
        RECT 73.305 32.195 73.635 32.555 ;
        RECT 73.805 32.165 74.300 32.335 ;
        RECT 74.505 32.165 75.360 32.335 ;
        RECT 73.175 30.975 73.635 32.025 ;
        RECT 73.115 30.190 73.440 30.975 ;
        RECT 73.805 30.805 73.975 32.165 ;
        RECT 74.145 31.255 74.495 31.875 ;
        RECT 74.665 31.655 75.020 31.875 ;
        RECT 74.665 31.065 74.835 31.655 ;
        RECT 75.190 31.455 75.360 32.165 ;
        RECT 76.235 32.095 76.565 32.555 ;
        RECT 76.775 32.195 77.125 32.365 ;
        RECT 75.565 31.625 76.355 31.875 ;
        RECT 76.775 31.805 77.035 32.195 ;
        RECT 77.345 32.105 78.295 32.385 ;
        RECT 78.465 32.115 78.655 32.555 ;
        RECT 78.825 32.175 79.895 32.345 ;
        RECT 76.525 31.455 76.695 31.635 ;
        RECT 73.805 30.635 74.200 30.805 ;
        RECT 74.370 30.675 74.835 31.065 ;
        RECT 75.005 31.285 76.695 31.455 ;
        RECT 74.030 30.505 74.200 30.635 ;
        RECT 75.005 30.505 75.175 31.285 ;
        RECT 76.865 31.115 77.035 31.805 ;
        RECT 75.535 30.945 77.035 31.115 ;
        RECT 77.225 31.145 77.435 31.935 ;
        RECT 77.605 31.315 77.955 31.935 ;
        RECT 78.125 31.325 78.295 32.105 ;
        RECT 78.825 31.945 78.995 32.175 ;
        RECT 78.465 31.775 78.995 31.945 ;
        RECT 78.465 31.495 78.685 31.775 ;
        RECT 79.165 31.605 79.405 32.005 ;
        RECT 78.125 31.155 78.530 31.325 ;
        RECT 78.865 31.235 79.405 31.605 ;
        RECT 79.575 31.820 79.895 32.175 ;
        RECT 80.140 32.095 80.445 32.555 ;
        RECT 80.615 31.845 80.870 32.375 ;
        RECT 79.575 31.645 79.900 31.820 ;
        RECT 79.575 31.345 80.490 31.645 ;
        RECT 79.750 31.315 80.490 31.345 ;
        RECT 77.225 30.985 77.900 31.145 ;
        RECT 78.360 31.065 78.530 31.155 ;
        RECT 77.225 30.975 78.190 30.985 ;
        RECT 76.865 30.805 77.035 30.945 ;
        RECT 73.610 30.005 73.860 30.465 ;
        RECT 74.030 30.175 74.280 30.505 ;
        RECT 74.495 30.175 75.175 30.505 ;
        RECT 75.345 30.605 76.420 30.775 ;
        RECT 76.865 30.635 77.425 30.805 ;
        RECT 77.730 30.685 78.190 30.975 ;
        RECT 78.360 30.895 79.580 31.065 ;
        RECT 75.345 30.265 75.515 30.605 ;
        RECT 75.750 30.005 76.080 30.435 ;
        RECT 76.250 30.265 76.420 30.605 ;
        RECT 76.715 30.005 77.085 30.465 ;
        RECT 77.255 30.175 77.425 30.635 ;
        RECT 78.360 30.515 78.530 30.895 ;
        RECT 79.750 30.725 79.920 31.315 ;
        RECT 80.660 31.195 80.870 31.845 ;
        RECT 81.135 32.005 81.305 32.385 ;
        RECT 81.485 32.175 81.815 32.555 ;
        RECT 81.135 31.835 81.800 32.005 ;
        RECT 81.995 31.880 82.255 32.385 ;
        RECT 81.065 31.285 81.395 31.655 ;
        RECT 81.630 31.580 81.800 31.835 ;
        RECT 77.660 30.175 78.530 30.515 ;
        RECT 79.120 30.555 79.920 30.725 ;
        RECT 78.700 30.005 78.950 30.465 ;
        RECT 79.120 30.265 79.290 30.555 ;
        RECT 79.470 30.005 79.800 30.385 ;
        RECT 80.140 30.005 80.445 31.145 ;
        RECT 80.615 30.315 80.870 31.195 ;
        RECT 81.630 31.250 81.915 31.580 ;
        RECT 81.630 31.105 81.800 31.250 ;
        RECT 81.135 30.935 81.800 31.105 ;
        RECT 82.085 31.080 82.255 31.880 ;
        RECT 82.885 31.830 83.175 32.555 ;
        RECT 83.350 31.815 83.605 32.385 ;
        RECT 83.775 32.155 84.105 32.555 ;
        RECT 84.530 32.020 85.060 32.385 ;
        RECT 84.530 31.985 84.705 32.020 ;
        RECT 83.775 31.815 84.705 31.985 ;
        RECT 81.135 30.175 81.305 30.935 ;
        RECT 81.485 30.005 81.815 30.765 ;
        RECT 81.985 30.175 82.255 31.080 ;
        RECT 82.885 30.005 83.175 31.170 ;
        RECT 83.350 31.145 83.520 31.815 ;
        RECT 83.775 31.645 83.945 31.815 ;
        RECT 83.690 31.315 83.945 31.645 ;
        RECT 84.170 31.315 84.365 31.645 ;
        RECT 83.350 30.175 83.685 31.145 ;
        RECT 83.855 30.005 84.025 31.145 ;
        RECT 84.195 30.345 84.365 31.315 ;
        RECT 84.535 30.685 84.705 31.815 ;
        RECT 84.875 31.025 85.045 31.825 ;
        RECT 85.250 31.535 85.525 32.385 ;
        RECT 85.245 31.365 85.525 31.535 ;
        RECT 85.250 31.225 85.525 31.365 ;
        RECT 85.695 31.025 85.885 32.385 ;
        RECT 86.065 32.020 86.575 32.555 ;
        RECT 86.795 31.745 87.040 32.350 ;
        RECT 87.575 32.005 87.745 32.295 ;
        RECT 87.915 32.175 88.245 32.555 ;
        RECT 87.575 31.835 88.240 32.005 ;
        RECT 86.085 31.575 87.315 31.745 ;
        RECT 84.875 30.855 85.885 31.025 ;
        RECT 86.055 31.010 86.805 31.200 ;
        RECT 84.535 30.515 85.660 30.685 ;
        RECT 86.055 30.345 86.225 31.010 ;
        RECT 86.975 30.765 87.315 31.575 ;
        RECT 87.490 31.015 87.840 31.665 ;
        RECT 88.010 30.845 88.240 31.835 ;
        RECT 84.195 30.175 86.225 30.345 ;
        RECT 86.395 30.005 86.565 30.765 ;
        RECT 86.800 30.355 87.315 30.765 ;
        RECT 87.575 30.675 88.240 30.845 ;
        RECT 87.575 30.175 87.745 30.675 ;
        RECT 87.915 30.005 88.245 30.505 ;
        RECT 88.415 30.175 88.640 32.295 ;
        RECT 88.855 32.175 89.185 32.555 ;
        RECT 89.355 32.005 89.525 32.335 ;
        RECT 89.825 32.175 90.840 32.375 ;
        RECT 88.830 31.815 89.525 32.005 ;
        RECT 88.830 30.845 89.000 31.815 ;
        RECT 89.170 31.015 89.580 31.635 ;
        RECT 89.750 31.065 89.970 31.935 ;
        RECT 90.150 31.625 90.500 31.995 ;
        RECT 90.670 31.445 90.840 32.175 ;
        RECT 91.010 32.115 91.420 32.555 ;
        RECT 91.710 31.915 91.960 32.345 ;
        RECT 92.160 32.095 92.480 32.555 ;
        RECT 93.040 32.165 93.890 32.335 ;
        RECT 91.010 31.575 91.420 31.905 ;
        RECT 91.710 31.575 92.130 31.915 ;
        RECT 90.420 31.405 90.840 31.445 ;
        RECT 90.420 31.235 91.770 31.405 ;
        RECT 88.830 30.675 89.525 30.845 ;
        RECT 89.750 30.685 90.250 31.065 ;
        RECT 88.855 30.005 89.185 30.505 ;
        RECT 89.355 30.175 89.525 30.675 ;
        RECT 90.420 30.390 90.590 31.235 ;
        RECT 91.520 31.075 91.770 31.235 ;
        RECT 90.760 30.805 91.010 31.065 ;
        RECT 91.940 30.805 92.130 31.575 ;
        RECT 90.760 30.555 92.130 30.805 ;
        RECT 92.300 31.745 93.550 31.915 ;
        RECT 92.300 30.985 92.470 31.745 ;
        RECT 93.220 31.625 93.550 31.745 ;
        RECT 92.640 31.165 92.820 31.575 ;
        RECT 93.720 31.405 93.890 32.165 ;
        RECT 94.090 32.075 94.750 32.555 ;
        RECT 94.930 31.960 95.250 32.290 ;
        RECT 94.080 31.635 94.740 31.905 ;
        RECT 94.080 31.575 94.410 31.635 ;
        RECT 94.560 31.405 94.890 31.465 ;
        RECT 92.990 31.235 94.890 31.405 ;
        RECT 92.300 30.675 92.820 30.985 ;
        RECT 92.990 30.725 93.160 31.235 ;
        RECT 95.060 31.065 95.250 31.960 ;
        RECT 93.330 30.895 95.250 31.065 ;
        RECT 94.930 30.875 95.250 30.895 ;
        RECT 95.450 31.645 95.700 32.295 ;
        RECT 95.880 32.095 96.165 32.555 ;
        RECT 96.345 31.845 96.600 32.375 ;
        RECT 97.145 32.010 102.490 32.555 ;
        RECT 102.665 32.010 108.010 32.555 ;
        RECT 95.450 31.315 96.250 31.645 ;
        RECT 92.990 30.555 94.200 30.725 ;
        RECT 89.760 30.220 90.590 30.390 ;
        RECT 90.830 30.005 91.210 30.385 ;
        RECT 91.390 30.265 91.560 30.555 ;
        RECT 92.990 30.475 93.160 30.555 ;
        RECT 91.730 30.005 92.060 30.385 ;
        RECT 92.530 30.225 93.160 30.475 ;
        RECT 93.340 30.005 93.760 30.385 ;
        RECT 93.960 30.265 94.200 30.555 ;
        RECT 94.430 30.005 94.760 30.695 ;
        RECT 94.930 30.265 95.100 30.875 ;
        RECT 95.450 30.725 95.700 31.315 ;
        RECT 96.420 31.195 96.600 31.845 ;
        RECT 96.420 31.025 96.685 31.195 ;
        RECT 98.730 31.180 99.070 32.010 ;
        RECT 96.420 30.985 96.600 31.025 ;
        RECT 95.370 30.215 95.700 30.725 ;
        RECT 95.880 30.005 96.165 30.805 ;
        RECT 96.345 30.315 96.600 30.985 ;
        RECT 100.550 30.440 100.900 31.690 ;
        RECT 104.250 31.180 104.590 32.010 ;
        RECT 108.645 31.830 108.935 32.555 ;
        RECT 109.105 32.010 114.450 32.555 ;
        RECT 106.070 30.440 106.420 31.690 ;
        RECT 110.690 31.180 111.030 32.010 ;
        RECT 114.625 31.785 117.215 32.555 ;
        RECT 117.385 31.805 118.595 32.555 ;
        RECT 97.145 30.005 102.490 30.440 ;
        RECT 102.665 30.005 108.010 30.440 ;
        RECT 108.645 30.005 108.935 31.170 ;
        RECT 112.510 30.440 112.860 31.690 ;
        RECT 114.625 31.265 115.835 31.785 ;
        RECT 116.005 31.095 117.215 31.615 ;
        RECT 109.105 30.005 114.450 30.440 ;
        RECT 114.625 30.005 117.215 31.095 ;
        RECT 117.385 31.095 117.905 31.635 ;
        RECT 118.075 31.265 118.595 31.805 ;
        RECT 117.385 30.005 118.595 31.095 ;
        RECT 5.520 29.835 118.680 30.005 ;
        RECT 5.605 28.745 6.815 29.835 ;
        RECT 6.985 29.400 12.330 29.835 ;
        RECT 5.605 28.035 6.125 28.575 ;
        RECT 6.295 28.205 6.815 28.745 ;
        RECT 5.605 27.285 6.815 28.035 ;
        RECT 8.570 27.830 8.910 28.660 ;
        RECT 10.390 28.150 10.740 29.400 ;
        RECT 12.505 28.745 16.015 29.835 ;
        RECT 12.505 28.055 14.155 28.575 ;
        RECT 14.325 28.225 16.015 28.745 ;
        RECT 17.145 28.695 17.375 29.835 ;
        RECT 17.545 28.685 17.875 29.665 ;
        RECT 18.045 28.695 18.255 29.835 ;
        RECT 17.125 28.275 17.455 28.525 ;
        RECT 6.985 27.285 12.330 27.830 ;
        RECT 12.505 27.285 16.015 28.055 ;
        RECT 17.145 27.285 17.375 28.105 ;
        RECT 17.625 28.085 17.875 28.685 ;
        RECT 18.485 28.670 18.775 29.835 ;
        RECT 18.950 28.695 19.285 29.665 ;
        RECT 19.455 28.695 19.625 29.835 ;
        RECT 19.795 29.495 21.825 29.665 ;
        RECT 17.545 27.455 17.875 28.085 ;
        RECT 18.045 27.285 18.255 28.105 ;
        RECT 18.950 28.025 19.120 28.695 ;
        RECT 19.795 28.525 19.965 29.495 ;
        RECT 19.290 28.195 19.545 28.525 ;
        RECT 19.770 28.195 19.965 28.525 ;
        RECT 20.135 29.155 21.260 29.325 ;
        RECT 19.375 28.025 19.545 28.195 ;
        RECT 20.135 28.025 20.305 29.155 ;
        RECT 18.485 27.285 18.775 28.010 ;
        RECT 18.950 27.455 19.205 28.025 ;
        RECT 19.375 27.855 20.305 28.025 ;
        RECT 20.475 28.815 21.485 28.985 ;
        RECT 20.475 28.015 20.645 28.815 ;
        RECT 20.130 27.820 20.305 27.855 ;
        RECT 19.375 27.285 19.705 27.685 ;
        RECT 20.130 27.455 20.660 27.820 ;
        RECT 20.850 27.795 21.125 28.615 ;
        RECT 20.845 27.625 21.125 27.795 ;
        RECT 20.850 27.455 21.125 27.625 ;
        RECT 21.295 27.455 21.485 28.815 ;
        RECT 21.655 28.830 21.825 29.495 ;
        RECT 21.995 29.075 22.165 29.835 ;
        RECT 22.400 29.075 22.915 29.485 ;
        RECT 21.655 28.640 22.405 28.830 ;
        RECT 22.575 28.265 22.915 29.075 ;
        RECT 23.145 28.695 23.355 29.835 ;
        RECT 21.685 28.095 22.915 28.265 ;
        RECT 23.525 28.685 23.855 29.665 ;
        RECT 24.025 28.695 24.255 29.835 ;
        RECT 24.465 28.745 27.975 29.835 ;
        RECT 28.145 28.745 29.355 29.835 ;
        RECT 29.615 29.090 29.885 29.835 ;
        RECT 30.515 29.830 36.790 29.835 ;
        RECT 30.055 28.920 30.345 29.660 ;
        RECT 30.515 29.105 30.770 29.830 ;
        RECT 30.955 28.935 31.215 29.660 ;
        RECT 31.385 29.105 31.630 29.830 ;
        RECT 31.815 28.935 32.075 29.660 ;
        RECT 32.245 29.105 32.490 29.830 ;
        RECT 32.675 28.935 32.935 29.660 ;
        RECT 33.105 29.105 33.350 29.830 ;
        RECT 33.520 28.935 33.780 29.660 ;
        RECT 33.950 29.105 34.210 29.830 ;
        RECT 34.380 28.935 34.640 29.660 ;
        RECT 34.810 29.105 35.070 29.830 ;
        RECT 35.240 28.935 35.500 29.660 ;
        RECT 35.670 29.105 35.930 29.830 ;
        RECT 36.100 28.935 36.360 29.660 ;
        RECT 36.530 29.035 36.790 29.830 ;
        RECT 30.955 28.920 36.360 28.935 ;
        RECT 21.665 27.285 22.175 27.820 ;
        RECT 22.395 27.490 22.640 28.095 ;
        RECT 23.145 27.285 23.355 28.105 ;
        RECT 23.525 28.085 23.775 28.685 ;
        RECT 23.945 28.275 24.275 28.525 ;
        RECT 23.525 27.455 23.855 28.085 ;
        RECT 24.025 27.285 24.255 28.105 ;
        RECT 24.465 28.055 26.115 28.575 ;
        RECT 26.285 28.225 27.975 28.745 ;
        RECT 24.465 27.285 27.975 28.055 ;
        RECT 28.145 28.035 28.665 28.575 ;
        RECT 28.835 28.205 29.355 28.745 ;
        RECT 29.615 28.695 36.360 28.920 ;
        RECT 29.615 28.135 30.780 28.695 ;
        RECT 36.960 28.525 37.210 29.660 ;
        RECT 37.390 29.025 37.650 29.835 ;
        RECT 37.825 28.525 38.070 29.665 ;
        RECT 38.250 29.025 38.545 29.835 ;
        RECT 38.785 28.695 38.995 29.835 ;
        RECT 39.165 28.685 39.495 29.665 ;
        RECT 39.665 28.695 39.895 29.835 ;
        RECT 40.105 28.745 42.695 29.835 ;
        RECT 30.950 28.275 38.070 28.525 ;
        RECT 29.585 28.105 30.780 28.135 ;
        RECT 28.145 27.285 29.355 28.035 ;
        RECT 29.585 27.965 36.360 28.105 ;
        RECT 29.615 27.935 36.360 27.965 ;
        RECT 29.615 27.285 29.915 27.765 ;
        RECT 30.085 27.480 30.345 27.935 ;
        RECT 30.515 27.285 30.775 27.765 ;
        RECT 30.955 27.480 31.215 27.935 ;
        RECT 31.385 27.285 31.635 27.765 ;
        RECT 31.815 27.480 32.075 27.935 ;
        RECT 32.245 27.285 32.495 27.765 ;
        RECT 32.675 27.480 32.935 27.935 ;
        RECT 33.105 27.285 33.350 27.765 ;
        RECT 33.520 27.480 33.795 27.935 ;
        RECT 33.965 27.285 34.210 27.765 ;
        RECT 34.380 27.480 34.640 27.935 ;
        RECT 34.810 27.285 35.070 27.765 ;
        RECT 35.240 27.480 35.500 27.935 ;
        RECT 35.670 27.285 35.930 27.765 ;
        RECT 36.100 27.480 36.360 27.935 ;
        RECT 36.530 27.285 36.790 27.845 ;
        RECT 36.960 27.465 37.210 28.275 ;
        RECT 37.390 27.285 37.650 27.810 ;
        RECT 37.820 27.465 38.070 28.275 ;
        RECT 38.240 27.965 38.555 28.525 ;
        RECT 38.250 27.285 38.555 27.795 ;
        RECT 38.785 27.285 38.995 28.105 ;
        RECT 39.165 28.085 39.415 28.685 ;
        RECT 39.585 28.275 39.915 28.525 ;
        RECT 39.165 27.455 39.495 28.085 ;
        RECT 39.665 27.285 39.895 28.105 ;
        RECT 40.105 28.055 41.315 28.575 ;
        RECT 41.485 28.225 42.695 28.745 ;
        RECT 42.905 28.695 43.135 29.835 ;
        RECT 43.305 28.685 43.635 29.665 ;
        RECT 43.805 28.695 44.015 29.835 ;
        RECT 42.885 28.275 43.215 28.525 ;
        RECT 40.105 27.285 42.695 28.055 ;
        RECT 42.905 27.285 43.135 28.105 ;
        RECT 43.385 28.085 43.635 28.685 ;
        RECT 44.245 28.670 44.535 29.835 ;
        RECT 44.710 28.695 45.045 29.665 ;
        RECT 45.215 28.695 45.385 29.835 ;
        RECT 45.555 29.495 47.585 29.665 ;
        RECT 43.305 27.455 43.635 28.085 ;
        RECT 43.805 27.285 44.015 28.105 ;
        RECT 44.710 28.025 44.880 28.695 ;
        RECT 45.555 28.525 45.725 29.495 ;
        RECT 45.050 28.195 45.305 28.525 ;
        RECT 45.530 28.195 45.725 28.525 ;
        RECT 45.895 29.155 47.020 29.325 ;
        RECT 45.135 28.025 45.305 28.195 ;
        RECT 45.895 28.025 46.065 29.155 ;
        RECT 44.245 27.285 44.535 28.010 ;
        RECT 44.710 27.455 44.965 28.025 ;
        RECT 45.135 27.855 46.065 28.025 ;
        RECT 46.235 28.815 47.245 28.985 ;
        RECT 46.235 28.015 46.405 28.815 ;
        RECT 46.610 28.475 46.885 28.615 ;
        RECT 46.605 28.305 46.885 28.475 ;
        RECT 45.890 27.820 46.065 27.855 ;
        RECT 45.135 27.285 45.465 27.685 ;
        RECT 45.890 27.455 46.420 27.820 ;
        RECT 46.610 27.455 46.885 28.305 ;
        RECT 47.055 27.455 47.245 28.815 ;
        RECT 47.415 28.830 47.585 29.495 ;
        RECT 47.755 29.075 47.925 29.835 ;
        RECT 48.160 29.075 48.675 29.485 ;
        RECT 48.845 29.400 54.190 29.835 ;
        RECT 47.415 28.640 48.165 28.830 ;
        RECT 48.335 28.265 48.675 29.075 ;
        RECT 47.445 28.095 48.675 28.265 ;
        RECT 47.425 27.285 47.935 27.820 ;
        RECT 48.155 27.490 48.400 28.095 ;
        RECT 50.430 27.830 50.770 28.660 ;
        RECT 52.250 28.150 52.600 29.400 ;
        RECT 54.365 28.745 57.875 29.835 ;
        RECT 54.365 28.055 56.015 28.575 ;
        RECT 56.185 28.225 57.875 28.745 ;
        RECT 58.045 28.695 58.305 29.835 ;
        RECT 58.545 29.325 60.160 29.655 ;
        RECT 58.555 28.525 58.725 29.085 ;
        RECT 58.985 28.985 60.160 29.155 ;
        RECT 60.330 29.035 60.610 29.835 ;
        RECT 58.985 28.695 59.315 28.985 ;
        RECT 59.990 28.865 60.160 28.985 ;
        RECT 59.485 28.525 59.730 28.815 ;
        RECT 59.990 28.695 60.650 28.865 ;
        RECT 60.820 28.695 61.095 29.665 ;
        RECT 60.480 28.525 60.650 28.695 ;
        RECT 58.050 28.275 58.385 28.525 ;
        RECT 58.555 28.195 59.270 28.525 ;
        RECT 59.485 28.195 60.310 28.525 ;
        RECT 60.480 28.195 60.755 28.525 ;
        RECT 58.555 28.105 58.805 28.195 ;
        RECT 48.845 27.285 54.190 27.830 ;
        RECT 54.365 27.285 57.875 28.055 ;
        RECT 58.045 27.285 58.305 28.105 ;
        RECT 58.475 27.685 58.805 28.105 ;
        RECT 60.480 28.025 60.650 28.195 ;
        RECT 58.985 27.855 60.650 28.025 ;
        RECT 60.925 27.960 61.095 28.695 ;
        RECT 58.985 27.455 59.245 27.855 ;
        RECT 59.415 27.285 59.745 27.685 ;
        RECT 59.915 27.505 60.085 27.855 ;
        RECT 60.255 27.285 60.630 27.685 ;
        RECT 60.820 27.615 61.095 27.960 ;
        RECT 61.265 28.695 61.540 29.665 ;
        RECT 61.750 29.035 62.030 29.835 ;
        RECT 62.200 29.325 63.815 29.655 ;
        RECT 62.200 28.985 63.375 29.155 ;
        RECT 62.200 28.865 62.370 28.985 ;
        RECT 61.710 28.695 62.370 28.865 ;
        RECT 61.265 27.960 61.435 28.695 ;
        RECT 61.710 28.525 61.880 28.695 ;
        RECT 62.630 28.525 62.875 28.815 ;
        RECT 63.045 28.695 63.375 28.985 ;
        RECT 63.635 28.525 63.805 29.085 ;
        RECT 64.055 28.695 64.315 29.835 ;
        RECT 64.485 28.745 66.155 29.835 ;
        RECT 61.605 28.195 61.880 28.525 ;
        RECT 62.050 28.195 62.875 28.525 ;
        RECT 63.090 28.195 63.805 28.525 ;
        RECT 63.975 28.275 64.310 28.525 ;
        RECT 61.710 28.025 61.880 28.195 ;
        RECT 63.555 28.105 63.805 28.195 ;
        RECT 61.265 27.615 61.540 27.960 ;
        RECT 61.710 27.855 63.375 28.025 ;
        RECT 61.730 27.285 62.105 27.685 ;
        RECT 62.275 27.505 62.445 27.855 ;
        RECT 62.615 27.285 62.945 27.685 ;
        RECT 63.115 27.455 63.375 27.855 ;
        RECT 63.555 27.685 63.885 28.105 ;
        RECT 64.055 27.285 64.315 28.105 ;
        RECT 64.485 28.055 65.235 28.575 ;
        RECT 65.405 28.225 66.155 28.745 ;
        RECT 66.825 28.695 67.055 29.835 ;
        RECT 67.225 28.685 67.555 29.665 ;
        RECT 67.725 28.695 67.935 29.835 ;
        RECT 68.165 28.745 69.835 29.835 ;
        RECT 66.805 28.275 67.135 28.525 ;
        RECT 64.485 27.285 66.155 28.055 ;
        RECT 66.825 27.285 67.055 28.105 ;
        RECT 67.305 28.085 67.555 28.685 ;
        RECT 67.225 27.455 67.555 28.085 ;
        RECT 67.725 27.285 67.935 28.105 ;
        RECT 68.165 28.055 68.915 28.575 ;
        RECT 69.085 28.225 69.835 28.745 ;
        RECT 70.005 28.670 70.295 29.835 ;
        RECT 70.465 28.745 73.975 29.835 ;
        RECT 70.465 28.055 72.115 28.575 ;
        RECT 72.285 28.225 73.975 28.745 ;
        RECT 75.070 28.645 75.325 29.525 ;
        RECT 75.495 28.695 75.800 29.835 ;
        RECT 76.140 29.455 76.470 29.835 ;
        RECT 76.650 29.285 76.820 29.575 ;
        RECT 76.990 29.375 77.240 29.835 ;
        RECT 76.020 29.115 76.820 29.285 ;
        RECT 77.410 29.325 78.280 29.665 ;
        RECT 68.165 27.285 69.835 28.055 ;
        RECT 70.005 27.285 70.295 28.010 ;
        RECT 70.465 27.285 73.975 28.055 ;
        RECT 75.070 27.995 75.280 28.645 ;
        RECT 76.020 28.525 76.190 29.115 ;
        RECT 77.410 28.945 77.580 29.325 ;
        RECT 78.515 29.205 78.685 29.665 ;
        RECT 78.855 29.375 79.225 29.835 ;
        RECT 79.520 29.235 79.690 29.575 ;
        RECT 79.860 29.405 80.190 29.835 ;
        RECT 80.425 29.235 80.595 29.575 ;
        RECT 76.360 28.775 77.580 28.945 ;
        RECT 77.750 28.865 78.210 29.155 ;
        RECT 78.515 29.035 79.075 29.205 ;
        RECT 79.520 29.065 80.595 29.235 ;
        RECT 80.765 29.335 81.445 29.665 ;
        RECT 81.660 29.335 81.910 29.665 ;
        RECT 82.080 29.375 82.330 29.835 ;
        RECT 78.905 28.895 79.075 29.035 ;
        RECT 77.750 28.855 78.715 28.865 ;
        RECT 77.410 28.685 77.580 28.775 ;
        RECT 78.040 28.695 78.715 28.855 ;
        RECT 75.450 28.495 76.190 28.525 ;
        RECT 75.450 28.195 76.365 28.495 ;
        RECT 76.040 28.020 76.365 28.195 ;
        RECT 75.070 27.465 75.325 27.995 ;
        RECT 75.495 27.285 75.800 27.745 ;
        RECT 76.045 27.665 76.365 28.020 ;
        RECT 76.535 28.235 77.075 28.605 ;
        RECT 77.410 28.515 77.815 28.685 ;
        RECT 76.535 27.835 76.775 28.235 ;
        RECT 77.255 28.065 77.475 28.345 ;
        RECT 76.945 27.895 77.475 28.065 ;
        RECT 76.945 27.665 77.115 27.895 ;
        RECT 77.645 27.735 77.815 28.515 ;
        RECT 77.985 27.905 78.335 28.525 ;
        RECT 78.505 27.905 78.715 28.695 ;
        RECT 78.905 28.725 80.405 28.895 ;
        RECT 78.905 28.035 79.075 28.725 ;
        RECT 80.765 28.555 80.935 29.335 ;
        RECT 81.740 29.205 81.910 29.335 ;
        RECT 79.245 28.385 80.935 28.555 ;
        RECT 81.105 28.775 81.570 29.165 ;
        RECT 81.740 29.035 82.135 29.205 ;
        RECT 79.245 28.205 79.415 28.385 ;
        RECT 76.045 27.495 77.115 27.665 ;
        RECT 77.285 27.285 77.475 27.725 ;
        RECT 77.645 27.455 78.595 27.735 ;
        RECT 78.905 27.645 79.165 28.035 ;
        RECT 79.585 27.965 80.375 28.215 ;
        RECT 78.815 27.475 79.165 27.645 ;
        RECT 79.375 27.285 79.705 27.745 ;
        RECT 80.580 27.675 80.750 28.385 ;
        RECT 81.105 28.185 81.275 28.775 ;
        RECT 80.920 27.965 81.275 28.185 ;
        RECT 81.445 27.965 81.795 28.585 ;
        RECT 81.965 27.675 82.135 29.035 ;
        RECT 82.500 28.865 82.825 29.650 ;
        RECT 82.305 27.815 82.765 28.865 ;
        RECT 80.580 27.505 81.435 27.675 ;
        RECT 81.640 27.505 82.135 27.675 ;
        RECT 82.305 27.285 82.635 27.645 ;
        RECT 82.995 27.545 83.165 29.665 ;
        RECT 83.335 29.335 83.665 29.835 ;
        RECT 83.835 29.165 84.090 29.665 ;
        RECT 83.340 28.995 84.090 29.165 ;
        RECT 83.340 28.005 83.570 28.995 ;
        RECT 83.740 28.175 84.090 28.825 ;
        RECT 84.305 28.695 84.535 29.835 ;
        RECT 84.705 28.685 85.035 29.665 ;
        RECT 85.205 28.695 85.415 29.835 ;
        RECT 85.645 29.400 90.990 29.835 ;
        RECT 84.285 28.275 84.615 28.525 ;
        RECT 83.340 27.835 84.090 28.005 ;
        RECT 83.335 27.285 83.665 27.665 ;
        RECT 83.835 27.545 84.090 27.835 ;
        RECT 84.305 27.285 84.535 28.105 ;
        RECT 84.785 28.085 85.035 28.685 ;
        RECT 84.705 27.455 85.035 28.085 ;
        RECT 85.205 27.285 85.415 28.105 ;
        RECT 87.230 27.830 87.570 28.660 ;
        RECT 89.050 28.150 89.400 29.400 ;
        RECT 91.165 28.745 94.675 29.835 ;
        RECT 91.165 28.055 92.815 28.575 ;
        RECT 92.985 28.225 94.675 28.745 ;
        RECT 95.765 28.670 96.055 29.835 ;
        RECT 96.225 29.400 101.570 29.835 ;
        RECT 101.745 29.400 107.090 29.835 ;
        RECT 107.265 29.400 112.610 29.835 ;
        RECT 85.645 27.285 90.990 27.830 ;
        RECT 91.165 27.285 94.675 28.055 ;
        RECT 95.765 27.285 96.055 28.010 ;
        RECT 97.810 27.830 98.150 28.660 ;
        RECT 99.630 28.150 99.980 29.400 ;
        RECT 103.330 27.830 103.670 28.660 ;
        RECT 105.150 28.150 105.500 29.400 ;
        RECT 108.850 27.830 109.190 28.660 ;
        RECT 110.670 28.150 111.020 29.400 ;
        RECT 112.785 28.745 116.295 29.835 ;
        RECT 112.785 28.055 114.435 28.575 ;
        RECT 114.605 28.225 116.295 28.745 ;
        RECT 117.385 28.745 118.595 29.835 ;
        RECT 117.385 28.205 117.905 28.745 ;
        RECT 96.225 27.285 101.570 27.830 ;
        RECT 101.745 27.285 107.090 27.830 ;
        RECT 107.265 27.285 112.610 27.830 ;
        RECT 112.785 27.285 116.295 28.055 ;
        RECT 118.075 28.035 118.595 28.575 ;
        RECT 117.385 27.285 118.595 28.035 ;
        RECT 5.520 27.115 118.680 27.285 ;
        RECT 5.605 26.365 6.815 27.115 ;
        RECT 6.985 26.570 12.330 27.115 ;
        RECT 5.605 25.825 6.125 26.365 ;
        RECT 6.295 25.655 6.815 26.195 ;
        RECT 8.570 25.740 8.910 26.570 ;
        RECT 12.505 26.365 13.715 27.115 ;
        RECT 13.890 26.565 14.145 26.855 ;
        RECT 14.315 26.735 14.645 27.115 ;
        RECT 13.890 26.395 14.640 26.565 ;
        RECT 5.605 24.565 6.815 25.655 ;
        RECT 10.390 25.000 10.740 26.250 ;
        RECT 12.505 25.825 13.025 26.365 ;
        RECT 13.195 25.655 13.715 26.195 ;
        RECT 6.985 24.565 12.330 25.000 ;
        RECT 12.505 24.565 13.715 25.655 ;
        RECT 13.890 25.575 14.240 26.225 ;
        RECT 14.410 25.405 14.640 26.395 ;
        RECT 13.890 25.235 14.640 25.405 ;
        RECT 13.890 24.735 14.145 25.235 ;
        RECT 14.315 24.565 14.645 25.065 ;
        RECT 14.815 24.735 14.985 26.855 ;
        RECT 15.345 26.755 15.675 27.115 ;
        RECT 15.845 26.725 16.340 26.895 ;
        RECT 16.545 26.725 17.400 26.895 ;
        RECT 15.215 25.535 15.675 26.585 ;
        RECT 15.155 24.750 15.480 25.535 ;
        RECT 15.845 25.365 16.015 26.725 ;
        RECT 16.185 25.815 16.535 26.435 ;
        RECT 16.705 26.215 17.060 26.435 ;
        RECT 16.705 25.625 16.875 26.215 ;
        RECT 17.230 26.015 17.400 26.725 ;
        RECT 18.275 26.655 18.605 27.115 ;
        RECT 18.815 26.755 19.165 26.925 ;
        RECT 17.605 26.185 18.395 26.435 ;
        RECT 18.815 26.365 19.075 26.755 ;
        RECT 19.385 26.665 20.335 26.945 ;
        RECT 20.505 26.675 20.695 27.115 ;
        RECT 20.865 26.735 21.935 26.905 ;
        RECT 18.565 26.015 18.735 26.195 ;
        RECT 15.845 25.195 16.240 25.365 ;
        RECT 16.410 25.235 16.875 25.625 ;
        RECT 17.045 25.845 18.735 26.015 ;
        RECT 16.070 25.065 16.240 25.195 ;
        RECT 17.045 25.065 17.215 25.845 ;
        RECT 18.905 25.675 19.075 26.365 ;
        RECT 17.575 25.505 19.075 25.675 ;
        RECT 19.265 25.705 19.475 26.495 ;
        RECT 19.645 25.875 19.995 26.495 ;
        RECT 20.165 25.885 20.335 26.665 ;
        RECT 20.865 26.505 21.035 26.735 ;
        RECT 20.505 26.335 21.035 26.505 ;
        RECT 20.505 26.055 20.725 26.335 ;
        RECT 21.205 26.165 21.445 26.565 ;
        RECT 20.165 25.715 20.570 25.885 ;
        RECT 20.905 25.795 21.445 26.165 ;
        RECT 21.615 26.380 21.935 26.735 ;
        RECT 22.180 26.655 22.485 27.115 ;
        RECT 22.655 26.405 22.910 26.935 ;
        RECT 23.085 26.570 28.430 27.115 ;
        RECT 21.615 26.205 21.940 26.380 ;
        RECT 21.615 25.905 22.530 26.205 ;
        RECT 21.790 25.875 22.530 25.905 ;
        RECT 19.265 25.545 19.940 25.705 ;
        RECT 20.400 25.625 20.570 25.715 ;
        RECT 19.265 25.535 20.230 25.545 ;
        RECT 18.905 25.365 19.075 25.505 ;
        RECT 15.650 24.565 15.900 25.025 ;
        RECT 16.070 24.735 16.320 25.065 ;
        RECT 16.535 24.735 17.215 25.065 ;
        RECT 17.385 25.165 18.460 25.335 ;
        RECT 18.905 25.195 19.465 25.365 ;
        RECT 19.770 25.245 20.230 25.535 ;
        RECT 20.400 25.455 21.620 25.625 ;
        RECT 17.385 24.825 17.555 25.165 ;
        RECT 17.790 24.565 18.120 24.995 ;
        RECT 18.290 24.825 18.460 25.165 ;
        RECT 18.755 24.565 19.125 25.025 ;
        RECT 19.295 24.735 19.465 25.195 ;
        RECT 20.400 25.075 20.570 25.455 ;
        RECT 21.790 25.285 21.960 25.875 ;
        RECT 22.700 25.755 22.910 26.405 ;
        RECT 19.700 24.735 20.570 25.075 ;
        RECT 21.160 25.115 21.960 25.285 ;
        RECT 20.740 24.565 20.990 25.025 ;
        RECT 21.160 24.825 21.330 25.115 ;
        RECT 21.510 24.565 21.840 24.945 ;
        RECT 22.180 24.565 22.485 25.705 ;
        RECT 22.655 24.875 22.910 25.755 ;
        RECT 24.670 25.740 25.010 26.570 ;
        RECT 28.605 26.345 31.195 27.115 ;
        RECT 31.365 26.390 31.655 27.115 ;
        RECT 31.825 26.375 32.210 26.945 ;
        RECT 32.380 26.655 32.705 27.115 ;
        RECT 33.225 26.485 33.505 26.945 ;
        RECT 26.490 25.000 26.840 26.250 ;
        RECT 28.605 25.825 29.815 26.345 ;
        RECT 29.985 25.655 31.195 26.175 ;
        RECT 23.085 24.565 28.430 25.000 ;
        RECT 28.605 24.565 31.195 25.655 ;
        RECT 31.365 24.565 31.655 25.730 ;
        RECT 31.825 25.705 32.105 26.375 ;
        RECT 32.380 26.315 33.505 26.485 ;
        RECT 32.380 26.205 32.830 26.315 ;
        RECT 32.275 25.875 32.830 26.205 ;
        RECT 33.695 26.145 34.095 26.945 ;
        RECT 34.495 26.655 34.765 27.115 ;
        RECT 34.935 26.485 35.220 26.945 ;
        RECT 31.825 24.735 32.210 25.705 ;
        RECT 32.380 25.415 32.830 25.875 ;
        RECT 33.000 25.585 34.095 26.145 ;
        RECT 32.380 25.195 33.505 25.415 ;
        RECT 32.380 24.565 32.705 25.025 ;
        RECT 33.225 24.735 33.505 25.195 ;
        RECT 33.695 24.735 34.095 25.585 ;
        RECT 34.265 26.315 35.220 26.485 ;
        RECT 35.505 26.345 38.095 27.115 ;
        RECT 38.355 26.565 38.525 26.855 ;
        RECT 38.695 26.735 39.025 27.115 ;
        RECT 38.355 26.395 39.020 26.565 ;
        RECT 34.265 25.415 34.475 26.315 ;
        RECT 34.645 25.585 35.335 26.145 ;
        RECT 35.505 25.825 36.715 26.345 ;
        RECT 36.885 25.655 38.095 26.175 ;
        RECT 34.265 25.195 35.220 25.415 ;
        RECT 34.495 24.565 34.765 25.025 ;
        RECT 34.935 24.735 35.220 25.195 ;
        RECT 35.505 24.565 38.095 25.655 ;
        RECT 38.270 25.575 38.620 26.225 ;
        RECT 38.790 25.405 39.020 26.395 ;
        RECT 38.355 25.235 39.020 25.405 ;
        RECT 38.355 24.735 38.525 25.235 ;
        RECT 38.695 24.565 39.025 25.065 ;
        RECT 39.195 24.735 39.420 26.855 ;
        RECT 39.635 26.735 39.965 27.115 ;
        RECT 40.135 26.565 40.305 26.895 ;
        RECT 40.605 26.735 41.620 26.935 ;
        RECT 39.610 26.375 40.305 26.565 ;
        RECT 39.610 25.405 39.780 26.375 ;
        RECT 39.950 25.575 40.360 26.195 ;
        RECT 40.530 25.625 40.750 26.495 ;
        RECT 40.930 26.185 41.280 26.555 ;
        RECT 41.450 26.005 41.620 26.735 ;
        RECT 41.790 26.675 42.200 27.115 ;
        RECT 42.490 26.475 42.740 26.905 ;
        RECT 42.940 26.655 43.260 27.115 ;
        RECT 43.820 26.725 44.670 26.895 ;
        RECT 41.790 26.135 42.200 26.465 ;
        RECT 42.490 26.135 42.910 26.475 ;
        RECT 41.200 25.965 41.620 26.005 ;
        RECT 41.200 25.795 42.550 25.965 ;
        RECT 39.610 25.235 40.305 25.405 ;
        RECT 40.530 25.245 41.030 25.625 ;
        RECT 39.635 24.565 39.965 25.065 ;
        RECT 40.135 24.735 40.305 25.235 ;
        RECT 41.200 24.950 41.370 25.795 ;
        RECT 42.300 25.635 42.550 25.795 ;
        RECT 41.540 25.365 41.790 25.625 ;
        RECT 42.720 25.365 42.910 26.135 ;
        RECT 41.540 25.115 42.910 25.365 ;
        RECT 43.080 26.305 44.330 26.475 ;
        RECT 43.080 25.545 43.250 26.305 ;
        RECT 44.000 26.185 44.330 26.305 ;
        RECT 43.420 25.725 43.600 26.135 ;
        RECT 44.500 25.965 44.670 26.725 ;
        RECT 44.870 26.635 45.530 27.115 ;
        RECT 45.710 26.520 46.030 26.850 ;
        RECT 44.860 26.195 45.520 26.465 ;
        RECT 44.860 26.135 45.190 26.195 ;
        RECT 45.340 25.965 45.670 26.025 ;
        RECT 43.770 25.795 45.670 25.965 ;
        RECT 43.080 25.235 43.600 25.545 ;
        RECT 43.770 25.285 43.940 25.795 ;
        RECT 45.840 25.625 46.030 26.520 ;
        RECT 44.110 25.455 46.030 25.625 ;
        RECT 45.710 25.435 46.030 25.455 ;
        RECT 46.230 26.205 46.480 26.855 ;
        RECT 46.660 26.655 46.945 27.115 ;
        RECT 47.125 26.775 47.380 26.935 ;
        RECT 47.125 26.605 47.465 26.775 ;
        RECT 47.125 26.405 47.380 26.605 ;
        RECT 47.925 26.570 53.270 27.115 ;
        RECT 46.230 25.875 47.030 26.205 ;
        RECT 43.770 25.115 44.980 25.285 ;
        RECT 40.540 24.780 41.370 24.950 ;
        RECT 41.610 24.565 41.990 24.945 ;
        RECT 42.170 24.825 42.340 25.115 ;
        RECT 43.770 25.035 43.940 25.115 ;
        RECT 42.510 24.565 42.840 24.945 ;
        RECT 43.310 24.785 43.940 25.035 ;
        RECT 44.120 24.565 44.540 24.945 ;
        RECT 44.740 24.825 44.980 25.115 ;
        RECT 45.210 24.565 45.540 25.255 ;
        RECT 45.710 24.825 45.880 25.435 ;
        RECT 46.230 25.285 46.480 25.875 ;
        RECT 47.200 25.545 47.380 26.405 ;
        RECT 49.510 25.740 49.850 26.570 ;
        RECT 53.445 26.345 56.955 27.115 ;
        RECT 57.125 26.390 57.415 27.115 ;
        RECT 57.585 26.365 58.795 27.115 ;
        RECT 59.295 26.715 59.625 27.115 ;
        RECT 59.795 26.545 60.125 26.885 ;
        RECT 61.175 26.715 61.505 27.115 ;
        RECT 59.140 26.375 61.505 26.545 ;
        RECT 61.675 26.390 62.005 26.900 ;
        RECT 62.185 26.735 63.075 26.905 ;
        RECT 46.150 24.775 46.480 25.285 ;
        RECT 46.660 24.565 46.945 25.365 ;
        RECT 47.125 24.875 47.380 25.545 ;
        RECT 51.330 25.000 51.680 26.250 ;
        RECT 53.445 25.825 55.095 26.345 ;
        RECT 55.265 25.655 56.955 26.175 ;
        RECT 57.585 25.825 58.105 26.365 ;
        RECT 47.925 24.565 53.270 25.000 ;
        RECT 53.445 24.565 56.955 25.655 ;
        RECT 57.125 24.565 57.415 25.730 ;
        RECT 58.275 25.655 58.795 26.195 ;
        RECT 57.585 24.565 58.795 25.655 ;
        RECT 59.140 25.375 59.310 26.375 ;
        RECT 61.335 26.205 61.505 26.375 ;
        RECT 59.480 25.545 59.725 26.205 ;
        RECT 59.940 25.545 60.205 26.205 ;
        RECT 60.400 25.545 60.685 26.205 ;
        RECT 60.860 25.875 61.165 26.205 ;
        RECT 61.335 25.875 61.645 26.205 ;
        RECT 60.860 25.545 61.075 25.875 ;
        RECT 59.140 25.205 59.595 25.375 ;
        RECT 59.265 24.775 59.595 25.205 ;
        RECT 59.775 25.205 61.065 25.375 ;
        RECT 59.775 24.785 60.025 25.205 ;
        RECT 60.255 24.565 60.585 25.035 ;
        RECT 60.815 24.785 61.065 25.205 ;
        RECT 61.255 24.565 61.505 25.705 ;
        RECT 61.815 25.625 62.005 26.390 ;
        RECT 62.185 26.180 62.735 26.565 ;
        RECT 62.905 26.010 63.075 26.735 ;
        RECT 61.675 24.775 62.005 25.625 ;
        RECT 62.185 25.940 63.075 26.010 ;
        RECT 63.245 26.410 63.465 26.895 ;
        RECT 63.635 26.575 63.885 27.115 ;
        RECT 64.055 26.465 64.315 26.945 ;
        RECT 64.485 26.570 69.830 27.115 ;
        RECT 70.005 26.570 75.350 27.115 ;
        RECT 63.245 25.985 63.575 26.410 ;
        RECT 62.185 25.915 63.080 25.940 ;
        RECT 62.185 25.900 63.090 25.915 ;
        RECT 62.185 25.885 63.095 25.900 ;
        RECT 62.185 25.880 63.105 25.885 ;
        RECT 62.185 25.870 63.110 25.880 ;
        RECT 62.185 25.860 63.115 25.870 ;
        RECT 62.185 25.855 63.125 25.860 ;
        RECT 62.185 25.845 63.135 25.855 ;
        RECT 62.185 25.840 63.145 25.845 ;
        RECT 62.185 25.390 62.445 25.840 ;
        RECT 62.810 25.835 63.145 25.840 ;
        RECT 62.810 25.830 63.160 25.835 ;
        RECT 62.810 25.820 63.175 25.830 ;
        RECT 62.810 25.815 63.200 25.820 ;
        RECT 63.745 25.815 63.975 26.210 ;
        RECT 62.810 25.810 63.975 25.815 ;
        RECT 62.840 25.775 63.975 25.810 ;
        RECT 62.875 25.750 63.975 25.775 ;
        RECT 62.905 25.720 63.975 25.750 ;
        RECT 62.925 25.690 63.975 25.720 ;
        RECT 62.945 25.660 63.975 25.690 ;
        RECT 63.015 25.650 63.975 25.660 ;
        RECT 63.040 25.640 63.975 25.650 ;
        RECT 63.060 25.625 63.975 25.640 ;
        RECT 63.080 25.610 63.975 25.625 ;
        RECT 63.085 25.600 63.870 25.610 ;
        RECT 63.100 25.565 63.870 25.600 ;
        RECT 62.615 25.245 62.945 25.490 ;
        RECT 63.115 25.315 63.870 25.565 ;
        RECT 64.145 25.435 64.315 26.465 ;
        RECT 66.070 25.740 66.410 26.570 ;
        RECT 62.615 25.220 62.800 25.245 ;
        RECT 62.185 25.120 62.800 25.220 ;
        RECT 62.185 24.565 62.790 25.120 ;
        RECT 62.965 24.735 63.445 25.075 ;
        RECT 63.615 24.565 63.870 25.110 ;
        RECT 64.040 24.735 64.315 25.435 ;
        RECT 67.890 25.000 68.240 26.250 ;
        RECT 71.590 25.740 71.930 26.570 ;
        RECT 75.525 26.375 75.910 26.945 ;
        RECT 76.080 26.655 76.405 27.115 ;
        RECT 76.925 26.485 77.205 26.945 ;
        RECT 73.410 25.000 73.760 26.250 ;
        RECT 75.525 25.705 75.805 26.375 ;
        RECT 76.080 26.315 77.205 26.485 ;
        RECT 76.080 26.205 76.530 26.315 ;
        RECT 75.975 25.875 76.530 26.205 ;
        RECT 77.395 26.145 77.795 26.945 ;
        RECT 78.195 26.655 78.465 27.115 ;
        RECT 78.635 26.485 78.920 26.945 ;
        RECT 64.485 24.565 69.830 25.000 ;
        RECT 70.005 24.565 75.350 25.000 ;
        RECT 75.525 24.735 75.910 25.705 ;
        RECT 76.080 25.415 76.530 25.875 ;
        RECT 76.700 25.585 77.795 26.145 ;
        RECT 76.080 25.195 77.205 25.415 ;
        RECT 76.080 24.565 76.405 25.025 ;
        RECT 76.925 24.735 77.205 25.195 ;
        RECT 77.395 24.735 77.795 25.585 ;
        RECT 77.965 26.315 78.920 26.485 ;
        RECT 77.965 25.415 78.175 26.315 ;
        RECT 79.245 26.295 79.475 27.115 ;
        RECT 79.645 26.315 79.975 26.945 ;
        RECT 78.345 25.585 79.035 26.145 ;
        RECT 79.225 25.875 79.555 26.125 ;
        RECT 79.725 25.715 79.975 26.315 ;
        RECT 80.145 26.295 80.355 27.115 ;
        RECT 80.585 26.345 82.255 27.115 ;
        RECT 82.885 26.390 83.175 27.115 ;
        RECT 83.345 26.570 88.690 27.115 ;
        RECT 88.865 26.570 94.210 27.115 ;
        RECT 94.385 26.570 99.730 27.115 ;
        RECT 99.905 26.570 105.250 27.115 ;
        RECT 80.585 25.825 81.335 26.345 ;
        RECT 77.965 25.195 78.920 25.415 ;
        RECT 78.195 24.565 78.465 25.025 ;
        RECT 78.635 24.735 78.920 25.195 ;
        RECT 79.245 24.565 79.475 25.705 ;
        RECT 79.645 24.735 79.975 25.715 ;
        RECT 80.145 24.565 80.355 25.705 ;
        RECT 81.505 25.655 82.255 26.175 ;
        RECT 84.930 25.740 85.270 26.570 ;
        RECT 80.585 24.565 82.255 25.655 ;
        RECT 82.885 24.565 83.175 25.730 ;
        RECT 86.750 25.000 87.100 26.250 ;
        RECT 90.450 25.740 90.790 26.570 ;
        RECT 92.270 25.000 92.620 26.250 ;
        RECT 95.970 25.740 96.310 26.570 ;
        RECT 97.790 25.000 98.140 26.250 ;
        RECT 101.490 25.740 101.830 26.570 ;
        RECT 105.425 26.345 108.015 27.115 ;
        RECT 108.645 26.390 108.935 27.115 ;
        RECT 109.105 26.570 114.450 27.115 ;
        RECT 103.310 25.000 103.660 26.250 ;
        RECT 105.425 25.825 106.635 26.345 ;
        RECT 106.805 25.655 108.015 26.175 ;
        RECT 110.690 25.740 111.030 26.570 ;
        RECT 114.625 26.345 117.215 27.115 ;
        RECT 117.385 26.365 118.595 27.115 ;
        RECT 83.345 24.565 88.690 25.000 ;
        RECT 88.865 24.565 94.210 25.000 ;
        RECT 94.385 24.565 99.730 25.000 ;
        RECT 99.905 24.565 105.250 25.000 ;
        RECT 105.425 24.565 108.015 25.655 ;
        RECT 108.645 24.565 108.935 25.730 ;
        RECT 112.510 25.000 112.860 26.250 ;
        RECT 114.625 25.825 115.835 26.345 ;
        RECT 116.005 25.655 117.215 26.175 ;
        RECT 109.105 24.565 114.450 25.000 ;
        RECT 114.625 24.565 117.215 25.655 ;
        RECT 117.385 25.655 117.905 26.195 ;
        RECT 118.075 25.825 118.595 26.365 ;
        RECT 117.385 24.565 118.595 25.655 ;
        RECT 5.520 24.395 118.680 24.565 ;
        RECT 5.605 23.305 6.815 24.395 ;
        RECT 6.985 23.960 12.330 24.395 ;
        RECT 12.505 23.960 17.850 24.395 ;
        RECT 5.605 22.595 6.125 23.135 ;
        RECT 6.295 22.765 6.815 23.305 ;
        RECT 5.605 21.845 6.815 22.595 ;
        RECT 8.570 22.390 8.910 23.220 ;
        RECT 10.390 22.710 10.740 23.960 ;
        RECT 14.090 22.390 14.430 23.220 ;
        RECT 15.910 22.710 16.260 23.960 ;
        RECT 18.485 23.230 18.775 24.395 ;
        RECT 18.945 23.960 24.290 24.395 ;
        RECT 6.985 21.845 12.330 22.390 ;
        RECT 12.505 21.845 17.850 22.390 ;
        RECT 18.485 21.845 18.775 22.570 ;
        RECT 20.530 22.390 20.870 23.220 ;
        RECT 22.350 22.710 22.700 23.960 ;
        RECT 24.465 23.305 27.055 24.395 ;
        RECT 27.230 23.725 27.485 24.225 ;
        RECT 27.655 23.895 27.985 24.395 ;
        RECT 27.230 23.555 27.980 23.725 ;
        RECT 24.465 22.615 25.675 23.135 ;
        RECT 25.845 22.785 27.055 23.305 ;
        RECT 27.230 22.735 27.580 23.385 ;
        RECT 18.945 21.845 24.290 22.390 ;
        RECT 24.465 21.845 27.055 22.615 ;
        RECT 27.750 22.565 27.980 23.555 ;
        RECT 27.230 22.395 27.980 22.565 ;
        RECT 27.230 22.105 27.485 22.395 ;
        RECT 27.655 21.845 27.985 22.225 ;
        RECT 28.155 22.105 28.325 24.225 ;
        RECT 28.495 23.425 28.820 24.210 ;
        RECT 28.990 23.935 29.240 24.395 ;
        RECT 29.410 23.895 29.660 24.225 ;
        RECT 29.875 23.895 30.555 24.225 ;
        RECT 29.410 23.765 29.580 23.895 ;
        RECT 29.185 23.595 29.580 23.765 ;
        RECT 28.555 22.375 29.015 23.425 ;
        RECT 29.185 22.235 29.355 23.595 ;
        RECT 29.750 23.335 30.215 23.725 ;
        RECT 29.525 22.525 29.875 23.145 ;
        RECT 30.045 22.745 30.215 23.335 ;
        RECT 30.385 23.115 30.555 23.895 ;
        RECT 30.725 23.795 30.895 24.135 ;
        RECT 31.130 23.965 31.460 24.395 ;
        RECT 31.630 23.795 31.800 24.135 ;
        RECT 32.095 23.935 32.465 24.395 ;
        RECT 30.725 23.625 31.800 23.795 ;
        RECT 32.635 23.765 32.805 24.225 ;
        RECT 33.040 23.885 33.910 24.225 ;
        RECT 34.080 23.935 34.330 24.395 ;
        RECT 32.245 23.595 32.805 23.765 ;
        RECT 32.245 23.455 32.415 23.595 ;
        RECT 30.915 23.285 32.415 23.455 ;
        RECT 33.110 23.425 33.570 23.715 ;
        RECT 30.385 22.945 32.075 23.115 ;
        RECT 30.045 22.525 30.400 22.745 ;
        RECT 30.570 22.235 30.740 22.945 ;
        RECT 30.945 22.525 31.735 22.775 ;
        RECT 31.905 22.765 32.075 22.945 ;
        RECT 32.245 22.595 32.415 23.285 ;
        RECT 28.685 21.845 29.015 22.205 ;
        RECT 29.185 22.065 29.680 22.235 ;
        RECT 29.885 22.065 30.740 22.235 ;
        RECT 31.615 21.845 31.945 22.305 ;
        RECT 32.155 22.205 32.415 22.595 ;
        RECT 32.605 23.415 33.570 23.425 ;
        RECT 33.740 23.505 33.910 23.885 ;
        RECT 34.500 23.845 34.670 24.135 ;
        RECT 34.850 24.015 35.180 24.395 ;
        RECT 34.500 23.675 35.300 23.845 ;
        RECT 32.605 23.255 33.280 23.415 ;
        RECT 33.740 23.335 34.960 23.505 ;
        RECT 32.605 22.465 32.815 23.255 ;
        RECT 33.740 23.245 33.910 23.335 ;
        RECT 32.985 22.465 33.335 23.085 ;
        RECT 33.505 23.075 33.910 23.245 ;
        RECT 33.505 22.295 33.675 23.075 ;
        RECT 33.845 22.625 34.065 22.905 ;
        RECT 34.245 22.795 34.785 23.165 ;
        RECT 35.130 23.085 35.300 23.675 ;
        RECT 35.520 23.255 35.825 24.395 ;
        RECT 35.995 23.205 36.250 24.085 ;
        RECT 36.425 23.960 41.770 24.395 ;
        RECT 35.130 23.055 35.870 23.085 ;
        RECT 33.845 22.455 34.375 22.625 ;
        RECT 32.155 22.035 32.505 22.205 ;
        RECT 32.725 22.015 33.675 22.295 ;
        RECT 33.845 21.845 34.035 22.285 ;
        RECT 34.205 22.225 34.375 22.455 ;
        RECT 34.545 22.395 34.785 22.795 ;
        RECT 34.955 22.755 35.870 23.055 ;
        RECT 34.955 22.580 35.280 22.755 ;
        RECT 34.955 22.225 35.275 22.580 ;
        RECT 36.040 22.555 36.250 23.205 ;
        RECT 34.205 22.055 35.275 22.225 ;
        RECT 35.520 21.845 35.825 22.305 ;
        RECT 35.995 22.025 36.250 22.555 ;
        RECT 38.010 22.390 38.350 23.220 ;
        RECT 39.830 22.710 40.180 23.960 ;
        RECT 41.945 23.305 43.615 24.395 ;
        RECT 41.945 22.615 42.695 23.135 ;
        RECT 42.865 22.785 43.615 23.305 ;
        RECT 44.245 23.230 44.535 24.395 ;
        RECT 44.705 23.305 46.375 24.395 ;
        RECT 44.705 22.615 45.455 23.135 ;
        RECT 45.625 22.785 46.375 23.305 ;
        RECT 46.585 23.255 46.815 24.395 ;
        RECT 46.985 23.245 47.315 24.225 ;
        RECT 47.485 23.255 47.695 24.395 ;
        RECT 47.985 23.255 48.195 24.395 ;
        RECT 46.565 22.835 46.895 23.085 ;
        RECT 36.425 21.845 41.770 22.390 ;
        RECT 41.945 21.845 43.615 22.615 ;
        RECT 44.245 21.845 44.535 22.570 ;
        RECT 44.705 21.845 46.375 22.615 ;
        RECT 46.585 21.845 46.815 22.665 ;
        RECT 47.065 22.645 47.315 23.245 ;
        RECT 48.365 23.245 48.695 24.225 ;
        RECT 48.865 23.255 49.095 24.395 ;
        RECT 49.305 23.320 49.575 24.225 ;
        RECT 49.745 23.635 50.075 24.395 ;
        RECT 50.255 23.465 50.425 24.225 ;
        RECT 46.985 22.015 47.315 22.645 ;
        RECT 47.485 21.845 47.695 22.665 ;
        RECT 47.985 21.845 48.195 22.665 ;
        RECT 48.365 22.645 48.615 23.245 ;
        RECT 48.785 22.835 49.115 23.085 ;
        RECT 48.365 22.015 48.695 22.645 ;
        RECT 48.865 21.845 49.095 22.665 ;
        RECT 49.305 22.520 49.475 23.320 ;
        RECT 49.760 23.295 50.425 23.465 ;
        RECT 49.760 23.150 49.930 23.295 ;
        RECT 50.685 23.255 50.965 24.395 ;
        RECT 51.135 23.245 51.465 24.225 ;
        RECT 51.635 23.255 51.895 24.395 ;
        RECT 52.250 23.425 52.640 23.600 ;
        RECT 53.125 23.595 53.455 24.395 ;
        RECT 53.625 23.605 54.160 24.225 ;
        RECT 52.250 23.255 53.675 23.425 ;
        RECT 49.645 22.820 49.930 23.150 ;
        RECT 49.760 22.565 49.930 22.820 ;
        RECT 50.165 22.745 50.495 23.115 ;
        RECT 50.695 22.815 51.030 23.085 ;
        RECT 51.200 22.645 51.370 23.245 ;
        RECT 51.540 22.835 51.875 23.085 ;
        RECT 49.305 22.015 49.565 22.520 ;
        RECT 49.760 22.395 50.425 22.565 ;
        RECT 49.745 21.845 50.075 22.225 ;
        RECT 50.255 22.015 50.425 22.395 ;
        RECT 50.685 21.845 50.995 22.645 ;
        RECT 51.200 22.015 51.895 22.645 ;
        RECT 52.125 22.525 52.480 23.085 ;
        RECT 52.650 22.355 52.820 23.255 ;
        RECT 52.990 22.525 53.255 23.085 ;
        RECT 53.505 22.755 53.675 23.255 ;
        RECT 53.845 22.585 54.160 23.605 ;
        RECT 54.480 23.765 54.765 24.225 ;
        RECT 54.935 23.935 55.205 24.395 ;
        RECT 54.480 23.545 55.435 23.765 ;
        RECT 54.365 22.815 55.055 23.375 ;
        RECT 55.225 22.645 55.435 23.545 ;
        RECT 52.230 21.845 52.470 22.355 ;
        RECT 52.650 22.025 52.930 22.355 ;
        RECT 53.160 21.845 53.375 22.355 ;
        RECT 53.545 22.015 54.160 22.585 ;
        RECT 54.480 22.475 55.435 22.645 ;
        RECT 55.605 23.375 56.005 24.225 ;
        RECT 56.195 23.765 56.475 24.225 ;
        RECT 56.995 23.935 57.320 24.395 ;
        RECT 56.195 23.545 57.320 23.765 ;
        RECT 55.605 22.815 56.700 23.375 ;
        RECT 56.870 23.085 57.320 23.545 ;
        RECT 57.490 23.255 57.875 24.225 ;
        RECT 54.480 22.015 54.765 22.475 ;
        RECT 54.935 21.845 55.205 22.305 ;
        RECT 55.605 22.015 56.005 22.815 ;
        RECT 56.870 22.755 57.425 23.085 ;
        RECT 56.870 22.645 57.320 22.755 ;
        RECT 56.195 22.475 57.320 22.645 ;
        RECT 57.595 22.585 57.875 23.255 ;
        RECT 56.195 22.015 56.475 22.475 ;
        RECT 56.995 21.845 57.320 22.305 ;
        RECT 57.490 22.015 57.875 22.585 ;
        RECT 58.045 23.895 58.305 24.225 ;
        RECT 58.615 24.015 58.945 24.395 ;
        RECT 58.045 23.215 58.215 23.895 ;
        RECT 59.185 23.845 59.375 24.225 ;
        RECT 59.625 24.015 59.955 24.395 ;
        RECT 60.165 23.845 60.335 24.225 ;
        RECT 60.530 24.015 60.860 24.395 ;
        RECT 61.120 23.845 61.290 24.225 ;
        RECT 61.715 24.015 62.045 24.395 ;
        RECT 58.385 23.385 58.735 23.715 ;
        RECT 59.185 23.675 59.925 23.845 ;
        RECT 59.005 23.335 59.585 23.505 ;
        RECT 59.005 23.215 59.175 23.335 ;
        RECT 58.045 23.045 59.175 23.215 ;
        RECT 59.755 23.165 59.925 23.675 ;
        RECT 58.045 22.345 58.215 23.045 ;
        RECT 59.355 22.995 59.925 23.165 ;
        RECT 60.095 23.675 62.045 23.845 ;
        RECT 58.565 22.705 59.185 22.875 ;
        RECT 58.565 22.525 58.775 22.705 ;
        RECT 59.355 22.515 59.525 22.995 ;
        RECT 60.095 22.685 60.265 23.675 ;
        RECT 60.855 23.085 61.040 23.395 ;
        RECT 61.310 23.085 61.505 23.395 ;
        RECT 58.045 22.015 58.305 22.345 ;
        RECT 58.615 21.845 58.945 22.225 ;
        RECT 59.125 22.185 59.525 22.515 ;
        RECT 59.715 22.355 60.265 22.685 ;
        RECT 60.435 22.185 60.605 23.085 ;
        RECT 59.125 22.015 60.605 22.185 ;
        RECT 60.855 22.755 61.085 23.085 ;
        RECT 61.310 22.755 61.565 23.085 ;
        RECT 61.875 22.755 62.045 23.675 ;
        RECT 60.855 22.175 61.040 22.755 ;
        RECT 61.310 22.180 61.505 22.755 ;
        RECT 61.715 21.845 62.045 22.225 ;
        RECT 62.215 22.015 62.475 24.225 ;
        RECT 62.645 23.425 62.915 24.195 ;
        RECT 63.085 23.615 63.415 24.395 ;
        RECT 63.620 23.790 63.805 24.195 ;
        RECT 63.975 23.970 64.310 24.395 ;
        RECT 63.620 23.615 64.285 23.790 ;
        RECT 62.645 23.255 63.775 23.425 ;
        RECT 62.645 22.345 62.815 23.255 ;
        RECT 62.985 22.505 63.345 23.085 ;
        RECT 63.525 22.755 63.775 23.255 ;
        RECT 63.945 22.585 64.285 23.615 ;
        RECT 64.575 23.465 64.745 24.225 ;
        RECT 64.925 23.635 65.255 24.395 ;
        RECT 64.575 23.295 65.240 23.465 ;
        RECT 65.425 23.320 65.695 24.225 ;
        RECT 65.070 23.150 65.240 23.295 ;
        RECT 64.505 22.745 64.835 23.115 ;
        RECT 65.070 22.820 65.355 23.150 ;
        RECT 63.600 22.415 64.285 22.585 ;
        RECT 65.070 22.565 65.240 22.820 ;
        RECT 62.645 22.015 62.905 22.345 ;
        RECT 63.115 21.845 63.390 22.325 ;
        RECT 63.600 22.015 63.805 22.415 ;
        RECT 64.575 22.395 65.240 22.565 ;
        RECT 65.525 22.520 65.695 23.320 ;
        RECT 65.865 23.305 69.375 24.395 ;
        RECT 63.975 21.845 64.310 22.245 ;
        RECT 64.575 22.015 64.745 22.395 ;
        RECT 64.925 21.845 65.255 22.225 ;
        RECT 65.435 22.015 65.695 22.520 ;
        RECT 65.865 22.615 67.515 23.135 ;
        RECT 67.685 22.785 69.375 23.305 ;
        RECT 70.005 23.230 70.295 24.395 ;
        RECT 70.465 23.960 75.810 24.395 ;
        RECT 75.985 23.960 81.330 24.395 ;
        RECT 81.505 23.960 86.850 24.395 ;
        RECT 87.025 23.960 92.370 24.395 ;
        RECT 65.865 21.845 69.375 22.615 ;
        RECT 70.005 21.845 70.295 22.570 ;
        RECT 72.050 22.390 72.390 23.220 ;
        RECT 73.870 22.710 74.220 23.960 ;
        RECT 77.570 22.390 77.910 23.220 ;
        RECT 79.390 22.710 79.740 23.960 ;
        RECT 83.090 22.390 83.430 23.220 ;
        RECT 84.910 22.710 85.260 23.960 ;
        RECT 88.610 22.390 88.950 23.220 ;
        RECT 90.430 22.710 90.780 23.960 ;
        RECT 92.545 23.305 95.135 24.395 ;
        RECT 92.545 22.615 93.755 23.135 ;
        RECT 93.925 22.785 95.135 23.305 ;
        RECT 95.765 23.230 96.055 24.395 ;
        RECT 96.225 23.960 101.570 24.395 ;
        RECT 101.745 23.960 107.090 24.395 ;
        RECT 107.265 23.960 112.610 24.395 ;
        RECT 70.465 21.845 75.810 22.390 ;
        RECT 75.985 21.845 81.330 22.390 ;
        RECT 81.505 21.845 86.850 22.390 ;
        RECT 87.025 21.845 92.370 22.390 ;
        RECT 92.545 21.845 95.135 22.615 ;
        RECT 95.765 21.845 96.055 22.570 ;
        RECT 97.810 22.390 98.150 23.220 ;
        RECT 99.630 22.710 99.980 23.960 ;
        RECT 103.330 22.390 103.670 23.220 ;
        RECT 105.150 22.710 105.500 23.960 ;
        RECT 108.850 22.390 109.190 23.220 ;
        RECT 110.670 22.710 111.020 23.960 ;
        RECT 112.785 23.305 116.295 24.395 ;
        RECT 112.785 22.615 114.435 23.135 ;
        RECT 114.605 22.785 116.295 23.305 ;
        RECT 117.385 23.305 118.595 24.395 ;
        RECT 117.385 22.765 117.905 23.305 ;
        RECT 96.225 21.845 101.570 22.390 ;
        RECT 101.745 21.845 107.090 22.390 ;
        RECT 107.265 21.845 112.610 22.390 ;
        RECT 112.785 21.845 116.295 22.615 ;
        RECT 118.075 22.595 118.595 23.135 ;
        RECT 117.385 21.845 118.595 22.595 ;
        RECT 5.520 21.675 118.680 21.845 ;
        RECT 5.605 20.925 6.815 21.675 ;
        RECT 6.985 21.130 12.330 21.675 ;
        RECT 12.505 21.130 17.850 21.675 ;
        RECT 18.025 21.130 23.370 21.675 ;
        RECT 23.545 21.130 28.890 21.675 ;
        RECT 5.605 20.385 6.125 20.925 ;
        RECT 6.295 20.215 6.815 20.755 ;
        RECT 8.570 20.300 8.910 21.130 ;
        RECT 5.605 19.125 6.815 20.215 ;
        RECT 10.390 19.560 10.740 20.810 ;
        RECT 14.090 20.300 14.430 21.130 ;
        RECT 15.910 19.560 16.260 20.810 ;
        RECT 19.610 20.300 19.950 21.130 ;
        RECT 21.430 19.560 21.780 20.810 ;
        RECT 25.130 20.300 25.470 21.130 ;
        RECT 29.065 20.905 30.735 21.675 ;
        RECT 31.365 20.950 31.655 21.675 ;
        RECT 31.825 21.130 37.170 21.675 ;
        RECT 37.345 21.130 42.690 21.675 ;
        RECT 26.950 19.560 27.300 20.810 ;
        RECT 29.065 20.385 29.815 20.905 ;
        RECT 29.985 20.215 30.735 20.735 ;
        RECT 33.410 20.300 33.750 21.130 ;
        RECT 6.985 19.125 12.330 19.560 ;
        RECT 12.505 19.125 17.850 19.560 ;
        RECT 18.025 19.125 23.370 19.560 ;
        RECT 23.545 19.125 28.890 19.560 ;
        RECT 29.065 19.125 30.735 20.215 ;
        RECT 31.365 19.125 31.655 20.290 ;
        RECT 35.230 19.560 35.580 20.810 ;
        RECT 38.930 20.300 39.270 21.130 ;
        RECT 42.865 20.905 44.535 21.675 ;
        RECT 44.710 21.125 44.965 21.415 ;
        RECT 45.135 21.295 45.465 21.675 ;
        RECT 44.710 20.955 45.460 21.125 ;
        RECT 40.750 19.560 41.100 20.810 ;
        RECT 42.865 20.385 43.615 20.905 ;
        RECT 43.785 20.215 44.535 20.735 ;
        RECT 31.825 19.125 37.170 19.560 ;
        RECT 37.345 19.125 42.690 19.560 ;
        RECT 42.865 19.125 44.535 20.215 ;
        RECT 44.710 20.135 45.060 20.785 ;
        RECT 45.230 19.965 45.460 20.955 ;
        RECT 44.710 19.795 45.460 19.965 ;
        RECT 44.710 19.295 44.965 19.795 ;
        RECT 45.135 19.125 45.465 19.625 ;
        RECT 45.635 19.295 45.805 21.415 ;
        RECT 46.165 21.315 46.495 21.675 ;
        RECT 46.665 21.285 47.160 21.455 ;
        RECT 47.365 21.285 48.220 21.455 ;
        RECT 46.035 20.095 46.495 21.145 ;
        RECT 45.975 19.310 46.300 20.095 ;
        RECT 46.665 19.925 46.835 21.285 ;
        RECT 47.005 20.375 47.355 20.995 ;
        RECT 47.525 20.775 47.880 20.995 ;
        RECT 47.525 20.185 47.695 20.775 ;
        RECT 48.050 20.575 48.220 21.285 ;
        RECT 49.095 21.215 49.425 21.675 ;
        RECT 49.635 21.315 49.985 21.485 ;
        RECT 48.425 20.745 49.215 20.995 ;
        RECT 49.635 20.925 49.895 21.315 ;
        RECT 50.205 21.225 51.155 21.505 ;
        RECT 51.325 21.235 51.515 21.675 ;
        RECT 51.685 21.295 52.755 21.465 ;
        RECT 49.385 20.575 49.555 20.755 ;
        RECT 46.665 19.755 47.060 19.925 ;
        RECT 47.230 19.795 47.695 20.185 ;
        RECT 47.865 20.405 49.555 20.575 ;
        RECT 46.890 19.625 47.060 19.755 ;
        RECT 47.865 19.625 48.035 20.405 ;
        RECT 49.725 20.235 49.895 20.925 ;
        RECT 48.395 20.065 49.895 20.235 ;
        RECT 50.085 20.265 50.295 21.055 ;
        RECT 50.465 20.435 50.815 21.055 ;
        RECT 50.985 20.445 51.155 21.225 ;
        RECT 51.685 21.065 51.855 21.295 ;
        RECT 51.325 20.895 51.855 21.065 ;
        RECT 51.325 20.615 51.545 20.895 ;
        RECT 52.025 20.725 52.265 21.125 ;
        RECT 50.985 20.275 51.390 20.445 ;
        RECT 51.725 20.355 52.265 20.725 ;
        RECT 52.435 20.940 52.755 21.295 ;
        RECT 53.000 21.215 53.305 21.675 ;
        RECT 53.475 20.965 53.730 21.495 ;
        RECT 54.365 21.295 55.255 21.465 ;
        RECT 52.435 20.765 52.760 20.940 ;
        RECT 52.435 20.465 53.350 20.765 ;
        RECT 52.610 20.435 53.350 20.465 ;
        RECT 50.085 20.105 50.760 20.265 ;
        RECT 51.220 20.185 51.390 20.275 ;
        RECT 50.085 20.095 51.050 20.105 ;
        RECT 49.725 19.925 49.895 20.065 ;
        RECT 46.470 19.125 46.720 19.585 ;
        RECT 46.890 19.295 47.140 19.625 ;
        RECT 47.355 19.295 48.035 19.625 ;
        RECT 48.205 19.725 49.280 19.895 ;
        RECT 49.725 19.755 50.285 19.925 ;
        RECT 50.590 19.805 51.050 20.095 ;
        RECT 51.220 20.015 52.440 20.185 ;
        RECT 48.205 19.385 48.375 19.725 ;
        RECT 48.610 19.125 48.940 19.555 ;
        RECT 49.110 19.385 49.280 19.725 ;
        RECT 49.575 19.125 49.945 19.585 ;
        RECT 50.115 19.295 50.285 19.755 ;
        RECT 51.220 19.635 51.390 20.015 ;
        RECT 52.610 19.845 52.780 20.435 ;
        RECT 53.520 20.315 53.730 20.965 ;
        RECT 54.365 20.740 54.915 21.125 ;
        RECT 55.085 20.570 55.255 21.295 ;
        RECT 50.520 19.295 51.390 19.635 ;
        RECT 51.980 19.675 52.780 19.845 ;
        RECT 51.560 19.125 51.810 19.585 ;
        RECT 51.980 19.385 52.150 19.675 ;
        RECT 52.330 19.125 52.660 19.505 ;
        RECT 53.000 19.125 53.305 20.265 ;
        RECT 53.475 19.435 53.730 20.315 ;
        RECT 54.365 20.500 55.255 20.570 ;
        RECT 55.425 20.995 55.645 21.455 ;
        RECT 55.815 21.135 56.065 21.675 ;
        RECT 56.235 21.025 56.495 21.505 ;
        RECT 55.425 20.970 55.675 20.995 ;
        RECT 55.425 20.545 55.755 20.970 ;
        RECT 54.365 20.475 55.260 20.500 ;
        RECT 54.365 20.460 55.270 20.475 ;
        RECT 54.365 20.445 55.275 20.460 ;
        RECT 54.365 20.440 55.285 20.445 ;
        RECT 54.365 20.430 55.290 20.440 ;
        RECT 54.365 20.420 55.295 20.430 ;
        RECT 54.365 20.415 55.305 20.420 ;
        RECT 54.365 20.405 55.315 20.415 ;
        RECT 54.365 20.400 55.325 20.405 ;
        RECT 54.365 19.950 54.625 20.400 ;
        RECT 54.990 20.395 55.325 20.400 ;
        RECT 54.990 20.390 55.340 20.395 ;
        RECT 54.990 20.380 55.355 20.390 ;
        RECT 54.990 20.375 55.380 20.380 ;
        RECT 55.925 20.375 56.155 20.770 ;
        RECT 54.990 20.370 56.155 20.375 ;
        RECT 55.020 20.335 56.155 20.370 ;
        RECT 55.055 20.310 56.155 20.335 ;
        RECT 55.085 20.280 56.155 20.310 ;
        RECT 55.105 20.250 56.155 20.280 ;
        RECT 55.125 20.220 56.155 20.250 ;
        RECT 55.195 20.210 56.155 20.220 ;
        RECT 55.220 20.200 56.155 20.210 ;
        RECT 55.240 20.185 56.155 20.200 ;
        RECT 55.260 20.170 56.155 20.185 ;
        RECT 55.265 20.160 56.050 20.170 ;
        RECT 55.280 20.125 56.050 20.160 ;
        RECT 54.795 19.805 55.125 20.050 ;
        RECT 55.295 19.875 56.050 20.125 ;
        RECT 56.325 19.995 56.495 21.025 ;
        RECT 57.125 20.950 57.415 21.675 ;
        RECT 57.585 21.175 57.845 21.505 ;
        RECT 58.055 21.195 58.330 21.675 ;
        RECT 54.795 19.780 54.980 19.805 ;
        RECT 54.365 19.680 54.980 19.780 ;
        RECT 54.365 19.125 54.970 19.680 ;
        RECT 55.145 19.295 55.625 19.635 ;
        RECT 55.795 19.125 56.050 19.670 ;
        RECT 56.220 19.295 56.495 19.995 ;
        RECT 57.125 19.125 57.415 20.290 ;
        RECT 57.585 20.265 57.755 21.175 ;
        RECT 58.540 21.105 58.745 21.505 ;
        RECT 58.915 21.275 59.250 21.675 ;
        RECT 59.510 21.105 59.685 21.505 ;
        RECT 59.855 21.295 60.185 21.675 ;
        RECT 60.430 21.175 60.660 21.505 ;
        RECT 57.925 20.435 58.285 21.015 ;
        RECT 58.540 20.935 59.225 21.105 ;
        RECT 59.510 20.935 60.140 21.105 ;
        RECT 58.465 20.265 58.715 20.765 ;
        RECT 57.585 20.095 58.715 20.265 ;
        RECT 57.585 19.325 57.855 20.095 ;
        RECT 58.885 19.905 59.225 20.935 ;
        RECT 59.970 20.765 60.140 20.935 ;
        RECT 59.425 20.085 59.790 20.765 ;
        RECT 59.970 20.435 60.320 20.765 ;
        RECT 59.970 19.915 60.140 20.435 ;
        RECT 58.025 19.125 58.355 19.905 ;
        RECT 58.560 19.730 59.225 19.905 ;
        RECT 59.510 19.745 60.140 19.915 ;
        RECT 60.490 19.885 60.660 21.175 ;
        RECT 60.860 20.065 61.140 21.340 ;
        RECT 61.365 21.335 61.635 21.340 ;
        RECT 61.325 21.165 61.635 21.335 ;
        RECT 62.095 21.295 62.425 21.675 ;
        RECT 62.595 21.420 62.930 21.465 ;
        RECT 61.365 20.065 61.635 21.165 ;
        RECT 61.825 20.065 62.165 21.095 ;
        RECT 62.595 20.955 62.935 21.420 ;
        RECT 63.415 21.205 63.585 21.675 ;
        RECT 63.755 21.025 64.085 21.505 ;
        RECT 64.255 21.205 64.425 21.675 ;
        RECT 64.595 21.025 64.925 21.505 ;
        RECT 62.335 20.435 62.595 20.765 ;
        RECT 62.335 19.885 62.505 20.435 ;
        RECT 62.765 20.265 62.935 20.955 ;
        RECT 58.560 19.325 58.745 19.730 ;
        RECT 58.915 19.125 59.250 19.550 ;
        RECT 59.510 19.295 59.685 19.745 ;
        RECT 60.490 19.715 62.505 19.885 ;
        RECT 59.855 19.125 60.185 19.565 ;
        RECT 60.490 19.295 60.660 19.715 ;
        RECT 60.895 19.125 61.565 19.535 ;
        RECT 61.780 19.295 61.950 19.715 ;
        RECT 62.150 19.125 62.480 19.535 ;
        RECT 62.675 19.295 62.935 20.265 ;
        RECT 63.160 20.855 64.925 21.025 ;
        RECT 65.095 20.865 65.265 21.675 ;
        RECT 65.465 21.295 66.535 21.465 ;
        RECT 65.465 20.940 65.785 21.295 ;
        RECT 63.160 20.305 63.570 20.855 ;
        RECT 65.460 20.685 65.785 20.940 ;
        RECT 63.755 20.475 65.785 20.685 ;
        RECT 65.440 20.465 65.785 20.475 ;
        RECT 65.955 20.725 66.195 21.125 ;
        RECT 66.365 21.065 66.535 21.295 ;
        RECT 66.705 21.235 66.895 21.675 ;
        RECT 67.065 21.225 68.015 21.505 ;
        RECT 68.235 21.315 68.585 21.485 ;
        RECT 66.365 20.895 66.895 21.065 ;
        RECT 63.160 20.135 64.885 20.305 ;
        RECT 63.415 19.125 63.585 19.965 ;
        RECT 63.795 19.295 64.045 20.135 ;
        RECT 64.255 19.125 64.425 19.965 ;
        RECT 64.595 19.295 64.885 20.135 ;
        RECT 65.095 19.125 65.265 20.185 ;
        RECT 65.440 19.845 65.610 20.465 ;
        RECT 65.955 20.355 66.495 20.725 ;
        RECT 66.675 20.615 66.895 20.895 ;
        RECT 67.065 20.445 67.235 21.225 ;
        RECT 66.830 20.275 67.235 20.445 ;
        RECT 67.405 20.435 67.755 21.055 ;
        RECT 66.830 20.185 67.000 20.275 ;
        RECT 67.925 20.265 68.135 21.055 ;
        RECT 65.780 20.015 67.000 20.185 ;
        RECT 67.460 20.105 68.135 20.265 ;
        RECT 65.440 19.675 66.240 19.845 ;
        RECT 65.560 19.125 65.890 19.505 ;
        RECT 66.070 19.385 66.240 19.675 ;
        RECT 66.830 19.635 67.000 20.015 ;
        RECT 67.170 20.095 68.135 20.105 ;
        RECT 68.325 20.925 68.585 21.315 ;
        RECT 68.795 21.215 69.125 21.675 ;
        RECT 70.000 21.285 70.855 21.455 ;
        RECT 71.060 21.285 71.555 21.455 ;
        RECT 71.725 21.315 72.055 21.675 ;
        RECT 68.325 20.235 68.495 20.925 ;
        RECT 68.665 20.575 68.835 20.755 ;
        RECT 69.005 20.745 69.795 20.995 ;
        RECT 70.000 20.575 70.170 21.285 ;
        RECT 70.340 20.775 70.695 20.995 ;
        RECT 68.665 20.405 70.355 20.575 ;
        RECT 67.170 19.805 67.630 20.095 ;
        RECT 68.325 20.065 69.825 20.235 ;
        RECT 68.325 19.925 68.495 20.065 ;
        RECT 67.935 19.755 68.495 19.925 ;
        RECT 66.410 19.125 66.660 19.585 ;
        RECT 66.830 19.295 67.700 19.635 ;
        RECT 67.935 19.295 68.105 19.755 ;
        RECT 68.940 19.725 70.015 19.895 ;
        RECT 68.275 19.125 68.645 19.585 ;
        RECT 68.940 19.385 69.110 19.725 ;
        RECT 69.280 19.125 69.610 19.555 ;
        RECT 69.845 19.385 70.015 19.725 ;
        RECT 70.185 19.625 70.355 20.405 ;
        RECT 70.525 20.185 70.695 20.775 ;
        RECT 70.865 20.375 71.215 20.995 ;
        RECT 70.525 19.795 70.990 20.185 ;
        RECT 71.385 19.925 71.555 21.285 ;
        RECT 71.725 20.095 72.185 21.145 ;
        RECT 71.160 19.755 71.555 19.925 ;
        RECT 71.160 19.625 71.330 19.755 ;
        RECT 70.185 19.295 70.865 19.625 ;
        RECT 71.080 19.295 71.330 19.625 ;
        RECT 71.500 19.125 71.750 19.585 ;
        RECT 71.920 19.310 72.245 20.095 ;
        RECT 72.415 19.295 72.585 21.415 ;
        RECT 72.755 21.295 73.085 21.675 ;
        RECT 73.255 21.125 73.510 21.415 ;
        RECT 73.685 21.130 79.030 21.675 ;
        RECT 72.760 20.955 73.510 21.125 ;
        RECT 72.760 19.965 72.990 20.955 ;
        RECT 73.160 20.135 73.510 20.785 ;
        RECT 75.270 20.300 75.610 21.130 ;
        RECT 79.205 20.905 82.715 21.675 ;
        RECT 82.885 20.950 83.175 21.675 ;
        RECT 83.345 21.130 88.690 21.675 ;
        RECT 88.865 21.130 94.210 21.675 ;
        RECT 94.385 21.130 99.730 21.675 ;
        RECT 99.905 21.130 105.250 21.675 ;
        RECT 72.760 19.795 73.510 19.965 ;
        RECT 72.755 19.125 73.085 19.625 ;
        RECT 73.255 19.295 73.510 19.795 ;
        RECT 77.090 19.560 77.440 20.810 ;
        RECT 79.205 20.385 80.855 20.905 ;
        RECT 81.025 20.215 82.715 20.735 ;
        RECT 84.930 20.300 85.270 21.130 ;
        RECT 73.685 19.125 79.030 19.560 ;
        RECT 79.205 19.125 82.715 20.215 ;
        RECT 82.885 19.125 83.175 20.290 ;
        RECT 86.750 19.560 87.100 20.810 ;
        RECT 90.450 20.300 90.790 21.130 ;
        RECT 92.270 19.560 92.620 20.810 ;
        RECT 95.970 20.300 96.310 21.130 ;
        RECT 97.790 19.560 98.140 20.810 ;
        RECT 101.490 20.300 101.830 21.130 ;
        RECT 105.425 20.905 108.015 21.675 ;
        RECT 108.645 20.950 108.935 21.675 ;
        RECT 109.105 21.130 114.450 21.675 ;
        RECT 103.310 19.560 103.660 20.810 ;
        RECT 105.425 20.385 106.635 20.905 ;
        RECT 106.805 20.215 108.015 20.735 ;
        RECT 110.690 20.300 111.030 21.130 ;
        RECT 114.625 20.905 117.215 21.675 ;
        RECT 117.385 20.925 118.595 21.675 ;
        RECT 83.345 19.125 88.690 19.560 ;
        RECT 88.865 19.125 94.210 19.560 ;
        RECT 94.385 19.125 99.730 19.560 ;
        RECT 99.905 19.125 105.250 19.560 ;
        RECT 105.425 19.125 108.015 20.215 ;
        RECT 108.645 19.125 108.935 20.290 ;
        RECT 112.510 19.560 112.860 20.810 ;
        RECT 114.625 20.385 115.835 20.905 ;
        RECT 116.005 20.215 117.215 20.735 ;
        RECT 109.105 19.125 114.450 19.560 ;
        RECT 114.625 19.125 117.215 20.215 ;
        RECT 117.385 20.215 117.905 20.755 ;
        RECT 118.075 20.385 118.595 20.925 ;
        RECT 117.385 19.125 118.595 20.215 ;
        RECT 5.520 18.955 118.680 19.125 ;
        RECT 5.605 17.865 6.815 18.955 ;
        RECT 6.985 18.520 12.330 18.955 ;
        RECT 12.505 18.520 17.850 18.955 ;
        RECT 5.605 17.155 6.125 17.695 ;
        RECT 6.295 17.325 6.815 17.865 ;
        RECT 5.605 16.405 6.815 17.155 ;
        RECT 8.570 16.950 8.910 17.780 ;
        RECT 10.390 17.270 10.740 18.520 ;
        RECT 14.090 16.950 14.430 17.780 ;
        RECT 15.910 17.270 16.260 18.520 ;
        RECT 18.485 17.790 18.775 18.955 ;
        RECT 18.945 18.520 24.290 18.955 ;
        RECT 24.465 18.520 29.810 18.955 ;
        RECT 29.985 18.520 35.330 18.955 ;
        RECT 35.505 18.520 40.850 18.955 ;
        RECT 6.985 16.405 12.330 16.950 ;
        RECT 12.505 16.405 17.850 16.950 ;
        RECT 18.485 16.405 18.775 17.130 ;
        RECT 20.530 16.950 20.870 17.780 ;
        RECT 22.350 17.270 22.700 18.520 ;
        RECT 26.050 16.950 26.390 17.780 ;
        RECT 27.870 17.270 28.220 18.520 ;
        RECT 31.570 16.950 31.910 17.780 ;
        RECT 33.390 17.270 33.740 18.520 ;
        RECT 37.090 16.950 37.430 17.780 ;
        RECT 38.910 17.270 39.260 18.520 ;
        RECT 41.025 17.865 43.615 18.955 ;
        RECT 41.025 17.175 42.235 17.695 ;
        RECT 42.405 17.345 43.615 17.865 ;
        RECT 44.245 17.790 44.535 18.955 ;
        RECT 44.705 17.865 46.375 18.955 ;
        RECT 46.550 18.285 46.805 18.785 ;
        RECT 46.975 18.455 47.305 18.955 ;
        RECT 46.550 18.115 47.300 18.285 ;
        RECT 44.705 17.175 45.455 17.695 ;
        RECT 45.625 17.345 46.375 17.865 ;
        RECT 46.550 17.295 46.900 17.945 ;
        RECT 18.945 16.405 24.290 16.950 ;
        RECT 24.465 16.405 29.810 16.950 ;
        RECT 29.985 16.405 35.330 16.950 ;
        RECT 35.505 16.405 40.850 16.950 ;
        RECT 41.025 16.405 43.615 17.175 ;
        RECT 44.245 16.405 44.535 17.130 ;
        RECT 44.705 16.405 46.375 17.175 ;
        RECT 47.070 17.125 47.300 18.115 ;
        RECT 46.550 16.955 47.300 17.125 ;
        RECT 46.550 16.665 46.805 16.955 ;
        RECT 46.975 16.405 47.305 16.785 ;
        RECT 47.475 16.665 47.645 18.785 ;
        RECT 47.815 17.985 48.140 18.770 ;
        RECT 48.310 18.495 48.560 18.955 ;
        RECT 48.730 18.455 48.980 18.785 ;
        RECT 49.195 18.455 49.875 18.785 ;
        RECT 48.730 18.325 48.900 18.455 ;
        RECT 48.505 18.155 48.900 18.325 ;
        RECT 47.875 16.935 48.335 17.985 ;
        RECT 48.505 16.795 48.675 18.155 ;
        RECT 49.070 17.895 49.535 18.285 ;
        RECT 48.845 17.085 49.195 17.705 ;
        RECT 49.365 17.305 49.535 17.895 ;
        RECT 49.705 17.675 49.875 18.455 ;
        RECT 50.045 18.355 50.215 18.695 ;
        RECT 50.450 18.525 50.780 18.955 ;
        RECT 50.950 18.355 51.120 18.695 ;
        RECT 51.415 18.495 51.785 18.955 ;
        RECT 50.045 18.185 51.120 18.355 ;
        RECT 51.955 18.325 52.125 18.785 ;
        RECT 52.360 18.445 53.230 18.785 ;
        RECT 53.400 18.495 53.650 18.955 ;
        RECT 51.565 18.155 52.125 18.325 ;
        RECT 51.565 18.015 51.735 18.155 ;
        RECT 50.235 17.845 51.735 18.015 ;
        RECT 52.430 17.985 52.890 18.275 ;
        RECT 49.705 17.505 51.395 17.675 ;
        RECT 49.365 17.085 49.720 17.305 ;
        RECT 49.890 16.795 50.060 17.505 ;
        RECT 50.265 17.085 51.055 17.335 ;
        RECT 51.225 17.325 51.395 17.505 ;
        RECT 51.565 17.155 51.735 17.845 ;
        RECT 48.005 16.405 48.335 16.765 ;
        RECT 48.505 16.625 49.000 16.795 ;
        RECT 49.205 16.625 50.060 16.795 ;
        RECT 50.935 16.405 51.265 16.865 ;
        RECT 51.475 16.765 51.735 17.155 ;
        RECT 51.925 17.975 52.890 17.985 ;
        RECT 53.060 18.065 53.230 18.445 ;
        RECT 53.820 18.405 53.990 18.695 ;
        RECT 54.170 18.575 54.500 18.955 ;
        RECT 53.820 18.235 54.620 18.405 ;
        RECT 51.925 17.815 52.600 17.975 ;
        RECT 53.060 17.895 54.280 18.065 ;
        RECT 51.925 17.025 52.135 17.815 ;
        RECT 53.060 17.805 53.230 17.895 ;
        RECT 52.305 17.025 52.655 17.645 ;
        RECT 52.825 17.635 53.230 17.805 ;
        RECT 52.825 16.855 52.995 17.635 ;
        RECT 53.165 17.185 53.385 17.465 ;
        RECT 53.565 17.355 54.105 17.725 ;
        RECT 54.450 17.645 54.620 18.235 ;
        RECT 54.840 17.815 55.145 18.955 ;
        RECT 55.315 17.765 55.570 18.645 ;
        RECT 55.750 18.285 56.005 18.785 ;
        RECT 56.175 18.455 56.505 18.955 ;
        RECT 55.750 18.115 56.500 18.285 ;
        RECT 54.450 17.615 55.190 17.645 ;
        RECT 53.165 17.015 53.695 17.185 ;
        RECT 51.475 16.595 51.825 16.765 ;
        RECT 52.045 16.575 52.995 16.855 ;
        RECT 53.165 16.405 53.355 16.845 ;
        RECT 53.525 16.785 53.695 17.015 ;
        RECT 53.865 16.955 54.105 17.355 ;
        RECT 54.275 17.315 55.190 17.615 ;
        RECT 54.275 17.140 54.600 17.315 ;
        RECT 54.275 16.785 54.595 17.140 ;
        RECT 55.360 17.115 55.570 17.765 ;
        RECT 55.750 17.295 56.100 17.945 ;
        RECT 56.270 17.125 56.500 18.115 ;
        RECT 53.525 16.615 54.595 16.785 ;
        RECT 54.840 16.405 55.145 16.865 ;
        RECT 55.315 16.585 55.570 17.115 ;
        RECT 55.750 16.955 56.500 17.125 ;
        RECT 55.750 16.665 56.005 16.955 ;
        RECT 56.175 16.405 56.505 16.785 ;
        RECT 56.675 16.665 56.845 18.785 ;
        RECT 57.015 17.985 57.340 18.770 ;
        RECT 57.510 18.495 57.760 18.955 ;
        RECT 57.930 18.455 58.180 18.785 ;
        RECT 58.395 18.455 59.075 18.785 ;
        RECT 57.930 18.325 58.100 18.455 ;
        RECT 57.705 18.155 58.100 18.325 ;
        RECT 57.075 16.935 57.535 17.985 ;
        RECT 57.705 16.795 57.875 18.155 ;
        RECT 58.270 17.895 58.735 18.285 ;
        RECT 58.045 17.085 58.395 17.705 ;
        RECT 58.565 17.305 58.735 17.895 ;
        RECT 58.905 17.675 59.075 18.455 ;
        RECT 59.245 18.355 59.415 18.695 ;
        RECT 59.650 18.525 59.980 18.955 ;
        RECT 60.150 18.355 60.320 18.695 ;
        RECT 60.615 18.495 60.985 18.955 ;
        RECT 59.245 18.185 60.320 18.355 ;
        RECT 61.155 18.325 61.325 18.785 ;
        RECT 61.560 18.445 62.430 18.785 ;
        RECT 62.600 18.495 62.850 18.955 ;
        RECT 60.765 18.155 61.325 18.325 ;
        RECT 60.765 18.015 60.935 18.155 ;
        RECT 59.435 17.845 60.935 18.015 ;
        RECT 61.630 17.985 62.090 18.275 ;
        RECT 58.905 17.505 60.595 17.675 ;
        RECT 58.565 17.085 58.920 17.305 ;
        RECT 59.090 16.795 59.260 17.505 ;
        RECT 59.465 17.085 60.255 17.335 ;
        RECT 60.425 17.325 60.595 17.505 ;
        RECT 60.765 17.155 60.935 17.845 ;
        RECT 57.205 16.405 57.535 16.765 ;
        RECT 57.705 16.625 58.200 16.795 ;
        RECT 58.405 16.625 59.260 16.795 ;
        RECT 60.135 16.405 60.465 16.865 ;
        RECT 60.675 16.765 60.935 17.155 ;
        RECT 61.125 17.975 62.090 17.985 ;
        RECT 62.260 18.065 62.430 18.445 ;
        RECT 63.020 18.405 63.190 18.695 ;
        RECT 63.370 18.575 63.700 18.955 ;
        RECT 63.020 18.235 63.820 18.405 ;
        RECT 61.125 17.815 61.800 17.975 ;
        RECT 62.260 17.895 63.480 18.065 ;
        RECT 61.125 17.025 61.335 17.815 ;
        RECT 62.260 17.805 62.430 17.895 ;
        RECT 61.505 17.025 61.855 17.645 ;
        RECT 62.025 17.635 62.430 17.805 ;
        RECT 62.025 16.855 62.195 17.635 ;
        RECT 62.365 17.185 62.585 17.465 ;
        RECT 62.765 17.355 63.305 17.725 ;
        RECT 63.650 17.645 63.820 18.235 ;
        RECT 64.040 17.815 64.345 18.955 ;
        RECT 64.515 17.765 64.770 18.645 ;
        RECT 65.005 17.815 65.215 18.955 ;
        RECT 63.650 17.615 64.390 17.645 ;
        RECT 62.365 17.015 62.895 17.185 ;
        RECT 60.675 16.595 61.025 16.765 ;
        RECT 61.245 16.575 62.195 16.855 ;
        RECT 62.365 16.405 62.555 16.845 ;
        RECT 62.725 16.785 62.895 17.015 ;
        RECT 63.065 16.955 63.305 17.355 ;
        RECT 63.475 17.315 64.390 17.615 ;
        RECT 63.475 17.140 63.800 17.315 ;
        RECT 63.475 16.785 63.795 17.140 ;
        RECT 64.560 17.115 64.770 17.765 ;
        RECT 65.385 17.805 65.715 18.785 ;
        RECT 65.885 17.815 66.115 18.955 ;
        RECT 67.285 17.815 67.515 18.955 ;
        RECT 67.685 17.805 68.015 18.785 ;
        RECT 68.185 17.815 68.395 18.955 ;
        RECT 68.625 17.865 69.835 18.955 ;
        RECT 62.725 16.615 63.795 16.785 ;
        RECT 64.040 16.405 64.345 16.865 ;
        RECT 64.515 16.585 64.770 17.115 ;
        RECT 65.005 16.405 65.215 17.225 ;
        RECT 65.385 17.205 65.635 17.805 ;
        RECT 65.805 17.395 66.135 17.645 ;
        RECT 67.265 17.395 67.595 17.645 ;
        RECT 65.385 16.575 65.715 17.205 ;
        RECT 65.885 16.405 66.115 17.225 ;
        RECT 67.285 16.405 67.515 17.225 ;
        RECT 67.765 17.205 68.015 17.805 ;
        RECT 67.685 16.575 68.015 17.205 ;
        RECT 68.185 16.405 68.395 17.225 ;
        RECT 68.625 17.155 69.145 17.695 ;
        RECT 69.315 17.325 69.835 17.865 ;
        RECT 70.005 17.790 70.295 18.955 ;
        RECT 70.465 18.520 75.810 18.955 ;
        RECT 75.985 18.520 81.330 18.955 ;
        RECT 81.505 18.520 86.850 18.955 ;
        RECT 87.025 18.520 92.370 18.955 ;
        RECT 68.625 16.405 69.835 17.155 ;
        RECT 70.005 16.405 70.295 17.130 ;
        RECT 72.050 16.950 72.390 17.780 ;
        RECT 73.870 17.270 74.220 18.520 ;
        RECT 77.570 16.950 77.910 17.780 ;
        RECT 79.390 17.270 79.740 18.520 ;
        RECT 83.090 16.950 83.430 17.780 ;
        RECT 84.910 17.270 85.260 18.520 ;
        RECT 88.610 16.950 88.950 17.780 ;
        RECT 90.430 17.270 90.780 18.520 ;
        RECT 92.545 17.865 95.135 18.955 ;
        RECT 92.545 17.175 93.755 17.695 ;
        RECT 93.925 17.345 95.135 17.865 ;
        RECT 95.765 17.790 96.055 18.955 ;
        RECT 96.225 18.520 101.570 18.955 ;
        RECT 101.745 18.520 107.090 18.955 ;
        RECT 107.265 18.520 112.610 18.955 ;
        RECT 70.465 16.405 75.810 16.950 ;
        RECT 75.985 16.405 81.330 16.950 ;
        RECT 81.505 16.405 86.850 16.950 ;
        RECT 87.025 16.405 92.370 16.950 ;
        RECT 92.545 16.405 95.135 17.175 ;
        RECT 95.765 16.405 96.055 17.130 ;
        RECT 97.810 16.950 98.150 17.780 ;
        RECT 99.630 17.270 99.980 18.520 ;
        RECT 103.330 16.950 103.670 17.780 ;
        RECT 105.150 17.270 105.500 18.520 ;
        RECT 108.850 16.950 109.190 17.780 ;
        RECT 110.670 17.270 111.020 18.520 ;
        RECT 112.785 17.865 116.295 18.955 ;
        RECT 112.785 17.175 114.435 17.695 ;
        RECT 114.605 17.345 116.295 17.865 ;
        RECT 117.385 17.865 118.595 18.955 ;
        RECT 117.385 17.325 117.905 17.865 ;
        RECT 96.225 16.405 101.570 16.950 ;
        RECT 101.745 16.405 107.090 16.950 ;
        RECT 107.265 16.405 112.610 16.950 ;
        RECT 112.785 16.405 116.295 17.175 ;
        RECT 118.075 17.155 118.595 17.695 ;
        RECT 117.385 16.405 118.595 17.155 ;
        RECT 5.520 16.235 118.680 16.405 ;
        RECT 5.605 15.485 6.815 16.235 ;
        RECT 6.985 15.690 12.330 16.235 ;
        RECT 12.505 15.690 17.850 16.235 ;
        RECT 18.025 15.690 23.370 16.235 ;
        RECT 23.545 15.690 28.890 16.235 ;
        RECT 5.605 14.945 6.125 15.485 ;
        RECT 6.295 14.775 6.815 15.315 ;
        RECT 8.570 14.860 8.910 15.690 ;
        RECT 5.605 13.685 6.815 14.775 ;
        RECT 10.390 14.120 10.740 15.370 ;
        RECT 14.090 14.860 14.430 15.690 ;
        RECT 15.910 14.120 16.260 15.370 ;
        RECT 19.610 14.860 19.950 15.690 ;
        RECT 21.430 14.120 21.780 15.370 ;
        RECT 25.130 14.860 25.470 15.690 ;
        RECT 29.065 15.465 30.735 16.235 ;
        RECT 31.365 15.510 31.655 16.235 ;
        RECT 31.825 15.690 37.170 16.235 ;
        RECT 37.345 15.690 42.690 16.235 ;
        RECT 42.865 15.690 48.210 16.235 ;
        RECT 26.950 14.120 27.300 15.370 ;
        RECT 29.065 14.945 29.815 15.465 ;
        RECT 29.985 14.775 30.735 15.295 ;
        RECT 33.410 14.860 33.750 15.690 ;
        RECT 6.985 13.685 12.330 14.120 ;
        RECT 12.505 13.685 17.850 14.120 ;
        RECT 18.025 13.685 23.370 14.120 ;
        RECT 23.545 13.685 28.890 14.120 ;
        RECT 29.065 13.685 30.735 14.775 ;
        RECT 31.365 13.685 31.655 14.850 ;
        RECT 35.230 14.120 35.580 15.370 ;
        RECT 38.930 14.860 39.270 15.690 ;
        RECT 40.750 14.120 41.100 15.370 ;
        RECT 44.450 14.860 44.790 15.690 ;
        RECT 48.385 15.465 51.895 16.235 ;
        RECT 52.985 15.495 53.450 16.040 ;
        RECT 46.270 14.120 46.620 15.370 ;
        RECT 48.385 14.945 50.035 15.465 ;
        RECT 50.205 14.775 51.895 15.295 ;
        RECT 31.825 13.685 37.170 14.120 ;
        RECT 37.345 13.685 42.690 14.120 ;
        RECT 42.865 13.685 48.210 14.120 ;
        RECT 48.385 13.685 51.895 14.775 ;
        RECT 52.985 14.535 53.155 15.495 ;
        RECT 53.955 15.415 54.125 16.235 ;
        RECT 54.295 15.585 54.625 16.065 ;
        RECT 54.795 15.845 55.145 16.235 ;
        RECT 55.315 15.665 55.545 16.065 ;
        RECT 55.035 15.585 55.545 15.665 ;
        RECT 54.295 15.495 55.545 15.585 ;
        RECT 55.715 15.495 56.035 15.975 ;
        RECT 57.125 15.510 57.415 16.235 ;
        RECT 54.295 15.415 55.205 15.495 ;
        RECT 53.325 14.875 53.570 15.325 ;
        RECT 53.830 15.045 54.525 15.245 ;
        RECT 54.695 15.075 55.295 15.245 ;
        RECT 54.695 14.875 54.865 15.075 ;
        RECT 55.525 14.905 55.695 15.325 ;
        RECT 53.325 14.705 54.865 14.875 ;
        RECT 55.035 14.735 55.695 14.905 ;
        RECT 55.035 14.535 55.205 14.735 ;
        RECT 55.865 14.565 56.035 15.495 ;
        RECT 57.590 15.395 57.850 16.235 ;
        RECT 58.025 15.490 58.280 16.065 ;
        RECT 58.450 15.855 58.780 16.235 ;
        RECT 58.995 15.685 59.165 16.065 ;
        RECT 58.450 15.515 59.165 15.685 ;
        RECT 52.985 14.365 55.205 14.535 ;
        RECT 55.375 14.365 56.035 14.565 ;
        RECT 52.985 13.685 53.285 14.195 ;
        RECT 53.455 13.855 53.785 14.365 ;
        RECT 55.375 14.195 55.545 14.365 ;
        RECT 53.955 13.685 54.585 14.195 ;
        RECT 55.165 14.025 55.545 14.195 ;
        RECT 55.715 13.685 56.015 14.195 ;
        RECT 57.125 13.685 57.415 14.850 ;
        RECT 57.590 13.685 57.850 14.835 ;
        RECT 58.025 14.760 58.195 15.490 ;
        RECT 58.450 15.325 58.620 15.515 ;
        RECT 59.485 15.415 59.695 16.235 ;
        RECT 59.865 15.435 60.195 16.065 ;
        RECT 58.365 14.995 58.620 15.325 ;
        RECT 58.450 14.785 58.620 14.995 ;
        RECT 58.900 14.965 59.255 15.335 ;
        RECT 59.865 14.835 60.115 15.435 ;
        RECT 60.365 15.415 60.595 16.235 ;
        RECT 60.805 15.690 66.150 16.235 ;
        RECT 66.325 15.690 71.670 16.235 ;
        RECT 71.845 15.690 77.190 16.235 ;
        RECT 77.365 15.690 82.710 16.235 ;
        RECT 60.285 14.995 60.615 15.245 ;
        RECT 62.390 14.860 62.730 15.690 ;
        RECT 58.025 13.855 58.280 14.760 ;
        RECT 58.450 14.615 59.165 14.785 ;
        RECT 58.450 13.685 58.780 14.445 ;
        RECT 58.995 13.855 59.165 14.615 ;
        RECT 59.485 13.685 59.695 14.825 ;
        RECT 59.865 13.855 60.195 14.835 ;
        RECT 60.365 13.685 60.595 14.825 ;
        RECT 64.210 14.120 64.560 15.370 ;
        RECT 67.910 14.860 68.250 15.690 ;
        RECT 69.730 14.120 70.080 15.370 ;
        RECT 73.430 14.860 73.770 15.690 ;
        RECT 75.250 14.120 75.600 15.370 ;
        RECT 78.950 14.860 79.290 15.690 ;
        RECT 82.885 15.510 83.175 16.235 ;
        RECT 83.345 15.690 88.690 16.235 ;
        RECT 88.865 15.690 94.210 16.235 ;
        RECT 94.385 15.690 99.730 16.235 ;
        RECT 99.905 15.690 105.250 16.235 ;
        RECT 80.770 14.120 81.120 15.370 ;
        RECT 84.930 14.860 85.270 15.690 ;
        RECT 60.805 13.685 66.150 14.120 ;
        RECT 66.325 13.685 71.670 14.120 ;
        RECT 71.845 13.685 77.190 14.120 ;
        RECT 77.365 13.685 82.710 14.120 ;
        RECT 82.885 13.685 83.175 14.850 ;
        RECT 86.750 14.120 87.100 15.370 ;
        RECT 90.450 14.860 90.790 15.690 ;
        RECT 92.270 14.120 92.620 15.370 ;
        RECT 95.970 14.860 96.310 15.690 ;
        RECT 97.790 14.120 98.140 15.370 ;
        RECT 101.490 14.860 101.830 15.690 ;
        RECT 105.425 15.465 108.015 16.235 ;
        RECT 108.645 15.510 108.935 16.235 ;
        RECT 109.105 15.690 114.450 16.235 ;
        RECT 103.310 14.120 103.660 15.370 ;
        RECT 105.425 14.945 106.635 15.465 ;
        RECT 106.805 14.775 108.015 15.295 ;
        RECT 110.690 14.860 111.030 15.690 ;
        RECT 114.625 15.465 117.215 16.235 ;
        RECT 117.385 15.485 118.595 16.235 ;
        RECT 83.345 13.685 88.690 14.120 ;
        RECT 88.865 13.685 94.210 14.120 ;
        RECT 94.385 13.685 99.730 14.120 ;
        RECT 99.905 13.685 105.250 14.120 ;
        RECT 105.425 13.685 108.015 14.775 ;
        RECT 108.645 13.685 108.935 14.850 ;
        RECT 112.510 14.120 112.860 15.370 ;
        RECT 114.625 14.945 115.835 15.465 ;
        RECT 116.005 14.775 117.215 15.295 ;
        RECT 109.105 13.685 114.450 14.120 ;
        RECT 114.625 13.685 117.215 14.775 ;
        RECT 117.385 14.775 117.905 15.315 ;
        RECT 118.075 14.945 118.595 15.485 ;
        RECT 117.385 13.685 118.595 14.775 ;
        RECT 5.520 13.515 118.680 13.685 ;
        RECT 5.605 12.425 6.815 13.515 ;
        RECT 6.985 13.080 12.330 13.515 ;
        RECT 12.505 13.080 17.850 13.515 ;
        RECT 5.605 11.715 6.125 12.255 ;
        RECT 6.295 11.885 6.815 12.425 ;
        RECT 5.605 10.965 6.815 11.715 ;
        RECT 8.570 11.510 8.910 12.340 ;
        RECT 10.390 11.830 10.740 13.080 ;
        RECT 14.090 11.510 14.430 12.340 ;
        RECT 15.910 11.830 16.260 13.080 ;
        RECT 18.485 12.350 18.775 13.515 ;
        RECT 18.945 13.080 24.290 13.515 ;
        RECT 24.465 13.080 29.810 13.515 ;
        RECT 6.985 10.965 12.330 11.510 ;
        RECT 12.505 10.965 17.850 11.510 ;
        RECT 18.485 10.965 18.775 11.690 ;
        RECT 20.530 11.510 20.870 12.340 ;
        RECT 22.350 11.830 22.700 13.080 ;
        RECT 26.050 11.510 26.390 12.340 ;
        RECT 27.870 11.830 28.220 13.080 ;
        RECT 29.985 12.425 31.195 13.515 ;
        RECT 29.985 11.715 30.505 12.255 ;
        RECT 30.675 11.885 31.195 12.425 ;
        RECT 31.365 12.350 31.655 13.515 ;
        RECT 31.825 13.080 37.170 13.515 ;
        RECT 37.345 13.080 42.690 13.515 ;
        RECT 18.945 10.965 24.290 11.510 ;
        RECT 24.465 10.965 29.810 11.510 ;
        RECT 29.985 10.965 31.195 11.715 ;
        RECT 31.365 10.965 31.655 11.690 ;
        RECT 33.410 11.510 33.750 12.340 ;
        RECT 35.230 11.830 35.580 13.080 ;
        RECT 38.930 11.510 39.270 12.340 ;
        RECT 40.750 11.830 41.100 13.080 ;
        RECT 42.865 12.425 44.075 13.515 ;
        RECT 42.865 11.715 43.385 12.255 ;
        RECT 43.555 11.885 44.075 12.425 ;
        RECT 44.245 12.350 44.535 13.515 ;
        RECT 44.705 13.080 50.050 13.515 ;
        RECT 50.225 13.080 55.570 13.515 ;
        RECT 31.825 10.965 37.170 11.510 ;
        RECT 37.345 10.965 42.690 11.510 ;
        RECT 42.865 10.965 44.075 11.715 ;
        RECT 44.245 10.965 44.535 11.690 ;
        RECT 46.290 11.510 46.630 12.340 ;
        RECT 48.110 11.830 48.460 13.080 ;
        RECT 51.810 11.510 52.150 12.340 ;
        RECT 53.630 11.830 53.980 13.080 ;
        RECT 55.745 12.425 56.955 13.515 ;
        RECT 55.745 11.715 56.265 12.255 ;
        RECT 56.435 11.885 56.955 12.425 ;
        RECT 57.125 12.350 57.415 13.515 ;
        RECT 57.585 13.080 62.930 13.515 ;
        RECT 63.105 13.080 68.450 13.515 ;
        RECT 44.705 10.965 50.050 11.510 ;
        RECT 50.225 10.965 55.570 11.510 ;
        RECT 55.745 10.965 56.955 11.715 ;
        RECT 57.125 10.965 57.415 11.690 ;
        RECT 59.170 11.510 59.510 12.340 ;
        RECT 60.990 11.830 61.340 13.080 ;
        RECT 64.690 11.510 65.030 12.340 ;
        RECT 66.510 11.830 66.860 13.080 ;
        RECT 68.625 12.425 69.835 13.515 ;
        RECT 68.625 11.715 69.145 12.255 ;
        RECT 69.315 11.885 69.835 12.425 ;
        RECT 70.005 12.350 70.295 13.515 ;
        RECT 70.465 13.080 75.810 13.515 ;
        RECT 75.985 13.080 81.330 13.515 ;
        RECT 57.585 10.965 62.930 11.510 ;
        RECT 63.105 10.965 68.450 11.510 ;
        RECT 68.625 10.965 69.835 11.715 ;
        RECT 70.005 10.965 70.295 11.690 ;
        RECT 72.050 11.510 72.390 12.340 ;
        RECT 73.870 11.830 74.220 13.080 ;
        RECT 77.570 11.510 77.910 12.340 ;
        RECT 79.390 11.830 79.740 13.080 ;
        RECT 81.505 12.425 82.715 13.515 ;
        RECT 81.505 11.715 82.025 12.255 ;
        RECT 82.195 11.885 82.715 12.425 ;
        RECT 82.885 12.350 83.175 13.515 ;
        RECT 83.345 13.080 88.690 13.515 ;
        RECT 88.865 13.080 94.210 13.515 ;
        RECT 70.465 10.965 75.810 11.510 ;
        RECT 75.985 10.965 81.330 11.510 ;
        RECT 81.505 10.965 82.715 11.715 ;
        RECT 82.885 10.965 83.175 11.690 ;
        RECT 84.930 11.510 85.270 12.340 ;
        RECT 86.750 11.830 87.100 13.080 ;
        RECT 90.450 11.510 90.790 12.340 ;
        RECT 92.270 11.830 92.620 13.080 ;
        RECT 94.385 12.425 95.595 13.515 ;
        RECT 94.385 11.715 94.905 12.255 ;
        RECT 95.075 11.885 95.595 12.425 ;
        RECT 95.765 12.350 96.055 13.515 ;
        RECT 96.225 13.080 101.570 13.515 ;
        RECT 101.745 13.080 107.090 13.515 ;
        RECT 83.345 10.965 88.690 11.510 ;
        RECT 88.865 10.965 94.210 11.510 ;
        RECT 94.385 10.965 95.595 11.715 ;
        RECT 95.765 10.965 96.055 11.690 ;
        RECT 97.810 11.510 98.150 12.340 ;
        RECT 99.630 11.830 99.980 13.080 ;
        RECT 103.330 11.510 103.670 12.340 ;
        RECT 105.150 11.830 105.500 13.080 ;
        RECT 107.265 12.425 108.475 13.515 ;
        RECT 107.265 11.715 107.785 12.255 ;
        RECT 107.955 11.885 108.475 12.425 ;
        RECT 108.645 12.350 108.935 13.515 ;
        RECT 109.105 13.080 114.450 13.515 ;
        RECT 96.225 10.965 101.570 11.510 ;
        RECT 101.745 10.965 107.090 11.510 ;
        RECT 107.265 10.965 108.475 11.715 ;
        RECT 108.645 10.965 108.935 11.690 ;
        RECT 110.690 11.510 111.030 12.340 ;
        RECT 112.510 11.830 112.860 13.080 ;
        RECT 114.625 12.425 117.215 13.515 ;
        RECT 114.625 11.735 115.835 12.255 ;
        RECT 116.005 11.905 117.215 12.425 ;
        RECT 117.385 12.425 118.595 13.515 ;
        RECT 117.385 11.885 117.905 12.425 ;
        RECT 109.105 10.965 114.450 11.510 ;
        RECT 114.625 10.965 117.215 11.735 ;
        RECT 118.075 11.715 118.595 12.255 ;
        RECT 117.385 10.965 118.595 11.715 ;
        RECT 5.520 10.795 118.680 10.965 ;
      LAYER met1 ;
        RECT 5.520 122.160 118.680 122.640 ;
        RECT 32.695 121.620 32.985 121.665 ;
        RECT 34.585 121.620 34.875 121.665 ;
        RECT 37.705 121.620 37.995 121.665 ;
        RECT 32.695 121.480 37.995 121.620 ;
        RECT 32.695 121.435 32.985 121.480 ;
        RECT 34.585 121.435 34.875 121.480 ;
        RECT 37.705 121.435 37.995 121.480 ;
        RECT 98.935 121.620 99.225 121.665 ;
        RECT 100.825 121.620 101.115 121.665 ;
        RECT 103.945 121.620 104.235 121.665 ;
        RECT 98.935 121.480 104.235 121.620 ;
        RECT 98.935 121.435 99.225 121.480 ;
        RECT 100.825 121.435 101.115 121.480 ;
        RECT 103.945 121.435 104.235 121.480 ;
        RECT 31.825 121.280 32.115 121.325 ;
        RECT 33.650 121.280 33.970 121.340 ;
        RECT 31.825 121.140 33.970 121.280 ;
        RECT 31.825 121.095 32.115 121.140 ;
        RECT 33.650 121.080 33.970 121.140 ;
        RECT 35.030 121.280 35.350 121.340 ;
        RECT 41.945 121.280 42.235 121.325 ;
        RECT 35.030 121.140 42.235 121.280 ;
        RECT 35.030 121.080 35.350 121.140 ;
        RECT 41.945 121.095 42.235 121.140 ;
        RECT 106.790 121.280 107.110 121.340 ;
        RECT 108.185 121.280 108.475 121.325 ;
        RECT 106.790 121.140 108.475 121.280 ;
        RECT 106.790 121.080 107.110 121.140 ;
        RECT 108.185 121.095 108.475 121.140 ;
        RECT 13.410 120.740 13.730 121.000 ;
        RECT 32.290 120.940 32.580 120.985 ;
        RECT 34.125 120.940 34.415 120.985 ;
        RECT 37.705 120.940 37.995 120.985 ;
        RECT 32.290 120.800 37.995 120.940 ;
        RECT 32.290 120.755 32.580 120.800 ;
        RECT 34.125 120.755 34.415 120.800 ;
        RECT 37.705 120.755 37.995 120.800 ;
        RECT 33.190 120.400 33.510 120.660 ;
        RECT 35.490 120.645 35.810 120.660 ;
        RECT 38.785 120.645 39.075 120.960 ;
        RECT 96.210 120.940 96.530 121.000 ;
        RECT 98.065 120.940 98.355 120.985 ;
        RECT 96.210 120.800 98.355 120.940 ;
        RECT 96.210 120.740 96.530 120.800 ;
        RECT 98.065 120.755 98.355 120.800 ;
        RECT 98.530 120.940 98.820 120.985 ;
        RECT 100.365 120.940 100.655 120.985 ;
        RECT 103.945 120.940 104.235 120.985 ;
        RECT 98.530 120.800 104.235 120.940 ;
        RECT 98.530 120.755 98.820 120.800 ;
        RECT 100.365 120.755 100.655 120.800 ;
        RECT 103.945 120.755 104.235 120.800 ;
        RECT 104.950 120.960 105.270 121.000 ;
        RECT 104.950 120.740 105.315 120.960 ;
        RECT 35.485 120.600 36.135 120.645 ;
        RECT 38.785 120.600 39.375 120.645 ;
        RECT 35.485 120.460 39.375 120.600 ;
        RECT 35.485 120.415 36.135 120.460 ;
        RECT 39.085 120.415 39.375 120.460 ;
        RECT 98.970 120.600 99.290 120.660 ;
        RECT 105.025 120.645 105.315 120.740 ;
        RECT 99.445 120.600 99.735 120.645 ;
        RECT 98.970 120.460 99.735 120.600 ;
        RECT 35.490 120.400 35.810 120.415 ;
        RECT 98.970 120.400 99.290 120.460 ;
        RECT 99.445 120.415 99.735 120.460 ;
        RECT 101.725 120.600 102.375 120.645 ;
        RECT 105.025 120.600 105.615 120.645 ;
        RECT 101.725 120.460 105.615 120.600 ;
        RECT 101.725 120.415 102.375 120.460 ;
        RECT 105.325 120.415 105.615 120.460 ;
        RECT 12.950 120.060 13.270 120.320 ;
        RECT 5.520 119.440 118.680 119.920 ;
        RECT 88.850 119.240 89.170 119.300 ;
        RECT 88.850 119.100 93.680 119.240 ;
        RECT 88.850 119.040 89.170 119.100 ;
        RECT 16.630 118.945 16.950 118.960 ;
        RECT 13.065 118.900 13.355 118.945 ;
        RECT 16.305 118.900 16.955 118.945 ;
        RECT 13.065 118.760 16.955 118.900 ;
        RECT 13.065 118.715 13.655 118.760 ;
        RECT 16.305 118.715 16.955 118.760 ;
        RECT 24.445 118.900 25.095 118.945 ;
        RECT 28.045 118.900 28.335 118.945 ;
        RECT 28.590 118.900 28.910 118.960 ;
        RECT 24.445 118.760 28.910 118.900 ;
        RECT 24.445 118.715 25.095 118.760 ;
        RECT 27.745 118.715 28.335 118.760 ;
        RECT 6.970 118.360 7.290 118.620 ;
        RECT 13.365 118.400 13.655 118.715 ;
        RECT 16.630 118.700 16.950 118.715 ;
        RECT 14.445 118.560 14.735 118.605 ;
        RECT 18.025 118.560 18.315 118.605 ;
        RECT 19.860 118.560 20.150 118.605 ;
        RECT 14.445 118.420 20.150 118.560 ;
        RECT 14.445 118.375 14.735 118.420 ;
        RECT 18.025 118.375 18.315 118.420 ;
        RECT 19.860 118.375 20.150 118.420 ;
        RECT 21.250 118.560 21.540 118.605 ;
        RECT 23.085 118.560 23.375 118.605 ;
        RECT 26.665 118.560 26.955 118.605 ;
        RECT 21.250 118.420 26.955 118.560 ;
        RECT 21.250 118.375 21.540 118.420 ;
        RECT 23.085 118.375 23.375 118.420 ;
        RECT 26.665 118.375 26.955 118.420 ;
        RECT 27.745 118.400 28.035 118.715 ;
        RECT 28.590 118.700 28.910 118.760 ;
        RECT 29.050 118.900 29.370 118.960 ;
        RECT 30.905 118.900 31.195 118.945 ;
        RECT 29.050 118.760 31.195 118.900 ;
        RECT 29.050 118.700 29.370 118.760 ;
        RECT 30.905 118.715 31.195 118.760 ;
        RECT 39.625 118.900 40.275 118.945 ;
        RECT 43.225 118.900 43.515 118.945 ;
        RECT 45.150 118.900 45.470 118.960 ;
        RECT 39.625 118.760 45.470 118.900 ;
        RECT 39.625 118.715 40.275 118.760 ;
        RECT 42.925 118.715 43.515 118.760 ;
        RECT 36.430 118.560 36.720 118.605 ;
        RECT 38.265 118.560 38.555 118.605 ;
        RECT 41.845 118.560 42.135 118.605 ;
        RECT 36.430 118.420 42.135 118.560 ;
        RECT 36.430 118.375 36.720 118.420 ;
        RECT 38.265 118.375 38.555 118.420 ;
        RECT 41.845 118.375 42.135 118.420 ;
        RECT 42.925 118.400 43.215 118.715 ;
        RECT 45.150 118.700 45.470 118.760 ;
        RECT 46.070 118.700 46.390 118.960 ;
        RECT 50.205 118.900 50.855 118.945 ;
        RECT 53.805 118.900 54.095 118.945 ;
        RECT 50.205 118.760 54.095 118.900 ;
        RECT 50.205 118.715 50.855 118.760 ;
        RECT 53.505 118.715 54.095 118.760 ;
        RECT 56.665 118.900 56.955 118.945 ;
        RECT 58.950 118.900 59.270 118.960 ;
        RECT 56.665 118.760 59.270 118.900 ;
        RECT 56.665 118.715 56.955 118.760 ;
        RECT 53.505 118.620 53.795 118.715 ;
        RECT 58.950 118.700 59.270 118.760 ;
        RECT 63.085 118.900 63.735 118.945 ;
        RECT 66.685 118.900 66.975 118.945 ;
        RECT 68.610 118.900 68.930 118.960 ;
        RECT 63.085 118.760 68.930 118.900 ;
        RECT 63.085 118.715 63.735 118.760 ;
        RECT 66.385 118.715 66.975 118.760 ;
        RECT 47.010 118.560 47.300 118.605 ;
        RECT 48.845 118.560 49.135 118.605 ;
        RECT 52.425 118.560 52.715 118.605 ;
        RECT 47.010 118.420 52.715 118.560 ;
        RECT 47.010 118.375 47.300 118.420 ;
        RECT 48.845 118.375 49.135 118.420 ;
        RECT 52.425 118.375 52.715 118.420 ;
        RECT 53.430 118.400 53.795 118.620 ;
        RECT 59.890 118.560 60.180 118.605 ;
        RECT 61.725 118.560 62.015 118.605 ;
        RECT 65.305 118.560 65.595 118.605 ;
        RECT 59.890 118.420 65.595 118.560 ;
        RECT 53.430 118.360 53.750 118.400 ;
        RECT 59.890 118.375 60.180 118.420 ;
        RECT 61.725 118.375 62.015 118.420 ;
        RECT 65.305 118.375 65.595 118.420 ;
        RECT 66.385 118.400 66.675 118.715 ;
        RECT 68.610 118.700 68.930 118.760 ;
        RECT 69.545 118.900 69.835 118.945 ;
        RECT 71.830 118.900 72.150 118.960 ;
        RECT 69.545 118.760 72.150 118.900 ;
        RECT 69.545 118.715 69.835 118.760 ;
        RECT 71.830 118.700 72.150 118.760 ;
        RECT 73.665 118.900 74.315 118.945 ;
        RECT 76.430 118.900 76.750 118.960 ;
        RECT 77.265 118.900 77.555 118.945 ;
        RECT 73.665 118.760 77.555 118.900 ;
        RECT 73.665 118.715 74.315 118.760 ;
        RECT 76.430 118.700 76.750 118.760 ;
        RECT 76.965 118.715 77.555 118.760 ;
        RECT 78.270 118.900 78.590 118.960 ;
        RECT 80.125 118.900 80.415 118.945 ;
        RECT 78.270 118.760 80.415 118.900 ;
        RECT 70.470 118.560 70.760 118.605 ;
        RECT 72.305 118.560 72.595 118.605 ;
        RECT 75.885 118.560 76.175 118.605 ;
        RECT 70.470 118.420 76.175 118.560 ;
        RECT 70.470 118.375 70.760 118.420 ;
        RECT 72.305 118.375 72.595 118.420 ;
        RECT 75.885 118.375 76.175 118.420 ;
        RECT 76.965 118.400 77.255 118.715 ;
        RECT 78.270 118.700 78.590 118.760 ;
        RECT 80.125 118.715 80.415 118.760 ;
        RECT 87.005 118.900 87.655 118.945 ;
        RECT 89.770 118.900 90.090 118.960 ;
        RECT 93.540 118.945 93.680 119.100 ;
        RECT 104.950 119.040 105.270 119.300 ;
        RECT 90.605 118.900 90.895 118.945 ;
        RECT 87.005 118.760 90.895 118.900 ;
        RECT 87.005 118.715 87.655 118.760 ;
        RECT 89.770 118.700 90.090 118.760 ;
        RECT 90.305 118.715 90.895 118.760 ;
        RECT 93.465 118.715 93.755 118.945 ;
        RECT 80.570 118.360 80.890 118.620 ;
        RECT 83.810 118.560 84.100 118.605 ;
        RECT 85.645 118.560 85.935 118.605 ;
        RECT 89.225 118.560 89.515 118.605 ;
        RECT 83.810 118.420 89.515 118.560 ;
        RECT 83.810 118.375 84.100 118.420 ;
        RECT 85.645 118.375 85.935 118.420 ;
        RECT 89.225 118.375 89.515 118.420 ;
        RECT 90.305 118.400 90.595 118.715 ;
        RECT 93.910 118.700 94.230 118.960 ;
        RECT 96.785 118.900 97.075 118.945 ;
        RECT 100.025 118.900 100.675 118.945 ;
        RECT 96.785 118.760 100.675 118.900 ;
        RECT 96.785 118.715 97.375 118.760 ;
        RECT 100.025 118.715 100.675 118.760 ;
        RECT 97.085 118.400 97.375 118.715 ;
        RECT 98.165 118.560 98.455 118.605 ;
        RECT 101.745 118.560 102.035 118.605 ;
        RECT 103.580 118.560 103.870 118.605 ;
        RECT 98.165 118.420 103.870 118.560 ;
        RECT 10.205 118.220 10.495 118.265 ;
        RECT 17.090 118.220 17.410 118.280 ;
        RECT 10.205 118.080 17.410 118.220 ;
        RECT 10.205 118.035 10.495 118.080 ;
        RECT 17.090 118.020 17.410 118.080 ;
        RECT 18.930 118.020 19.250 118.280 ;
        RECT 20.325 118.220 20.615 118.265 ;
        RECT 20.770 118.220 21.090 118.280 ;
        RECT 20.325 118.080 21.090 118.220 ;
        RECT 20.325 118.035 20.615 118.080 ;
        RECT 20.770 118.020 21.090 118.080 ;
        RECT 22.150 118.020 22.470 118.280 ;
        RECT 33.650 118.220 33.970 118.280 ;
        RECT 35.965 118.220 36.255 118.265 ;
        RECT 33.650 118.080 36.255 118.220 ;
        RECT 33.650 118.020 33.970 118.080 ;
        RECT 35.965 118.035 36.255 118.080 ;
        RECT 37.345 118.220 37.635 118.265 ;
        RECT 44.690 118.220 45.010 118.280 ;
        RECT 37.345 118.080 45.010 118.220 ;
        RECT 37.345 118.035 37.635 118.080 ;
        RECT 44.690 118.020 45.010 118.080 ;
        RECT 46.530 118.020 46.850 118.280 ;
        RECT 47.925 118.220 48.215 118.265 ;
        RECT 57.110 118.220 57.430 118.280 ;
        RECT 47.925 118.080 57.430 118.220 ;
        RECT 47.925 118.035 48.215 118.080 ;
        RECT 57.110 118.020 57.430 118.080 ;
        RECT 59.410 118.020 59.730 118.280 ;
        RECT 60.805 118.220 61.095 118.265 ;
        RECT 69.070 118.220 69.390 118.280 ;
        RECT 60.805 118.080 69.390 118.220 ;
        RECT 60.805 118.035 61.095 118.080 ;
        RECT 69.070 118.020 69.390 118.080 ;
        RECT 70.005 118.035 70.295 118.265 ;
        RECT 71.385 118.220 71.675 118.265 ;
        RECT 75.050 118.220 75.370 118.280 ;
        RECT 83.345 118.220 83.635 118.265 ;
        RECT 71.385 118.080 75.370 118.220 ;
        RECT 71.385 118.035 71.675 118.080 ;
        RECT 14.445 117.880 14.735 117.925 ;
        RECT 17.565 117.880 17.855 117.925 ;
        RECT 19.455 117.880 19.745 117.925 ;
        RECT 14.445 117.740 19.745 117.880 ;
        RECT 14.445 117.695 14.735 117.740 ;
        RECT 17.565 117.695 17.855 117.740 ;
        RECT 19.455 117.695 19.745 117.740 ;
        RECT 21.655 117.880 21.945 117.925 ;
        RECT 23.545 117.880 23.835 117.925 ;
        RECT 26.665 117.880 26.955 117.925 ;
        RECT 21.655 117.740 26.955 117.880 ;
        RECT 21.655 117.695 21.945 117.740 ;
        RECT 23.545 117.695 23.835 117.740 ;
        RECT 26.665 117.695 26.955 117.740 ;
        RECT 36.835 117.880 37.125 117.925 ;
        RECT 38.725 117.880 39.015 117.925 ;
        RECT 41.845 117.880 42.135 117.925 ;
        RECT 36.835 117.740 42.135 117.880 ;
        RECT 36.835 117.695 37.125 117.740 ;
        RECT 38.725 117.695 39.015 117.740 ;
        RECT 41.845 117.695 42.135 117.740 ;
        RECT 47.415 117.880 47.705 117.925 ;
        RECT 49.305 117.880 49.595 117.925 ;
        RECT 52.425 117.880 52.715 117.925 ;
        RECT 47.415 117.740 52.715 117.880 ;
        RECT 47.415 117.695 47.705 117.740 ;
        RECT 49.305 117.695 49.595 117.740 ;
        RECT 52.425 117.695 52.715 117.740 ;
        RECT 60.295 117.880 60.585 117.925 ;
        RECT 62.185 117.880 62.475 117.925 ;
        RECT 65.305 117.880 65.595 117.925 ;
        RECT 60.295 117.740 65.595 117.880 ;
        RECT 60.295 117.695 60.585 117.740 ;
        RECT 62.185 117.695 62.475 117.740 ;
        RECT 65.305 117.695 65.595 117.740 ;
        RECT 7.905 117.540 8.195 117.585 ;
        RECT 53.890 117.540 54.210 117.600 ;
        RECT 7.905 117.400 54.210 117.540 ;
        RECT 7.905 117.355 8.195 117.400 ;
        RECT 53.890 117.340 54.210 117.400 ;
        RECT 59.410 117.540 59.730 117.600 ;
        RECT 70.080 117.540 70.220 118.035 ;
        RECT 75.050 118.020 75.370 118.080 ;
        RECT 82.730 118.080 83.635 118.220 ;
        RECT 82.730 117.940 82.870 118.080 ;
        RECT 83.345 118.035 83.635 118.080 ;
        RECT 84.710 118.020 85.030 118.280 ;
        RECT 96.670 118.220 96.990 118.280 ;
        RECT 97.220 118.220 97.360 118.400 ;
        RECT 98.165 118.375 98.455 118.420 ;
        RECT 101.745 118.375 102.035 118.420 ;
        RECT 103.580 118.375 103.870 118.420 ;
        RECT 105.410 118.360 105.730 118.620 ;
        RECT 96.670 118.080 97.360 118.220 ;
        RECT 97.590 118.220 97.910 118.280 ;
        RECT 102.665 118.220 102.955 118.265 ;
        RECT 97.590 118.080 102.955 118.220 ;
        RECT 96.670 118.020 96.990 118.080 ;
        RECT 97.590 118.020 97.910 118.080 ;
        RECT 102.665 118.035 102.955 118.080 ;
        RECT 104.045 118.035 104.335 118.265 ;
        RECT 70.875 117.880 71.165 117.925 ;
        RECT 72.765 117.880 73.055 117.925 ;
        RECT 75.885 117.880 76.175 117.925 ;
        RECT 82.410 117.880 82.870 117.940 ;
        RECT 70.875 117.740 76.175 117.880 ;
        RECT 70.875 117.695 71.165 117.740 ;
        RECT 72.765 117.695 73.055 117.740 ;
        RECT 75.885 117.695 76.175 117.740 ;
        RECT 76.520 117.740 82.870 117.880 ;
        RECT 84.215 117.880 84.505 117.925 ;
        RECT 86.105 117.880 86.395 117.925 ;
        RECT 89.225 117.880 89.515 117.925 ;
        RECT 84.215 117.740 89.515 117.880 ;
        RECT 76.520 117.600 76.660 117.740 ;
        RECT 82.410 117.680 82.730 117.740 ;
        RECT 84.215 117.695 84.505 117.740 ;
        RECT 86.105 117.695 86.395 117.740 ;
        RECT 89.225 117.695 89.515 117.740 ;
        RECT 98.165 117.880 98.455 117.925 ;
        RECT 101.285 117.880 101.575 117.925 ;
        RECT 103.175 117.880 103.465 117.925 ;
        RECT 98.165 117.740 103.465 117.880 ;
        RECT 98.165 117.695 98.455 117.740 ;
        RECT 101.285 117.695 101.575 117.740 ;
        RECT 103.175 117.695 103.465 117.740 ;
        RECT 104.120 117.600 104.260 118.035 ;
        RECT 76.430 117.540 76.750 117.600 ;
        RECT 59.410 117.400 76.750 117.540 ;
        RECT 59.410 117.340 59.730 117.400 ;
        RECT 76.430 117.340 76.750 117.400 ;
        RECT 81.045 117.540 81.335 117.585 ;
        RECT 82.870 117.540 83.190 117.600 ;
        RECT 81.045 117.400 83.190 117.540 ;
        RECT 81.045 117.355 81.335 117.400 ;
        RECT 82.870 117.340 83.190 117.400 ;
        RECT 96.210 117.540 96.530 117.600 ;
        RECT 104.030 117.540 104.350 117.600 ;
        RECT 96.210 117.400 104.350 117.540 ;
        RECT 96.210 117.340 96.530 117.400 ;
        RECT 104.030 117.340 104.350 117.400 ;
        RECT 5.520 116.720 118.680 117.200 ;
        RECT 28.590 116.520 28.910 116.580 ;
        RECT 29.985 116.520 30.275 116.565 ;
        RECT 28.590 116.380 30.275 116.520 ;
        RECT 28.590 116.320 28.910 116.380 ;
        RECT 29.985 116.335 30.275 116.380 ;
        RECT 32.745 116.520 33.035 116.565 ;
        RECT 35.490 116.520 35.810 116.580 ;
        RECT 32.745 116.380 35.810 116.520 ;
        RECT 32.745 116.335 33.035 116.380 ;
        RECT 35.490 116.320 35.810 116.380 ;
        RECT 44.690 116.320 45.010 116.580 ;
        RECT 57.110 116.320 57.430 116.580 ;
        RECT 69.070 116.520 69.390 116.580 ;
        RECT 70.465 116.520 70.755 116.565 ;
        RECT 69.070 116.380 70.755 116.520 ;
        RECT 69.070 116.320 69.390 116.380 ;
        RECT 70.465 116.335 70.755 116.380 ;
        RECT 75.065 116.520 75.355 116.565 ;
        RECT 75.970 116.520 76.290 116.580 ;
        RECT 75.065 116.380 76.290 116.520 ;
        RECT 75.065 116.335 75.355 116.380 ;
        RECT 75.970 116.320 76.290 116.380 ;
        RECT 84.710 116.520 85.030 116.580 ;
        RECT 86.565 116.520 86.855 116.565 ;
        RECT 84.710 116.380 86.855 116.520 ;
        RECT 84.710 116.320 85.030 116.380 ;
        RECT 86.565 116.335 86.855 116.380 ;
        RECT 88.405 116.520 88.695 116.565 ;
        RECT 89.770 116.520 90.090 116.580 ;
        RECT 88.405 116.380 90.090 116.520 ;
        RECT 88.405 116.335 88.695 116.380 ;
        RECT 89.770 116.320 90.090 116.380 ;
        RECT 93.005 116.520 93.295 116.565 ;
        RECT 96.670 116.520 96.990 116.580 ;
        RECT 93.005 116.380 96.990 116.520 ;
        RECT 93.005 116.335 93.295 116.380 ;
        RECT 96.670 116.320 96.990 116.380 ;
        RECT 11.225 116.180 11.515 116.225 ;
        RECT 14.345 116.180 14.635 116.225 ;
        RECT 16.235 116.180 16.525 116.225 ;
        RECT 11.225 116.040 16.525 116.180 ;
        RECT 11.225 115.995 11.515 116.040 ;
        RECT 14.345 115.995 14.635 116.040 ;
        RECT 16.235 115.995 16.525 116.040 ;
        RECT 19.815 116.180 20.105 116.225 ;
        RECT 21.705 116.180 21.995 116.225 ;
        RECT 24.825 116.180 25.115 116.225 ;
        RECT 19.815 116.040 25.115 116.180 ;
        RECT 19.815 115.995 20.105 116.040 ;
        RECT 21.705 115.995 21.995 116.040 ;
        RECT 24.825 115.995 25.115 116.040 ;
        RECT 34.535 116.180 34.825 116.225 ;
        RECT 36.425 116.180 36.715 116.225 ;
        RECT 39.545 116.180 39.835 116.225 ;
        RECT 34.535 116.040 39.835 116.180 ;
        RECT 34.535 115.995 34.825 116.040 ;
        RECT 36.425 115.995 36.715 116.040 ;
        RECT 39.545 115.995 39.835 116.040 ;
        RECT 47.415 116.180 47.705 116.225 ;
        RECT 49.305 116.180 49.595 116.225 ;
        RECT 52.425 116.180 52.715 116.225 ;
        RECT 47.415 116.040 52.715 116.180 ;
        RECT 47.415 115.995 47.705 116.040 ;
        RECT 49.305 115.995 49.595 116.040 ;
        RECT 52.425 115.995 52.715 116.040 ;
        RECT 60.295 116.180 60.585 116.225 ;
        RECT 62.185 116.180 62.475 116.225 ;
        RECT 65.305 116.180 65.595 116.225 ;
        RECT 60.295 116.040 65.595 116.180 ;
        RECT 60.295 115.995 60.585 116.040 ;
        RECT 62.185 115.995 62.475 116.040 ;
        RECT 65.305 115.995 65.595 116.040 ;
        RECT 68.610 116.180 68.930 116.240 ;
        RECT 72.305 116.180 72.595 116.225 ;
        RECT 76.855 116.180 77.145 116.225 ;
        RECT 78.745 116.180 79.035 116.225 ;
        RECT 81.865 116.180 82.155 116.225 ;
        RECT 68.610 116.040 72.595 116.180 ;
        RECT 68.610 115.980 68.930 116.040 ;
        RECT 72.305 115.995 72.595 116.040 ;
        RECT 74.680 116.040 76.660 116.180 ;
        RECT 6.985 115.840 7.275 115.885 ;
        RECT 12.030 115.840 12.350 115.900 ;
        RECT 6.985 115.700 12.350 115.840 ;
        RECT 6.985 115.655 7.275 115.700 ;
        RECT 12.030 115.640 12.350 115.700 ;
        RECT 17.105 115.840 17.395 115.885 ;
        RECT 18.945 115.840 19.235 115.885 ;
        RECT 20.770 115.840 21.090 115.900 ;
        RECT 33.650 115.840 33.970 115.900 ;
        RECT 46.530 115.840 46.850 115.900 ;
        RECT 17.105 115.700 46.850 115.840 ;
        RECT 17.105 115.655 17.395 115.700 ;
        RECT 18.945 115.655 19.235 115.700 ;
        RECT 20.770 115.640 21.090 115.700 ;
        RECT 33.650 115.640 33.970 115.700 ;
        RECT 46.530 115.640 46.850 115.700 ;
        RECT 52.970 115.840 53.290 115.900 ;
        RECT 56.665 115.840 56.955 115.885 ;
        RECT 52.970 115.700 56.955 115.840 ;
        RECT 52.970 115.640 53.290 115.700 ;
        RECT 56.665 115.655 56.955 115.700 ;
        RECT 59.410 115.640 59.730 115.900 ;
        RECT 64.470 115.840 64.790 115.900 ;
        RECT 69.545 115.840 69.835 115.885 ;
        RECT 64.470 115.700 69.835 115.840 ;
        RECT 64.470 115.640 64.790 115.700 ;
        RECT 69.545 115.655 69.835 115.700 ;
        RECT 10.145 115.205 10.435 115.520 ;
        RECT 11.225 115.500 11.515 115.545 ;
        RECT 14.805 115.500 15.095 115.545 ;
        RECT 16.640 115.500 16.930 115.545 ;
        RECT 11.225 115.360 16.930 115.500 ;
        RECT 11.225 115.315 11.515 115.360 ;
        RECT 14.805 115.315 15.095 115.360 ;
        RECT 16.640 115.315 16.930 115.360 ;
        RECT 19.410 115.500 19.700 115.545 ;
        RECT 21.245 115.500 21.535 115.545 ;
        RECT 24.825 115.500 25.115 115.545 ;
        RECT 19.410 115.360 25.115 115.500 ;
        RECT 19.410 115.315 19.700 115.360 ;
        RECT 21.245 115.315 21.535 115.360 ;
        RECT 24.825 115.315 25.115 115.360 ;
        RECT 9.845 115.160 10.435 115.205 ;
        RECT 12.950 115.205 13.270 115.220 ;
        RECT 12.950 115.160 13.735 115.205 ;
        RECT 9.845 115.020 13.735 115.160 ;
        RECT 9.845 114.975 10.135 115.020 ;
        RECT 12.950 114.975 13.735 115.020 ;
        RECT 12.950 114.960 13.270 114.975 ;
        RECT 15.710 114.960 16.030 115.220 ;
        RECT 20.325 115.160 20.615 115.205 ;
        RECT 21.690 115.160 22.010 115.220 ;
        RECT 20.325 115.020 22.010 115.160 ;
        RECT 20.325 114.975 20.615 115.020 ;
        RECT 21.690 114.960 22.010 115.020 ;
        RECT 22.605 115.160 23.255 115.205 ;
        RECT 23.530 115.160 23.850 115.220 ;
        RECT 25.905 115.205 26.195 115.520 ;
        RECT 30.430 115.500 30.750 115.560 ;
        RECT 32.285 115.500 32.575 115.545 ;
        RECT 30.430 115.360 32.575 115.500 ;
        RECT 30.430 115.300 30.750 115.360 ;
        RECT 32.285 115.315 32.575 115.360 ;
        RECT 34.130 115.500 34.420 115.545 ;
        RECT 35.965 115.500 36.255 115.545 ;
        RECT 39.545 115.500 39.835 115.545 ;
        RECT 34.130 115.360 39.835 115.500 ;
        RECT 34.130 115.315 34.420 115.360 ;
        RECT 35.965 115.315 36.255 115.360 ;
        RECT 39.545 115.315 39.835 115.360 ;
        RECT 25.905 115.160 26.495 115.205 ;
        RECT 22.605 115.020 26.495 115.160 ;
        RECT 22.605 114.975 23.255 115.020 ;
        RECT 23.530 114.960 23.850 115.020 ;
        RECT 26.205 114.975 26.495 115.020 ;
        RECT 29.065 114.975 29.355 115.205 ;
        RECT 23.990 114.820 24.310 114.880 ;
        RECT 29.140 114.820 29.280 114.975 ;
        RECT 35.030 114.960 35.350 115.220 ;
        RECT 37.325 115.160 37.975 115.205 ;
        RECT 40.090 115.160 40.410 115.220 ;
        RECT 40.625 115.205 40.915 115.520 ;
        RECT 45.625 115.500 45.915 115.545 ;
        RECT 46.070 115.500 46.390 115.560 ;
        RECT 45.625 115.360 46.390 115.500 ;
        RECT 45.625 115.315 45.915 115.360 ;
        RECT 46.070 115.300 46.390 115.360 ;
        RECT 47.010 115.500 47.300 115.545 ;
        RECT 48.845 115.500 49.135 115.545 ;
        RECT 52.425 115.500 52.715 115.545 ;
        RECT 47.010 115.360 52.715 115.500 ;
        RECT 47.010 115.315 47.300 115.360 ;
        RECT 48.845 115.315 49.135 115.360 ;
        RECT 52.425 115.315 52.715 115.360 ;
        RECT 40.625 115.160 41.215 115.205 ;
        RECT 37.325 115.020 41.215 115.160 ;
        RECT 37.325 114.975 37.975 115.020 ;
        RECT 40.090 114.960 40.410 115.020 ;
        RECT 40.925 114.975 41.215 115.020 ;
        RECT 43.785 114.975 44.075 115.205 ;
        RECT 47.925 115.160 48.215 115.205 ;
        RECT 49.290 115.160 49.610 115.220 ;
        RECT 47.925 115.020 49.610 115.160 ;
        RECT 47.925 114.975 48.215 115.020 ;
        RECT 23.990 114.680 29.280 114.820 ;
        RECT 39.170 114.820 39.490 114.880 ;
        RECT 43.860 114.820 44.000 114.975 ;
        RECT 49.290 114.960 49.610 115.020 ;
        RECT 50.205 115.160 50.855 115.205 ;
        RECT 51.130 115.160 51.450 115.220 ;
        RECT 53.505 115.205 53.795 115.520 ;
        RECT 58.030 115.300 58.350 115.560 ;
        RECT 59.890 115.500 60.180 115.545 ;
        RECT 61.725 115.500 62.015 115.545 ;
        RECT 65.305 115.500 65.595 115.545 ;
        RECT 59.890 115.360 65.595 115.500 ;
        RECT 59.890 115.315 60.180 115.360 ;
        RECT 61.725 115.315 62.015 115.360 ;
        RECT 65.305 115.315 65.595 115.360 ;
        RECT 53.505 115.160 54.095 115.205 ;
        RECT 50.205 115.020 54.095 115.160 ;
        RECT 50.205 114.975 50.855 115.020 ;
        RECT 51.130 114.960 51.450 115.020 ;
        RECT 53.805 114.975 54.095 115.020 ;
        RECT 60.790 114.960 61.110 115.220 ;
        RECT 66.385 115.205 66.675 115.520 ;
        RECT 71.385 115.500 71.675 115.545 ;
        RECT 72.290 115.500 72.610 115.560 ;
        RECT 71.385 115.360 72.610 115.500 ;
        RECT 71.385 115.315 71.675 115.360 ;
        RECT 72.290 115.300 72.610 115.360 ;
        RECT 72.750 115.500 73.070 115.560 ;
        RECT 74.680 115.545 74.820 116.040 ;
        RECT 75.970 115.640 76.290 115.900 ;
        RECT 76.520 115.840 76.660 116.040 ;
        RECT 76.855 116.040 82.155 116.180 ;
        RECT 76.855 115.995 77.145 116.040 ;
        RECT 78.745 115.995 79.035 116.040 ;
        RECT 81.865 115.995 82.155 116.040 ;
        RECT 82.730 116.040 88.160 116.180 ;
        RECT 80.570 115.840 80.890 115.900 ;
        RECT 82.730 115.840 82.870 116.040 ;
        RECT 76.520 115.700 82.870 115.840 ;
        RECT 83.330 115.840 83.650 115.900 ;
        RECT 86.105 115.840 86.395 115.885 ;
        RECT 83.330 115.700 86.395 115.840 ;
        RECT 80.570 115.640 80.890 115.700 ;
        RECT 83.330 115.640 83.650 115.700 ;
        RECT 86.105 115.655 86.395 115.700 ;
        RECT 74.605 115.500 74.895 115.545 ;
        RECT 72.750 115.360 74.895 115.500 ;
        RECT 72.750 115.300 73.070 115.360 ;
        RECT 74.605 115.315 74.895 115.360 ;
        RECT 76.450 115.500 76.740 115.545 ;
        RECT 78.285 115.500 78.575 115.545 ;
        RECT 81.865 115.500 82.155 115.545 ;
        RECT 76.450 115.360 82.155 115.500 ;
        RECT 76.450 115.315 76.740 115.360 ;
        RECT 78.285 115.315 78.575 115.360 ;
        RECT 81.865 115.315 82.155 115.360 ;
        RECT 82.870 115.520 83.190 115.560 ;
        RECT 82.870 115.300 83.235 115.520 ;
        RECT 87.010 115.500 87.330 115.560 ;
        RECT 88.020 115.545 88.160 116.040 ;
        RECT 90.705 115.995 90.995 116.225 ;
        RECT 97.095 116.180 97.385 116.225 ;
        RECT 98.985 116.180 99.275 116.225 ;
        RECT 102.105 116.180 102.395 116.225 ;
        RECT 97.095 116.040 102.395 116.180 ;
        RECT 97.095 115.995 97.385 116.040 ;
        RECT 98.985 115.995 99.275 116.040 ;
        RECT 102.105 115.995 102.395 116.040 ;
        RECT 107.675 116.180 107.965 116.225 ;
        RECT 109.565 116.180 109.855 116.225 ;
        RECT 112.685 116.180 112.975 116.225 ;
        RECT 107.675 116.040 112.975 116.180 ;
        RECT 107.675 115.995 107.965 116.040 ;
        RECT 109.565 115.995 109.855 116.040 ;
        RECT 112.685 115.995 112.975 116.040 ;
        RECT 90.780 115.840 90.920 115.995 ;
        RECT 97.590 115.840 97.910 115.900 ;
        RECT 90.780 115.700 97.910 115.840 ;
        RECT 97.590 115.640 97.910 115.700 ;
        RECT 102.650 115.840 102.970 115.900 ;
        RECT 104.030 115.840 104.350 115.900 ;
        RECT 106.805 115.840 107.095 115.885 ;
        RECT 102.650 115.700 103.800 115.840 ;
        RECT 102.650 115.640 102.970 115.700 ;
        RECT 87.485 115.500 87.775 115.545 ;
        RECT 87.010 115.360 87.775 115.500 ;
        RECT 87.010 115.300 87.330 115.360 ;
        RECT 87.485 115.315 87.775 115.360 ;
        RECT 87.945 115.315 88.235 115.545 ;
        RECT 89.785 115.500 90.075 115.545 ;
        RECT 91.610 115.500 91.930 115.560 ;
        RECT 92.545 115.500 92.835 115.545 ;
        RECT 89.785 115.360 91.930 115.500 ;
        RECT 89.785 115.315 90.075 115.360 ;
        RECT 63.085 115.160 63.735 115.205 ;
        RECT 66.385 115.160 66.975 115.205 ;
        RECT 67.690 115.160 68.010 115.220 ;
        RECT 63.085 115.020 68.010 115.160 ;
        RECT 63.085 114.975 63.735 115.020 ;
        RECT 66.685 114.975 66.975 115.020 ;
        RECT 67.690 114.960 68.010 115.020 ;
        RECT 77.350 114.960 77.670 115.220 ;
        RECT 82.945 115.205 83.235 115.300 ;
        RECT 79.645 115.160 80.295 115.205 ;
        RECT 82.945 115.160 83.535 115.205 ;
        RECT 79.645 115.020 83.535 115.160 ;
        RECT 88.020 115.160 88.160 115.315 ;
        RECT 91.610 115.300 91.930 115.360 ;
        RECT 92.160 115.360 92.835 115.500 ;
        RECT 92.160 115.220 92.300 115.360 ;
        RECT 92.545 115.315 92.835 115.360 ;
        RECT 94.370 115.300 94.690 115.560 ;
        RECT 96.210 115.300 96.530 115.560 ;
        RECT 96.690 115.500 96.980 115.545 ;
        RECT 98.525 115.500 98.815 115.545 ;
        RECT 102.105 115.500 102.395 115.545 ;
        RECT 96.690 115.360 102.395 115.500 ;
        RECT 96.690 115.315 96.980 115.360 ;
        RECT 98.525 115.315 98.815 115.360 ;
        RECT 102.105 115.315 102.395 115.360 ;
        RECT 92.070 115.160 92.390 115.220 ;
        RECT 97.605 115.160 97.895 115.205 ;
        RECT 88.020 115.020 92.390 115.160 ;
        RECT 79.645 114.975 80.295 115.020 ;
        RECT 83.245 114.975 83.535 115.020 ;
        RECT 92.070 114.960 92.390 115.020 ;
        RECT 95.380 115.020 97.895 115.160 ;
        RECT 95.380 114.865 95.520 115.020 ;
        RECT 97.605 114.975 97.895 115.020 ;
        RECT 99.885 115.160 100.535 115.205 ;
        RECT 101.270 115.160 101.590 115.220 ;
        RECT 103.185 115.205 103.475 115.520 ;
        RECT 103.660 115.500 103.800 115.700 ;
        RECT 104.030 115.700 107.095 115.840 ;
        RECT 104.030 115.640 104.350 115.700 ;
        RECT 106.805 115.655 107.095 115.700 ;
        RECT 114.150 115.840 114.470 115.900 ;
        RECT 116.925 115.840 117.215 115.885 ;
        RECT 114.150 115.700 117.215 115.840 ;
        RECT 114.150 115.640 114.470 115.700 ;
        RECT 116.925 115.655 117.215 115.700 ;
        RECT 106.345 115.500 106.635 115.545 ;
        RECT 103.660 115.360 106.635 115.500 ;
        RECT 106.345 115.315 106.635 115.360 ;
        RECT 107.270 115.500 107.560 115.545 ;
        RECT 109.105 115.500 109.395 115.545 ;
        RECT 112.685 115.500 112.975 115.545 ;
        RECT 107.270 115.360 112.975 115.500 ;
        RECT 107.270 115.315 107.560 115.360 ;
        RECT 109.105 115.315 109.395 115.360 ;
        RECT 112.685 115.315 112.975 115.360 ;
        RECT 103.185 115.160 103.775 115.205 ;
        RECT 99.885 115.020 103.775 115.160 ;
        RECT 99.885 114.975 100.535 115.020 ;
        RECT 101.270 114.960 101.590 115.020 ;
        RECT 103.485 114.975 103.775 115.020 ;
        RECT 108.185 114.975 108.475 115.205 ;
        RECT 109.550 115.160 109.870 115.220 ;
        RECT 113.765 115.205 114.055 115.520 ;
        RECT 110.465 115.160 111.115 115.205 ;
        RECT 113.765 115.160 114.355 115.205 ;
        RECT 109.550 115.020 114.355 115.160 ;
        RECT 39.170 114.680 44.000 114.820 ;
        RECT 23.990 114.620 24.310 114.680 ;
        RECT 39.170 114.620 39.490 114.680 ;
        RECT 95.305 114.635 95.595 114.865 ;
        RECT 100.810 114.820 101.130 114.880 ;
        RECT 108.260 114.820 108.400 114.975 ;
        RECT 109.550 114.960 109.870 115.020 ;
        RECT 110.465 114.975 111.115 115.020 ;
        RECT 114.065 114.975 114.355 115.020 ;
        RECT 100.810 114.680 108.400 114.820 ;
        RECT 100.810 114.620 101.130 114.680 ;
        RECT 5.520 114.000 118.680 114.480 ;
        RECT 13.870 113.600 14.190 113.860 ;
        RECT 16.630 113.800 16.950 113.860 ;
        RECT 18.025 113.800 18.315 113.845 ;
        RECT 16.630 113.660 18.315 113.800 ;
        RECT 16.630 113.600 16.950 113.660 ;
        RECT 18.025 113.615 18.315 113.660 ;
        RECT 18.930 113.800 19.250 113.860 ;
        RECT 20.325 113.800 20.615 113.845 ;
        RECT 18.930 113.660 20.615 113.800 ;
        RECT 18.930 113.600 19.250 113.660 ;
        RECT 20.325 113.615 20.615 113.660 ;
        RECT 21.690 113.600 22.010 113.860 ;
        RECT 23.530 113.600 23.850 113.860 ;
        RECT 32.745 113.800 33.035 113.845 ;
        RECT 33.190 113.800 33.510 113.860 ;
        RECT 32.745 113.660 33.510 113.800 ;
        RECT 32.745 113.615 33.035 113.660 ;
        RECT 33.190 113.600 33.510 113.660 ;
        RECT 35.030 113.800 35.350 113.860 ;
        RECT 38.265 113.800 38.555 113.845 ;
        RECT 35.030 113.660 38.555 113.800 ;
        RECT 35.030 113.600 35.350 113.660 ;
        RECT 38.265 113.615 38.555 113.660 ;
        RECT 40.090 113.600 40.410 113.860 ;
        RECT 45.150 113.600 45.470 113.860 ;
        RECT 49.290 113.600 49.610 113.860 ;
        RECT 53.430 113.800 53.750 113.860 ;
        RECT 56.205 113.800 56.495 113.845 ;
        RECT 53.430 113.660 56.495 113.800 ;
        RECT 53.430 113.600 53.750 113.660 ;
        RECT 56.205 113.615 56.495 113.660 ;
        RECT 60.790 113.800 61.110 113.860 ;
        RECT 63.565 113.800 63.855 113.845 ;
        RECT 60.790 113.660 63.855 113.800 ;
        RECT 60.790 113.600 61.110 113.660 ;
        RECT 63.565 113.615 63.855 113.660 ;
        RECT 67.690 113.600 68.010 113.860 ;
        RECT 75.050 113.600 75.370 113.860 ;
        RECT 77.350 113.800 77.670 113.860 ;
        RECT 81.045 113.800 81.335 113.845 ;
        RECT 77.350 113.660 81.335 113.800 ;
        RECT 77.350 113.600 77.670 113.660 ;
        RECT 81.045 113.615 81.335 113.660 ;
        RECT 98.525 113.800 98.815 113.845 ;
        RECT 98.970 113.800 99.290 113.860 ;
        RECT 98.525 113.660 99.290 113.800 ;
        RECT 98.525 113.615 98.815 113.660 ;
        RECT 98.970 113.600 99.290 113.660 ;
        RECT 100.810 113.600 101.130 113.860 ;
        RECT 101.270 113.800 101.590 113.860 ;
        RECT 101.745 113.800 102.035 113.845 ;
        RECT 101.270 113.660 102.035 113.800 ;
        RECT 101.270 113.600 101.590 113.660 ;
        RECT 101.745 113.615 102.035 113.660 ;
        RECT 109.550 113.600 109.870 113.860 ;
        RECT 5.130 113.460 5.450 113.520 ;
        RECT 12.950 113.505 13.270 113.520 ;
        RECT 6.985 113.460 7.275 113.505 ;
        RECT 5.130 113.320 7.275 113.460 ;
        RECT 5.130 113.260 5.450 113.320 ;
        RECT 6.985 113.275 7.275 113.320 ;
        RECT 9.845 113.460 10.135 113.505 ;
        RECT 12.950 113.460 13.735 113.505 ;
        RECT 9.845 113.320 13.735 113.460 ;
        RECT 13.960 113.460 14.100 113.600 ;
        RECT 30.430 113.460 30.750 113.520 ;
        RECT 57.110 113.460 57.430 113.520 ;
        RECT 13.960 113.320 40.780 113.460 ;
        RECT 9.845 113.275 10.435 113.320 ;
        RECT 10.145 112.960 10.435 113.275 ;
        RECT 12.950 113.275 13.735 113.320 ;
        RECT 12.950 113.260 13.270 113.275 ;
        RECT 18.560 113.165 18.700 113.320 ;
        RECT 11.225 113.120 11.515 113.165 ;
        RECT 14.805 113.120 15.095 113.165 ;
        RECT 16.640 113.120 16.930 113.165 ;
        RECT 11.225 112.980 16.930 113.120 ;
        RECT 11.225 112.935 11.515 112.980 ;
        RECT 14.805 112.935 15.095 112.980 ;
        RECT 16.640 112.935 16.930 112.980 ;
        RECT 18.485 112.935 18.775 113.165 ;
        RECT 21.245 113.120 21.535 113.165 ;
        RECT 21.690 113.120 22.010 113.180 ;
        RECT 21.245 112.980 22.010 113.120 ;
        RECT 21.245 112.935 21.535 112.980 ;
        RECT 21.690 112.920 22.010 112.980 ;
        RECT 22.610 112.920 22.930 113.180 ;
        RECT 23.160 113.165 23.300 113.320 ;
        RECT 30.430 113.260 30.750 113.320 ;
        RECT 23.085 112.935 23.375 113.165 ;
        RECT 26.765 113.120 27.055 113.165 ;
        RECT 29.510 113.120 29.830 113.180 ;
        RECT 26.765 112.980 29.830 113.120 ;
        RECT 26.765 112.935 27.055 112.980 ;
        RECT 29.510 112.920 29.830 112.980 ;
        RECT 31.825 113.120 32.115 113.165 ;
        RECT 33.190 113.120 33.510 113.180 ;
        RECT 31.825 112.980 33.510 113.120 ;
        RECT 31.825 112.935 32.115 112.980 ;
        RECT 33.190 112.920 33.510 112.980 ;
        RECT 38.250 113.120 38.570 113.180 ;
        RECT 40.640 113.165 40.780 113.320 ;
        RECT 50.300 113.320 57.430 113.460 ;
        RECT 50.300 113.165 50.440 113.320 ;
        RECT 57.110 113.260 57.430 113.320 ;
        RECT 92.070 113.460 92.390 113.520 ;
        RECT 105.410 113.460 105.730 113.520 ;
        RECT 92.070 113.320 109.320 113.460 ;
        RECT 92.070 113.260 92.390 113.320 ;
        RECT 39.185 113.120 39.475 113.165 ;
        RECT 38.250 112.980 39.475 113.120 ;
        RECT 38.250 112.920 38.570 112.980 ;
        RECT 39.185 112.935 39.475 112.980 ;
        RECT 40.565 113.120 40.855 113.165 ;
        RECT 45.625 113.120 45.915 113.165 ;
        RECT 40.565 112.980 45.915 113.120 ;
        RECT 40.565 112.935 40.855 112.980 ;
        RECT 45.625 112.935 45.915 112.980 ;
        RECT 50.225 112.935 50.515 113.165 ;
        RECT 52.985 113.120 53.275 113.165 ;
        RECT 53.890 113.120 54.210 113.180 ;
        RECT 54.365 113.120 54.655 113.165 ;
        RECT 52.985 112.980 53.660 113.120 ;
        RECT 52.985 112.935 53.275 112.980 ;
        RECT 13.870 112.780 14.190 112.840 ;
        RECT 15.725 112.780 16.015 112.825 ;
        RECT 13.870 112.640 16.015 112.780 ;
        RECT 13.870 112.580 14.190 112.640 ;
        RECT 15.725 112.595 16.015 112.640 ;
        RECT 17.105 112.780 17.395 112.825 ;
        RECT 45.700 112.780 45.840 112.935 ;
        RECT 51.590 112.780 51.910 112.840 ;
        RECT 17.105 112.640 21.460 112.780 ;
        RECT 45.700 112.640 51.910 112.780 ;
        RECT 53.520 112.780 53.660 112.980 ;
        RECT 53.890 112.980 54.655 113.120 ;
        RECT 53.890 112.920 54.210 112.980 ;
        RECT 54.365 112.935 54.655 112.980 ;
        RECT 54.810 113.120 55.130 113.180 ;
        RECT 55.745 113.120 56.035 113.165 ;
        RECT 54.810 112.980 56.035 113.120 ;
        RECT 54.810 112.920 55.130 112.980 ;
        RECT 55.745 112.935 56.035 112.980 ;
        RECT 64.010 113.120 64.330 113.180 ;
        RECT 64.485 113.120 64.775 113.165 ;
        RECT 64.010 112.980 64.775 113.120 ;
        RECT 64.010 112.920 64.330 112.980 ;
        RECT 64.485 112.935 64.775 112.980 ;
        RECT 68.165 113.120 68.455 113.165 ;
        RECT 71.845 113.120 72.135 113.165 ;
        RECT 72.750 113.120 73.070 113.180 ;
        RECT 68.165 112.980 73.070 113.120 ;
        RECT 68.165 112.935 68.455 112.980 ;
        RECT 71.845 112.935 72.135 112.980 ;
        RECT 72.750 112.920 73.070 112.980 ;
        RECT 73.210 112.920 73.530 113.180 ;
        RECT 75.970 112.920 76.290 113.180 ;
        RECT 81.030 113.120 81.350 113.180 ;
        RECT 81.965 113.120 82.255 113.165 ;
        RECT 81.030 112.980 82.255 113.120 ;
        RECT 81.030 112.920 81.350 112.980 ;
        RECT 81.965 112.935 82.255 112.980 ;
        RECT 97.605 113.120 97.895 113.165 ;
        RECT 98.510 113.120 98.830 113.180 ;
        RECT 101.360 113.165 101.500 113.320 ;
        RECT 105.410 113.260 105.730 113.320 ;
        RECT 97.605 112.980 98.830 113.120 ;
        RECT 97.605 112.935 97.895 112.980 ;
        RECT 98.510 112.920 98.830 112.980 ;
        RECT 99.905 112.935 100.195 113.165 ;
        RECT 101.285 112.935 101.575 113.165 ;
        RECT 103.570 113.120 103.890 113.180 ;
        RECT 109.180 113.165 109.320 113.320 ;
        RECT 104.505 113.120 104.795 113.165 ;
        RECT 103.570 112.980 104.795 113.120 ;
        RECT 73.300 112.780 73.440 112.920 ;
        RECT 53.520 112.640 73.440 112.780 ;
        RECT 99.980 112.780 100.120 112.935 ;
        RECT 103.570 112.920 103.890 112.980 ;
        RECT 104.505 112.935 104.795 112.980 ;
        RECT 109.105 113.120 109.395 113.165 ;
        RECT 111.405 113.120 111.695 113.165 ;
        RECT 109.105 112.980 111.695 113.120 ;
        RECT 109.105 112.935 109.395 112.980 ;
        RECT 111.405 112.935 111.695 112.980 ;
        RECT 101.730 112.780 102.050 112.840 ;
        RECT 99.980 112.640 102.050 112.780 ;
        RECT 17.105 112.595 17.395 112.640 ;
        RECT 21.320 112.500 21.460 112.640 ;
        RECT 51.590 112.580 51.910 112.640 ;
        RECT 101.730 112.580 102.050 112.640 ;
        RECT 11.225 112.440 11.515 112.485 ;
        RECT 14.345 112.440 14.635 112.485 ;
        RECT 16.235 112.440 16.525 112.485 ;
        RECT 11.225 112.300 16.525 112.440 ;
        RECT 11.225 112.255 11.515 112.300 ;
        RECT 14.345 112.255 14.635 112.300 ;
        RECT 16.235 112.255 16.525 112.300 ;
        RECT 21.230 112.240 21.550 112.500 ;
        RECT 22.150 112.440 22.470 112.500 ;
        RECT 25.845 112.440 26.135 112.485 ;
        RECT 22.150 112.300 26.135 112.440 ;
        RECT 22.150 112.240 22.470 112.300 ;
        RECT 25.845 112.255 26.135 112.300 ;
        RECT 54.825 112.100 55.115 112.145 ;
        RECT 58.950 112.100 59.270 112.160 ;
        RECT 54.825 111.960 59.270 112.100 ;
        RECT 54.825 111.915 55.115 111.960 ;
        RECT 58.950 111.900 59.270 111.960 ;
        RECT 105.410 111.900 105.730 112.160 ;
        RECT 111.850 111.900 112.170 112.160 ;
        RECT 5.520 111.280 118.680 111.760 ;
        RECT 105.410 111.080 105.730 111.140 ;
        RECT 108.090 111.080 108.380 111.125 ;
        RECT 105.410 110.940 108.380 111.080 ;
        RECT 105.410 110.880 105.730 110.940 ;
        RECT 108.090 110.895 108.380 110.940 ;
        RECT 92.545 110.740 92.835 110.785 ;
        RECT 96.210 110.740 96.530 110.800 ;
        RECT 107.675 110.740 107.965 110.785 ;
        RECT 109.565 110.740 109.855 110.785 ;
        RECT 112.685 110.740 112.975 110.785 ;
        RECT 12.580 110.600 13.640 110.740 ;
        RECT 12.580 110.400 12.720 110.600 ;
        RECT 9.820 110.260 12.720 110.400 ;
        RECT 9.820 110.105 9.960 110.260 ;
        RECT 12.950 110.200 13.270 110.460 ;
        RECT 13.500 110.400 13.640 110.600 ;
        RECT 89.860 110.600 107.020 110.740 ;
        RECT 28.590 110.400 28.910 110.460 ;
        RECT 13.500 110.260 28.910 110.400 ;
        RECT 28.590 110.200 28.910 110.260 ;
        RECT 51.130 110.400 51.450 110.460 ;
        RECT 52.065 110.400 52.355 110.445 ;
        RECT 51.130 110.260 52.355 110.400 ;
        RECT 51.130 110.200 51.450 110.260 ;
        RECT 52.065 110.215 52.355 110.260 ;
        RECT 82.410 110.400 82.730 110.460 ;
        RECT 89.860 110.400 90.000 110.600 ;
        RECT 92.545 110.555 92.835 110.600 ;
        RECT 96.210 110.540 96.530 110.600 ;
        RECT 82.410 110.260 90.000 110.400 ;
        RECT 82.410 110.200 82.730 110.260 ;
        RECT 106.880 110.120 107.020 110.600 ;
        RECT 107.675 110.600 112.975 110.740 ;
        RECT 107.675 110.555 107.965 110.600 ;
        RECT 109.565 110.555 109.855 110.600 ;
        RECT 112.685 110.555 112.975 110.600 ;
        RECT 116.925 110.400 117.215 110.445 ;
        RECT 118.750 110.400 119.070 110.460 ;
        RECT 116.925 110.260 119.070 110.400 ;
        RECT 116.925 110.215 117.215 110.260 ;
        RECT 118.750 110.200 119.070 110.260 ;
        RECT 9.745 109.875 10.035 110.105 ;
        RECT 11.110 109.860 11.430 110.120 ;
        RECT 13.410 109.860 13.730 110.120 ;
        RECT 51.590 110.060 51.910 110.120 ;
        RECT 54.810 110.060 55.130 110.120 ;
        RECT 51.590 109.920 55.130 110.060 ;
        RECT 51.590 109.860 51.910 109.920 ;
        RECT 54.810 109.860 55.130 109.920 ;
        RECT 97.130 110.060 97.450 110.120 ;
        RECT 98.065 110.060 98.355 110.105 ;
        RECT 97.130 109.920 98.355 110.060 ;
        RECT 97.130 109.860 97.450 109.920 ;
        RECT 98.065 109.875 98.355 109.920 ;
        RECT 106.790 109.860 107.110 110.120 ;
        RECT 107.270 110.060 107.560 110.105 ;
        RECT 109.105 110.060 109.395 110.105 ;
        RECT 112.685 110.060 112.975 110.105 ;
        RECT 107.270 109.920 112.975 110.060 ;
        RECT 107.270 109.875 107.560 109.920 ;
        RECT 109.105 109.875 109.395 109.920 ;
        RECT 112.685 109.875 112.975 109.920 ;
        RECT 13.870 109.720 14.190 109.780 ;
        RECT 31.365 109.720 31.655 109.765 ;
        RECT 10.740 109.580 14.190 109.720 ;
        RECT 10.740 109.425 10.880 109.580 ;
        RECT 13.870 109.520 14.190 109.580 ;
        RECT 30.060 109.580 31.655 109.720 ;
        RECT 10.665 109.195 10.955 109.425 ;
        RECT 12.045 109.380 12.335 109.425 ;
        RECT 15.710 109.380 16.030 109.440 ;
        RECT 12.045 109.240 16.030 109.380 ;
        RECT 12.045 109.195 12.335 109.240 ;
        RECT 15.710 109.180 16.030 109.240 ;
        RECT 21.230 109.380 21.550 109.440 ;
        RECT 30.060 109.425 30.200 109.580 ;
        RECT 31.365 109.535 31.655 109.580 ;
        RECT 40.090 109.520 40.410 109.780 ;
        RECT 83.790 109.720 84.110 109.780 ;
        RECT 86.105 109.720 86.395 109.765 ;
        RECT 83.790 109.580 86.395 109.720 ;
        RECT 83.790 109.520 84.110 109.580 ;
        RECT 86.105 109.535 86.395 109.580 ;
        RECT 110.465 109.720 111.115 109.765 ;
        RECT 111.850 109.720 112.170 109.780 ;
        RECT 113.765 109.765 114.055 110.080 ;
        RECT 113.765 109.720 114.355 109.765 ;
        RECT 110.465 109.580 114.355 109.720 ;
        RECT 110.465 109.535 111.115 109.580 ;
        RECT 111.850 109.520 112.170 109.580 ;
        RECT 114.065 109.535 114.355 109.580 ;
        RECT 29.985 109.380 30.275 109.425 ;
        RECT 21.230 109.240 30.275 109.380 ;
        RECT 21.230 109.180 21.550 109.240 ;
        RECT 29.985 109.195 30.275 109.240 ;
        RECT 98.050 109.380 98.370 109.440 ;
        RECT 98.525 109.380 98.815 109.425 ;
        RECT 98.050 109.240 98.815 109.380 ;
        RECT 98.050 109.180 98.370 109.240 ;
        RECT 98.525 109.195 98.815 109.240 ;
        RECT 5.520 108.560 118.680 109.040 ;
        RECT 11.110 108.360 11.430 108.420 ;
        RECT 31.350 108.360 31.670 108.420 ;
        RECT 11.110 108.220 31.670 108.360 ;
        RECT 11.110 108.160 11.430 108.220 ;
        RECT 31.350 108.160 31.670 108.220 ;
        RECT 97.130 108.360 97.450 108.420 ;
        RECT 97.130 108.220 109.320 108.360 ;
        RECT 97.130 108.160 97.450 108.220 ;
        RECT 41.930 108.065 42.250 108.080 ;
        RECT 50.210 108.065 50.530 108.080 ;
        RECT 38.660 108.020 38.950 108.065 ;
        RECT 41.920 108.020 42.250 108.065 ;
        RECT 38.660 107.880 42.250 108.020 ;
        RECT 38.660 107.835 38.950 107.880 ;
        RECT 41.920 107.835 42.250 107.880 ;
        RECT 41.930 107.820 42.250 107.835 ;
        RECT 42.840 108.020 43.130 108.065 ;
        RECT 44.700 108.020 44.990 108.065 ;
        RECT 42.840 107.880 44.990 108.020 ;
        RECT 42.840 107.835 43.130 107.880 ;
        RECT 44.700 107.835 44.990 107.880 ;
        RECT 47.470 108.020 47.760 108.065 ;
        RECT 49.330 108.020 49.620 108.065 ;
        RECT 47.470 107.880 49.620 108.020 ;
        RECT 47.470 107.835 47.760 107.880 ;
        RECT 49.330 107.835 49.620 107.880 ;
        RECT 19.865 107.680 20.155 107.725 ;
        RECT 23.530 107.680 23.850 107.740 ;
        RECT 19.865 107.540 23.850 107.680 ;
        RECT 19.865 107.495 20.155 107.540 ;
        RECT 23.530 107.480 23.850 107.540 ;
        RECT 23.990 107.680 24.310 107.740 ;
        RECT 24.925 107.680 25.215 107.725 ;
        RECT 23.990 107.540 25.215 107.680 ;
        RECT 23.990 107.480 24.310 107.540 ;
        RECT 24.925 107.495 25.215 107.540 ;
        RECT 31.810 107.480 32.130 107.740 ;
        RECT 40.520 107.680 40.810 107.725 ;
        RECT 42.840 107.680 43.055 107.835 ;
        RECT 40.520 107.540 43.055 107.680 ;
        RECT 49.405 107.680 49.620 107.835 ;
        RECT 50.210 108.020 50.540 108.065 ;
        RECT 53.510 108.020 53.800 108.065 ;
        RECT 50.210 107.880 53.800 108.020 ;
        RECT 50.210 107.835 50.540 107.880 ;
        RECT 53.510 107.835 53.800 107.880 ;
        RECT 85.645 108.020 85.935 108.065 ;
        RECT 90.690 108.020 91.010 108.080 ;
        RECT 104.490 108.065 104.810 108.080 ;
        RECT 85.645 107.880 91.010 108.020 ;
        RECT 85.645 107.835 85.935 107.880 ;
        RECT 50.210 107.820 50.530 107.835 ;
        RECT 90.690 107.820 91.010 107.880 ;
        RECT 101.220 108.020 101.510 108.065 ;
        RECT 104.480 108.020 104.810 108.065 ;
        RECT 101.220 107.880 104.810 108.020 ;
        RECT 101.220 107.835 101.510 107.880 ;
        RECT 104.480 107.835 104.810 107.880 ;
        RECT 104.490 107.820 104.810 107.835 ;
        RECT 105.400 108.020 105.690 108.065 ;
        RECT 107.260 108.020 107.550 108.065 ;
        RECT 105.400 107.880 107.550 108.020 ;
        RECT 105.400 107.835 105.690 107.880 ;
        RECT 107.260 107.835 107.550 107.880 ;
        RECT 51.650 107.680 51.940 107.725 ;
        RECT 49.405 107.540 51.940 107.680 ;
        RECT 40.520 107.495 40.810 107.540 ;
        RECT 51.650 107.495 51.940 107.540 ;
        RECT 64.930 107.480 65.250 107.740 ;
        RECT 66.785 107.495 67.075 107.725 ;
        RECT 80.585 107.680 80.875 107.725 ;
        RECT 83.330 107.680 83.650 107.740 ;
        RECT 87.945 107.680 88.235 107.725 ;
        RECT 80.585 107.540 83.650 107.680 ;
        RECT 80.585 107.495 80.875 107.540 ;
        RECT 20.310 107.140 20.630 107.400 ;
        RECT 20.785 107.155 21.075 107.385 ;
        RECT 43.785 107.340 44.075 107.385 ;
        RECT 44.690 107.340 45.010 107.400 ;
        RECT 43.785 107.200 45.010 107.340 ;
        RECT 43.785 107.155 44.075 107.200 ;
        RECT 19.850 107.000 20.170 107.060 ;
        RECT 20.860 107.000 21.000 107.155 ;
        RECT 44.690 107.140 45.010 107.200 ;
        RECT 45.625 107.340 45.915 107.385 ;
        RECT 46.530 107.340 46.850 107.400 ;
        RECT 47.450 107.340 47.770 107.400 ;
        RECT 45.625 107.200 47.770 107.340 ;
        RECT 45.625 107.155 45.915 107.200 ;
        RECT 46.530 107.140 46.850 107.200 ;
        RECT 47.450 107.140 47.770 107.200 ;
        RECT 48.370 107.140 48.690 107.400 ;
        RECT 63.550 107.340 63.870 107.400 ;
        RECT 66.860 107.340 67.000 107.495 ;
        RECT 83.330 107.480 83.650 107.540 ;
        RECT 83.880 107.540 88.235 107.680 ;
        RECT 63.550 107.200 67.000 107.340 ;
        RECT 82.870 107.340 83.190 107.400 ;
        RECT 83.880 107.340 84.020 107.540 ;
        RECT 87.945 107.495 88.235 107.540 ;
        RECT 82.870 107.200 84.020 107.340 ;
        RECT 63.550 107.140 63.870 107.200 ;
        RECT 82.870 107.140 83.190 107.200 ;
        RECT 84.725 107.155 85.015 107.385 ;
        RECT 85.185 107.340 85.475 107.385 ;
        RECT 87.010 107.340 87.330 107.400 ;
        RECT 85.185 107.200 87.330 107.340 ;
        RECT 88.020 107.340 88.160 107.495 ;
        RECT 92.990 107.480 93.310 107.740 ;
        RECT 96.210 107.480 96.530 107.740 ;
        RECT 97.130 107.480 97.450 107.740 ;
        RECT 103.080 107.680 103.370 107.725 ;
        RECT 105.400 107.680 105.615 107.835 ;
        RECT 103.080 107.540 105.615 107.680 ;
        RECT 106.345 107.680 106.635 107.725 ;
        RECT 109.180 107.680 109.320 108.220 ;
        RECT 109.565 107.680 109.855 107.725 ;
        RECT 106.345 107.540 108.860 107.680 ;
        RECT 109.180 107.540 111.620 107.680 ;
        RECT 103.080 107.495 103.370 107.540 ;
        RECT 106.345 107.495 106.635 107.540 ;
        RECT 97.220 107.340 97.360 107.480 ;
        RECT 88.020 107.200 97.360 107.340 ;
        RECT 107.250 107.340 107.570 107.400 ;
        RECT 108.185 107.340 108.475 107.385 ;
        RECT 107.250 107.200 108.475 107.340 ;
        RECT 108.720 107.340 108.860 107.540 ;
        RECT 109.565 107.495 109.855 107.540 ;
        RECT 111.480 107.340 111.620 107.540 ;
        RECT 111.850 107.480 112.170 107.740 ;
        RECT 113.230 107.340 113.550 107.400 ;
        RECT 108.720 107.200 111.160 107.340 ;
        RECT 111.480 107.200 113.550 107.340 ;
        RECT 85.185 107.155 85.475 107.200 ;
        RECT 19.850 106.860 21.000 107.000 ;
        RECT 40.520 107.000 40.810 107.045 ;
        RECT 43.300 107.000 43.590 107.045 ;
        RECT 45.160 107.000 45.450 107.045 ;
        RECT 40.520 106.860 45.450 107.000 ;
        RECT 19.850 106.800 20.170 106.860 ;
        RECT 40.520 106.815 40.810 106.860 ;
        RECT 43.300 106.815 43.590 106.860 ;
        RECT 45.160 106.815 45.450 106.860 ;
        RECT 47.010 107.000 47.300 107.045 ;
        RECT 48.870 107.000 49.160 107.045 ;
        RECT 51.650 107.000 51.940 107.045 ;
        RECT 47.010 106.860 51.940 107.000 ;
        RECT 84.800 107.000 84.940 107.155 ;
        RECT 87.010 107.140 87.330 107.200 ;
        RECT 107.250 107.140 107.570 107.200 ;
        RECT 108.185 107.155 108.475 107.200 ;
        RECT 89.310 107.000 89.630 107.060 ;
        RECT 111.020 107.045 111.160 107.200 ;
        RECT 113.230 107.140 113.550 107.200 ;
        RECT 84.800 106.860 89.630 107.000 ;
        RECT 47.010 106.815 47.300 106.860 ;
        RECT 48.870 106.815 49.160 106.860 ;
        RECT 51.650 106.815 51.940 106.860 ;
        RECT 89.310 106.800 89.630 106.860 ;
        RECT 103.080 107.000 103.370 107.045 ;
        RECT 105.860 107.000 106.150 107.045 ;
        RECT 107.720 107.000 108.010 107.045 ;
        RECT 103.080 106.860 108.010 107.000 ;
        RECT 103.080 106.815 103.370 106.860 ;
        RECT 105.860 106.815 106.150 106.860 ;
        RECT 107.720 106.815 108.010 106.860 ;
        RECT 110.945 106.815 111.235 107.045 ;
        RECT 17.550 106.660 17.870 106.720 ;
        RECT 18.025 106.660 18.315 106.705 ;
        RECT 17.550 106.520 18.315 106.660 ;
        RECT 17.550 106.460 17.870 106.520 ;
        RECT 18.025 106.475 18.315 106.520 ;
        RECT 23.070 106.660 23.390 106.720 ;
        RECT 24.005 106.660 24.295 106.705 ;
        RECT 23.070 106.520 24.295 106.660 ;
        RECT 23.070 106.460 23.390 106.520 ;
        RECT 24.005 106.475 24.295 106.520 ;
        RECT 32.730 106.460 33.050 106.720 ;
        RECT 36.655 106.660 36.945 106.705 ;
        RECT 39.170 106.660 39.490 106.720 ;
        RECT 36.655 106.520 39.490 106.660 ;
        RECT 36.655 106.475 36.945 106.520 ;
        RECT 39.170 106.460 39.490 106.520 ;
        RECT 53.430 106.660 53.750 106.720 ;
        RECT 55.515 106.660 55.805 106.705 ;
        RECT 53.430 106.520 55.805 106.660 ;
        RECT 53.430 106.460 53.750 106.520 ;
        RECT 55.515 106.475 55.805 106.520 ;
        RECT 59.410 106.660 59.730 106.720 ;
        RECT 61.710 106.660 62.030 106.720 ;
        RECT 59.410 106.520 62.030 106.660 ;
        RECT 59.410 106.460 59.730 106.520 ;
        RECT 61.710 106.460 62.030 106.520 ;
        RECT 62.170 106.660 62.490 106.720 ;
        RECT 64.025 106.660 64.315 106.705 ;
        RECT 62.170 106.520 64.315 106.660 ;
        RECT 62.170 106.460 62.490 106.520 ;
        RECT 64.025 106.475 64.315 106.520 ;
        RECT 66.310 106.460 66.630 106.720 ;
        RECT 78.270 106.660 78.590 106.720 ;
        RECT 79.665 106.660 79.955 106.705 ;
        RECT 78.270 106.520 79.955 106.660 ;
        RECT 78.270 106.460 78.590 106.520 ;
        RECT 79.665 106.475 79.955 106.520 ;
        RECT 87.470 106.460 87.790 106.720 ;
        RECT 88.405 106.660 88.695 106.705 ;
        RECT 89.770 106.660 90.090 106.720 ;
        RECT 88.405 106.520 90.090 106.660 ;
        RECT 88.405 106.475 88.695 106.520 ;
        RECT 89.770 106.460 90.090 106.520 ;
        RECT 93.910 106.460 94.230 106.720 ;
        RECT 95.290 106.460 95.610 106.720 ;
        RECT 97.590 106.460 97.910 106.720 ;
        RECT 99.215 106.660 99.505 106.705 ;
        RECT 102.190 106.660 102.510 106.720 ;
        RECT 99.215 106.520 102.510 106.660 ;
        RECT 99.215 106.475 99.505 106.520 ;
        RECT 102.190 106.460 102.510 106.520 ;
        RECT 109.550 106.660 109.870 106.720 ;
        RECT 110.025 106.660 110.315 106.705 ;
        RECT 109.550 106.520 110.315 106.660 ;
        RECT 109.550 106.460 109.870 106.520 ;
        RECT 110.025 106.475 110.315 106.520 ;
        RECT 5.520 105.840 118.680 106.320 ;
        RECT 41.930 105.440 42.250 105.700 ;
        RECT 44.690 105.440 45.010 105.700 ;
        RECT 85.415 105.640 85.705 105.685 ;
        RECT 87.010 105.640 87.330 105.700 ;
        RECT 85.415 105.500 87.330 105.640 ;
        RECT 85.415 105.455 85.705 105.500 ;
        RECT 87.010 105.440 87.330 105.500 ;
        RECT 104.490 105.640 104.810 105.700 ;
        RECT 116.005 105.640 116.295 105.685 ;
        RECT 104.490 105.500 116.295 105.640 ;
        RECT 104.490 105.440 104.810 105.500 ;
        RECT 116.005 105.455 116.295 105.500 ;
        RECT 21.710 105.300 22.000 105.345 ;
        RECT 23.570 105.300 23.860 105.345 ;
        RECT 26.350 105.300 26.640 105.345 ;
        RECT 21.710 105.160 26.640 105.300 ;
        RECT 21.710 105.115 22.000 105.160 ;
        RECT 23.570 105.115 23.860 105.160 ;
        RECT 26.350 105.115 26.640 105.160 ;
        RECT 31.370 105.300 31.660 105.345 ;
        RECT 33.230 105.300 33.520 105.345 ;
        RECT 36.010 105.300 36.300 105.345 ;
        RECT 49.290 105.300 49.610 105.360 ;
        RECT 31.370 105.160 36.300 105.300 ;
        RECT 31.370 105.115 31.660 105.160 ;
        RECT 33.230 105.115 33.520 105.160 ;
        RECT 36.010 105.115 36.300 105.160 ;
        RECT 47.080 105.160 49.610 105.300 ;
        RECT 30.905 104.960 31.195 105.005 ;
        RECT 21.320 104.820 31.195 104.960 ;
        RECT 21.320 104.680 21.460 104.820 ;
        RECT 30.905 104.775 31.195 104.820 ;
        RECT 32.730 104.760 33.050 105.020 ;
        RECT 39.170 104.960 39.490 105.020 ;
        RECT 47.080 105.005 47.220 105.160 ;
        RECT 49.290 105.100 49.610 105.160 ;
        RECT 51.150 105.300 51.440 105.345 ;
        RECT 53.010 105.300 53.300 105.345 ;
        RECT 55.790 105.300 56.080 105.345 ;
        RECT 51.150 105.160 56.080 105.300 ;
        RECT 51.150 105.115 51.440 105.160 ;
        RECT 53.010 105.115 53.300 105.160 ;
        RECT 55.790 105.115 56.080 105.160 ;
        RECT 60.810 105.300 61.100 105.345 ;
        RECT 62.670 105.300 62.960 105.345 ;
        RECT 65.450 105.300 65.740 105.345 ;
        RECT 60.810 105.160 65.740 105.300 ;
        RECT 60.810 105.115 61.100 105.160 ;
        RECT 62.670 105.115 62.960 105.160 ;
        RECT 65.450 105.115 65.740 105.160 ;
        RECT 76.910 105.300 77.200 105.345 ;
        RECT 78.770 105.300 79.060 105.345 ;
        RECT 81.550 105.300 81.840 105.345 ;
        RECT 76.910 105.160 81.840 105.300 ;
        RECT 76.910 105.115 77.200 105.160 ;
        RECT 78.770 105.115 79.060 105.160 ;
        RECT 81.550 105.115 81.840 105.160 ;
        RECT 86.570 105.300 86.860 105.345 ;
        RECT 88.430 105.300 88.720 105.345 ;
        RECT 91.210 105.300 91.500 105.345 ;
        RECT 86.570 105.160 91.500 105.300 ;
        RECT 86.570 105.115 86.860 105.160 ;
        RECT 88.430 105.115 88.720 105.160 ;
        RECT 91.210 105.115 91.500 105.160 ;
        RECT 100.320 105.300 100.610 105.345 ;
        RECT 103.100 105.300 103.390 105.345 ;
        RECT 104.960 105.300 105.250 105.345 ;
        RECT 100.320 105.160 105.250 105.300 ;
        RECT 100.320 105.115 100.610 105.160 ;
        RECT 103.100 105.115 103.390 105.160 ;
        RECT 104.960 105.115 105.250 105.160 ;
        RECT 106.350 105.300 106.640 105.345 ;
        RECT 108.210 105.300 108.500 105.345 ;
        RECT 110.990 105.300 111.280 105.345 ;
        RECT 106.350 105.160 111.280 105.300 ;
        RECT 106.350 105.115 106.640 105.160 ;
        RECT 108.210 105.115 108.500 105.160 ;
        RECT 110.990 105.115 111.280 105.160 ;
        RECT 39.170 104.820 46.300 104.960 ;
        RECT 39.170 104.760 39.490 104.820 ;
        RECT 17.550 104.420 17.870 104.680 ;
        RECT 18.945 104.435 19.235 104.665 ;
        RECT 14.790 104.280 15.110 104.340 ;
        RECT 19.020 104.280 19.160 104.435 ;
        RECT 21.230 104.420 21.550 104.680 ;
        RECT 23.070 104.420 23.390 104.680 ;
        RECT 26.350 104.620 26.640 104.665 ;
        RECT 36.010 104.620 36.300 104.665 ;
        RECT 24.105 104.480 26.640 104.620 ;
        RECT 24.105 104.325 24.320 104.480 ;
        RECT 26.350 104.435 26.640 104.480 ;
        RECT 33.765 104.480 36.300 104.620 ;
        RECT 14.790 104.140 19.160 104.280 ;
        RECT 22.170 104.280 22.460 104.325 ;
        RECT 24.030 104.280 24.320 104.325 ;
        RECT 22.170 104.140 24.320 104.280 ;
        RECT 14.790 104.080 15.110 104.140 ;
        RECT 22.170 104.095 22.460 104.140 ;
        RECT 24.030 104.095 24.320 104.140 ;
        RECT 24.950 104.280 25.240 104.325 ;
        RECT 27.210 104.280 27.530 104.340 ;
        RECT 33.765 104.325 33.980 104.480 ;
        RECT 36.010 104.435 36.300 104.480 ;
        RECT 42.405 104.620 42.695 104.665 ;
        RECT 43.785 104.620 44.075 104.665 ;
        RECT 42.405 104.480 44.075 104.620 ;
        RECT 42.405 104.435 42.695 104.480 ;
        RECT 43.785 104.435 44.075 104.480 ;
        RECT 28.210 104.280 28.500 104.325 ;
        RECT 24.950 104.140 28.500 104.280 ;
        RECT 24.950 104.095 25.240 104.140 ;
        RECT 27.210 104.080 27.530 104.140 ;
        RECT 28.210 104.095 28.500 104.140 ;
        RECT 31.830 104.280 32.120 104.325 ;
        RECT 33.690 104.280 33.980 104.325 ;
        RECT 31.830 104.140 33.980 104.280 ;
        RECT 31.830 104.095 32.120 104.140 ;
        RECT 33.690 104.095 33.980 104.140 ;
        RECT 34.610 104.280 34.900 104.325 ;
        RECT 37.870 104.280 38.160 104.325 ;
        RECT 43.325 104.280 43.615 104.325 ;
        RECT 34.610 104.140 43.615 104.280 ;
        RECT 43.860 104.280 44.000 104.435 ;
        RECT 45.610 104.420 45.930 104.680 ;
        RECT 46.160 104.620 46.300 104.820 ;
        RECT 47.005 104.775 47.295 105.005 ;
        RECT 47.450 104.960 47.770 105.020 ;
        RECT 50.685 104.960 50.975 105.005 ;
        RECT 53.430 104.960 53.750 105.020 ;
        RECT 47.450 104.820 50.975 104.960 ;
        RECT 47.450 104.760 47.770 104.820 ;
        RECT 50.685 104.775 50.975 104.820 ;
        RECT 51.680 104.820 53.750 104.960 ;
        RECT 47.925 104.620 48.215 104.665 ;
        RECT 46.160 104.480 48.215 104.620 ;
        RECT 47.925 104.435 48.215 104.480 ;
        RECT 48.385 104.620 48.675 104.665 ;
        RECT 51.680 104.620 51.820 104.820 ;
        RECT 53.430 104.760 53.750 104.820 ;
        RECT 60.345 104.960 60.635 105.005 ;
        RECT 61.710 104.960 62.030 105.020 ;
        RECT 60.345 104.820 62.030 104.960 ;
        RECT 60.345 104.775 60.635 104.820 ;
        RECT 61.710 104.760 62.030 104.820 ;
        RECT 62.170 104.760 62.490 105.020 ;
        RECT 63.550 104.960 63.870 105.020 ;
        RECT 76.430 104.960 76.750 105.020 ;
        RECT 93.910 104.960 94.230 105.020 ;
        RECT 103.585 104.960 103.875 105.005 ;
        RECT 63.550 104.820 71.600 104.960 ;
        RECT 63.550 104.760 63.870 104.820 ;
        RECT 48.385 104.480 51.820 104.620 ;
        RECT 52.050 104.620 52.370 104.680 ;
        RECT 71.460 104.665 71.600 104.820 ;
        RECT 76.430 104.820 86.320 104.960 ;
        RECT 76.430 104.760 76.750 104.820 ;
        RECT 52.525 104.620 52.815 104.665 ;
        RECT 55.790 104.620 56.080 104.665 ;
        RECT 65.450 104.620 65.740 104.665 ;
        RECT 52.050 104.480 52.815 104.620 ;
        RECT 48.385 104.435 48.675 104.480 ;
        RECT 52.050 104.420 52.370 104.480 ;
        RECT 52.525 104.435 52.815 104.480 ;
        RECT 53.545 104.480 56.080 104.620 ;
        RECT 49.750 104.280 50.070 104.340 ;
        RECT 53.545 104.325 53.760 104.480 ;
        RECT 55.790 104.435 56.080 104.480 ;
        RECT 63.205 104.480 65.740 104.620 ;
        RECT 57.570 104.325 57.890 104.340 ;
        RECT 63.205 104.325 63.420 104.480 ;
        RECT 65.450 104.435 65.740 104.480 ;
        RECT 71.385 104.620 71.675 104.665 ;
        RECT 73.210 104.620 73.530 104.680 ;
        RECT 75.050 104.620 75.370 104.680 ;
        RECT 71.385 104.480 75.370 104.620 ;
        RECT 71.385 104.435 71.675 104.480 ;
        RECT 73.210 104.420 73.530 104.480 ;
        RECT 75.050 104.420 75.370 104.480 ;
        RECT 78.270 104.420 78.590 104.680 ;
        RECT 86.180 104.665 86.320 104.820 ;
        RECT 93.910 104.820 103.875 104.960 ;
        RECT 93.910 104.760 94.230 104.820 ;
        RECT 103.585 104.775 103.875 104.820 ;
        RECT 105.425 104.960 105.715 105.005 ;
        RECT 105.885 104.960 106.175 105.005 ;
        RECT 107.250 104.960 107.570 105.020 ;
        RECT 105.425 104.820 107.570 104.960 ;
        RECT 105.425 104.775 105.715 104.820 ;
        RECT 105.885 104.775 106.175 104.820 ;
        RECT 107.250 104.760 107.570 104.820 ;
        RECT 81.550 104.620 81.840 104.665 ;
        RECT 79.305 104.480 81.840 104.620 ;
        RECT 43.860 104.140 50.070 104.280 ;
        RECT 34.610 104.095 34.900 104.140 ;
        RECT 37.870 104.095 38.160 104.140 ;
        RECT 43.325 104.095 43.615 104.140 ;
        RECT 49.750 104.080 50.070 104.140 ;
        RECT 51.610 104.280 51.900 104.325 ;
        RECT 53.470 104.280 53.760 104.325 ;
        RECT 51.610 104.140 53.760 104.280 ;
        RECT 51.610 104.095 51.900 104.140 ;
        RECT 53.470 104.095 53.760 104.140 ;
        RECT 54.390 104.280 54.680 104.325 ;
        RECT 57.570 104.280 57.940 104.325 ;
        RECT 54.390 104.140 57.940 104.280 ;
        RECT 54.390 104.095 54.680 104.140 ;
        RECT 57.570 104.095 57.940 104.140 ;
        RECT 61.270 104.280 61.560 104.325 ;
        RECT 63.130 104.280 63.420 104.325 ;
        RECT 61.270 104.140 63.420 104.280 ;
        RECT 61.270 104.095 61.560 104.140 ;
        RECT 63.130 104.095 63.420 104.140 ;
        RECT 64.050 104.280 64.340 104.325 ;
        RECT 66.310 104.280 66.630 104.340 ;
        RECT 79.305 104.325 79.520 104.480 ;
        RECT 81.550 104.435 81.840 104.480 ;
        RECT 86.105 104.620 86.395 104.665 ;
        RECT 86.550 104.620 86.870 104.680 ;
        RECT 86.105 104.480 86.870 104.620 ;
        RECT 86.105 104.435 86.395 104.480 ;
        RECT 86.550 104.420 86.870 104.480 ;
        RECT 87.930 104.420 88.250 104.680 ;
        RECT 91.210 104.620 91.500 104.665 ;
        RECT 88.965 104.480 91.500 104.620 ;
        RECT 67.310 104.280 67.600 104.325 ;
        RECT 64.050 104.140 67.600 104.280 ;
        RECT 64.050 104.095 64.340 104.140 ;
        RECT 57.570 104.080 57.890 104.095 ;
        RECT 66.310 104.080 66.630 104.140 ;
        RECT 67.310 104.095 67.600 104.140 ;
        RECT 77.370 104.280 77.660 104.325 ;
        RECT 79.230 104.280 79.520 104.325 ;
        RECT 77.370 104.140 79.520 104.280 ;
        RECT 77.370 104.095 77.660 104.140 ;
        RECT 79.230 104.095 79.520 104.140 ;
        RECT 80.150 104.280 80.440 104.325 ;
        RECT 81.950 104.280 82.270 104.340 ;
        RECT 88.965 104.325 89.180 104.480 ;
        RECT 91.210 104.435 91.500 104.480 ;
        RECT 100.320 104.620 100.610 104.665 ;
        RECT 100.320 104.480 102.855 104.620 ;
        RECT 100.320 104.435 100.610 104.480 ;
        RECT 83.410 104.280 83.700 104.325 ;
        RECT 80.150 104.140 83.700 104.280 ;
        RECT 80.150 104.095 80.440 104.140 ;
        RECT 81.950 104.080 82.270 104.140 ;
        RECT 83.410 104.095 83.700 104.140 ;
        RECT 87.030 104.280 87.320 104.325 ;
        RECT 88.890 104.280 89.180 104.325 ;
        RECT 87.030 104.140 89.180 104.280 ;
        RECT 87.030 104.095 87.320 104.140 ;
        RECT 88.890 104.095 89.180 104.140 ;
        RECT 89.770 104.325 90.090 104.340 ;
        RECT 89.770 104.280 90.100 104.325 ;
        RECT 93.070 104.280 93.360 104.325 ;
        RECT 89.770 104.140 93.360 104.280 ;
        RECT 89.770 104.095 90.100 104.140 ;
        RECT 93.070 104.095 93.360 104.140 ;
        RECT 97.590 104.280 97.910 104.340 ;
        RECT 102.640 104.325 102.855 104.480 ;
        RECT 107.710 104.420 108.030 104.680 ;
        RECT 110.990 104.620 111.280 104.665 ;
        RECT 108.745 104.480 111.280 104.620 ;
        RECT 108.745 104.325 108.960 104.480 ;
        RECT 110.990 104.435 111.280 104.480 ;
        RECT 113.690 104.620 114.010 104.680 ;
        RECT 115.545 104.620 115.835 104.665 ;
        RECT 113.690 104.480 115.835 104.620 ;
        RECT 113.690 104.420 114.010 104.480 ;
        RECT 115.545 104.435 115.835 104.480 ;
        RECT 98.460 104.280 98.750 104.325 ;
        RECT 101.720 104.280 102.010 104.325 ;
        RECT 97.590 104.140 102.010 104.280 ;
        RECT 89.770 104.080 90.090 104.095 ;
        RECT 97.590 104.080 97.910 104.140 ;
        RECT 98.460 104.095 98.750 104.140 ;
        RECT 101.720 104.095 102.010 104.140 ;
        RECT 102.640 104.280 102.930 104.325 ;
        RECT 104.500 104.280 104.790 104.325 ;
        RECT 102.640 104.140 104.790 104.280 ;
        RECT 102.640 104.095 102.930 104.140 ;
        RECT 104.500 104.095 104.790 104.140 ;
        RECT 106.810 104.280 107.100 104.325 ;
        RECT 108.670 104.280 108.960 104.325 ;
        RECT 106.810 104.140 108.960 104.280 ;
        RECT 106.810 104.095 107.100 104.140 ;
        RECT 108.670 104.095 108.960 104.140 ;
        RECT 109.550 104.325 109.870 104.340 ;
        RECT 109.550 104.280 109.880 104.325 ;
        RECT 112.850 104.280 113.140 104.325 ;
        RECT 109.550 104.140 113.140 104.280 ;
        RECT 109.550 104.095 109.880 104.140 ;
        RECT 112.850 104.095 113.140 104.140 ;
        RECT 109.550 104.080 109.870 104.095 ;
        RECT 16.630 103.740 16.950 104.000 ;
        RECT 19.390 103.740 19.710 104.000 ;
        RECT 30.430 103.985 30.750 104.000 ;
        RECT 30.215 103.755 30.750 103.985 ;
        RECT 30.430 103.740 30.750 103.755 ;
        RECT 39.630 103.985 39.950 104.000 ;
        RECT 39.630 103.755 40.165 103.985 ;
        RECT 48.830 103.940 49.150 104.000 ;
        RECT 50.225 103.940 50.515 103.985 ;
        RECT 48.830 103.800 50.515 103.940 ;
        RECT 39.630 103.740 39.950 103.755 ;
        RECT 48.830 103.740 49.150 103.800 ;
        RECT 50.225 103.755 50.515 103.800 ;
        RECT 53.890 103.940 54.210 104.000 ;
        RECT 59.655 103.940 59.945 103.985 ;
        RECT 53.890 103.800 59.945 103.940 ;
        RECT 53.890 103.740 54.210 103.800 ;
        RECT 59.655 103.755 59.945 103.800 ;
        RECT 68.610 103.940 68.930 104.000 ;
        RECT 69.315 103.940 69.605 103.985 ;
        RECT 68.610 103.800 69.605 103.940 ;
        RECT 68.610 103.740 68.930 103.800 ;
        RECT 69.315 103.755 69.605 103.800 ;
        RECT 70.910 103.740 71.230 104.000 ;
        RECT 90.690 103.940 91.010 104.000 ;
        RECT 96.670 103.985 96.990 104.000 ;
        RECT 95.075 103.940 95.365 103.985 ;
        RECT 90.690 103.800 95.365 103.940 ;
        RECT 90.690 103.740 91.010 103.800 ;
        RECT 95.075 103.755 95.365 103.800 ;
        RECT 96.455 103.755 96.990 103.985 ;
        RECT 96.670 103.740 96.990 103.755 ;
        RECT 110.470 103.940 110.790 104.000 ;
        RECT 114.855 103.940 115.145 103.985 ;
        RECT 110.470 103.800 115.145 103.940 ;
        RECT 110.470 103.740 110.790 103.800 ;
        RECT 114.855 103.755 115.145 103.800 ;
        RECT 5.520 103.120 118.680 103.600 ;
        RECT 21.230 102.920 21.550 102.980 ;
        RECT 14.880 102.780 21.550 102.920 ;
        RECT 12.490 102.040 12.810 102.300 ;
        RECT 14.330 102.040 14.650 102.300 ;
        RECT 14.880 102.285 15.020 102.780 ;
        RECT 21.230 102.720 21.550 102.780 ;
        RECT 23.990 102.920 24.310 102.980 ;
        RECT 24.465 102.920 24.755 102.965 ;
        RECT 23.990 102.780 24.755 102.920 ;
        RECT 23.990 102.720 24.310 102.780 ;
        RECT 24.465 102.735 24.755 102.780 ;
        RECT 27.210 102.920 27.530 102.980 ;
        RECT 29.065 102.920 29.355 102.965 ;
        RECT 27.210 102.780 29.355 102.920 ;
        RECT 27.210 102.720 27.530 102.780 ;
        RECT 29.065 102.735 29.355 102.780 ;
        RECT 31.810 102.720 32.130 102.980 ;
        RECT 39.170 102.920 39.490 102.980 ;
        RECT 40.105 102.920 40.395 102.965 ;
        RECT 39.170 102.780 40.395 102.920 ;
        RECT 39.170 102.720 39.490 102.780 ;
        RECT 40.105 102.735 40.395 102.780 ;
        RECT 41.945 102.920 42.235 102.965 ;
        RECT 45.610 102.920 45.930 102.980 ;
        RECT 41.945 102.780 45.930 102.920 ;
        RECT 41.945 102.735 42.235 102.780 ;
        RECT 45.610 102.720 45.930 102.780 ;
        RECT 47.925 102.920 48.215 102.965 ;
        RECT 48.370 102.920 48.690 102.980 ;
        RECT 47.925 102.780 48.690 102.920 ;
        RECT 47.925 102.735 48.215 102.780 ;
        RECT 48.370 102.720 48.690 102.780 ;
        RECT 50.210 102.720 50.530 102.980 ;
        RECT 52.050 102.720 52.370 102.980 ;
        RECT 52.525 102.735 52.815 102.965 ;
        RECT 53.890 102.920 54.210 102.980 ;
        RECT 54.365 102.920 54.655 102.965 ;
        RECT 53.890 102.780 54.655 102.920 ;
        RECT 15.730 102.580 16.020 102.625 ;
        RECT 17.590 102.580 17.880 102.625 ;
        RECT 15.730 102.440 17.880 102.580 ;
        RECT 15.730 102.395 16.020 102.440 ;
        RECT 17.590 102.395 17.880 102.440 ;
        RECT 18.510 102.580 18.800 102.625 ;
        RECT 19.390 102.580 19.710 102.640 ;
        RECT 21.770 102.580 22.060 102.625 ;
        RECT 18.510 102.440 22.060 102.580 ;
        RECT 18.510 102.395 18.800 102.440 ;
        RECT 14.805 102.055 15.095 102.285 ;
        RECT 16.630 102.040 16.950 102.300 ;
        RECT 17.665 102.240 17.880 102.395 ;
        RECT 19.390 102.380 19.710 102.440 ;
        RECT 21.770 102.395 22.060 102.440 ;
        RECT 26.305 102.580 26.595 102.625 ;
        RECT 26.750 102.580 27.070 102.640 ;
        RECT 30.430 102.580 30.750 102.640 ;
        RECT 34.125 102.580 34.415 102.625 ;
        RECT 26.305 102.440 34.415 102.580 ;
        RECT 26.305 102.395 26.595 102.440 ;
        RECT 26.750 102.380 27.070 102.440 ;
        RECT 30.430 102.380 30.750 102.440 ;
        RECT 34.125 102.395 34.415 102.440 ;
        RECT 19.910 102.240 20.200 102.285 ;
        RECT 29.525 102.240 29.815 102.285 ;
        RECT 32.730 102.240 33.050 102.300 ;
        RECT 17.665 102.100 20.200 102.240 ;
        RECT 19.910 102.055 20.200 102.100 ;
        RECT 23.160 102.100 33.050 102.240 ;
        RECT 14.420 101.900 14.560 102.040 ;
        RECT 23.160 101.900 23.300 102.100 ;
        RECT 29.525 102.055 29.815 102.100 ;
        RECT 32.730 102.040 33.050 102.100 ;
        RECT 33.650 102.240 33.970 102.300 ;
        RECT 39.630 102.240 39.950 102.300 ;
        RECT 33.650 102.100 39.950 102.240 ;
        RECT 33.650 102.040 33.970 102.100 ;
        RECT 39.630 102.040 39.950 102.100 ;
        RECT 48.830 102.040 49.150 102.300 ;
        RECT 49.750 102.040 50.070 102.300 ;
        RECT 51.145 102.240 51.435 102.285 ;
        RECT 52.600 102.240 52.740 102.735 ;
        RECT 53.890 102.720 54.210 102.780 ;
        RECT 54.365 102.735 54.655 102.780 ;
        RECT 57.570 102.920 57.890 102.980 ;
        RECT 58.045 102.920 58.335 102.965 ;
        RECT 57.570 102.780 58.335 102.920 ;
        RECT 57.570 102.720 57.890 102.780 ;
        RECT 58.045 102.735 58.335 102.780 ;
        RECT 81.950 102.720 82.270 102.980 ;
        RECT 83.330 102.720 83.650 102.980 ;
        RECT 87.930 102.920 88.250 102.980 ;
        RECT 88.405 102.920 88.695 102.965 ;
        RECT 87.930 102.780 88.695 102.920 ;
        RECT 87.930 102.720 88.250 102.780 ;
        RECT 88.405 102.735 88.695 102.780 ;
        RECT 90.690 102.720 91.010 102.980 ;
        RECT 92.990 102.720 93.310 102.980 ;
        RECT 106.805 102.920 107.095 102.965 ;
        RECT 107.710 102.920 108.030 102.980 ;
        RECT 106.805 102.780 108.030 102.920 ;
        RECT 106.805 102.735 107.095 102.780 ;
        RECT 107.710 102.720 108.030 102.780 ;
        RECT 111.850 102.920 112.170 102.980 ;
        RECT 112.785 102.920 113.075 102.965 ;
        RECT 111.850 102.780 113.075 102.920 ;
        RECT 111.850 102.720 112.170 102.780 ;
        RECT 112.785 102.735 113.075 102.780 ;
        RECT 53.430 102.580 53.750 102.640 ;
        RECT 54.825 102.580 55.115 102.625 ;
        RECT 53.430 102.440 55.115 102.580 ;
        RECT 53.430 102.380 53.750 102.440 ;
        RECT 54.825 102.395 55.115 102.440 ;
        RECT 62.170 102.580 62.490 102.640 ;
        RECT 65.410 102.580 65.700 102.625 ;
        RECT 67.270 102.580 67.560 102.625 ;
        RECT 62.170 102.440 64.700 102.580 ;
        RECT 62.170 102.380 62.490 102.440 ;
        RECT 51.145 102.100 52.740 102.240 ;
        RECT 58.505 102.240 58.795 102.285 ;
        RECT 59.870 102.240 60.190 102.300 ;
        RECT 58.505 102.100 60.190 102.240 ;
        RECT 51.145 102.055 51.435 102.100 ;
        RECT 58.505 102.055 58.795 102.100 ;
        RECT 59.870 102.040 60.190 102.100 ;
        RECT 63.090 102.040 63.410 102.300 ;
        RECT 64.560 102.285 64.700 102.440 ;
        RECT 65.410 102.440 67.560 102.580 ;
        RECT 65.410 102.395 65.700 102.440 ;
        RECT 67.270 102.395 67.560 102.440 ;
        RECT 68.190 102.580 68.480 102.625 ;
        RECT 70.910 102.580 71.230 102.640 ;
        RECT 71.450 102.580 71.740 102.625 ;
        RECT 68.190 102.440 71.740 102.580 ;
        RECT 68.190 102.395 68.480 102.440 ;
        RECT 64.485 102.055 64.775 102.285 ;
        RECT 67.345 102.240 67.560 102.395 ;
        RECT 70.910 102.380 71.230 102.440 ;
        RECT 71.450 102.395 71.740 102.440 ;
        RECT 86.550 102.580 86.870 102.640 ;
        RECT 94.390 102.580 94.680 102.625 ;
        RECT 96.250 102.580 96.540 102.625 ;
        RECT 86.550 102.440 93.680 102.580 ;
        RECT 86.550 102.380 86.870 102.440 ;
        RECT 69.590 102.240 69.880 102.285 ;
        RECT 67.345 102.100 69.880 102.240 ;
        RECT 69.590 102.055 69.880 102.100 ;
        RECT 75.050 102.240 75.370 102.300 ;
        RECT 77.365 102.240 77.655 102.285 ;
        RECT 75.050 102.100 77.655 102.240 ;
        RECT 75.050 102.040 75.370 102.100 ;
        RECT 77.365 102.055 77.655 102.100 ;
        RECT 78.745 102.240 79.035 102.285 ;
        RECT 82.425 102.240 82.715 102.285 ;
        RECT 82.870 102.240 83.190 102.300 ;
        RECT 78.745 102.100 83.190 102.240 ;
        RECT 78.745 102.055 79.035 102.100 ;
        RECT 82.425 102.055 82.715 102.100 ;
        RECT 82.870 102.040 83.190 102.100 ;
        RECT 85.185 102.240 85.475 102.285 ;
        RECT 85.185 102.100 86.780 102.240 ;
        RECT 85.185 102.055 85.475 102.100 ;
        RECT 86.640 101.960 86.780 102.100 ;
        RECT 87.470 102.040 87.790 102.300 ;
        RECT 91.150 102.040 91.470 102.300 ;
        RECT 93.540 102.285 93.680 102.440 ;
        RECT 94.390 102.440 96.540 102.580 ;
        RECT 94.390 102.395 94.680 102.440 ;
        RECT 96.250 102.395 96.540 102.440 ;
        RECT 97.170 102.580 97.460 102.625 ;
        RECT 98.050 102.580 98.370 102.640 ;
        RECT 100.430 102.580 100.720 102.625 ;
        RECT 97.170 102.440 100.720 102.580 ;
        RECT 97.170 102.395 97.460 102.440 ;
        RECT 93.465 102.055 93.755 102.285 ;
        RECT 95.290 102.040 95.610 102.300 ;
        RECT 96.325 102.240 96.540 102.395 ;
        RECT 98.050 102.380 98.370 102.440 ;
        RECT 100.430 102.395 100.720 102.440 ;
        RECT 102.190 102.580 102.510 102.640 ;
        RECT 110.945 102.580 111.235 102.625 ;
        RECT 102.190 102.440 111.235 102.580 ;
        RECT 102.190 102.380 102.510 102.440 ;
        RECT 110.945 102.395 111.235 102.440 ;
        RECT 98.570 102.240 98.860 102.285 ;
        RECT 96.325 102.100 98.860 102.240 ;
        RECT 98.570 102.055 98.860 102.100 ;
        RECT 14.420 101.760 23.300 101.900 ;
        RECT 23.530 101.945 23.850 101.960 ;
        RECT 23.530 101.900 24.065 101.945 ;
        RECT 26.765 101.900 27.055 101.945 ;
        RECT 23.530 101.760 27.055 101.900 ;
        RECT 23.530 101.715 24.065 101.760 ;
        RECT 26.765 101.715 27.055 101.760 ;
        RECT 27.670 101.900 27.990 101.960 ;
        RECT 35.045 101.900 35.335 101.945 ;
        RECT 39.185 101.900 39.475 101.945 ;
        RECT 49.290 101.900 49.610 101.960 ;
        RECT 53.430 101.900 53.750 101.960 ;
        RECT 55.285 101.900 55.575 101.945 ;
        RECT 66.325 101.900 66.615 101.945 ;
        RECT 27.670 101.760 55.575 101.900 ;
        RECT 23.530 101.700 23.850 101.715 ;
        RECT 27.670 101.700 27.990 101.760 ;
        RECT 35.045 101.715 35.335 101.760 ;
        RECT 39.185 101.715 39.475 101.760 ;
        RECT 49.290 101.700 49.610 101.760 ;
        RECT 53.430 101.700 53.750 101.760 ;
        RECT 55.285 101.715 55.575 101.760 ;
        RECT 64.100 101.760 66.615 101.900 ;
        RECT 64.100 101.605 64.240 101.760 ;
        RECT 66.325 101.715 66.615 101.760 ;
        RECT 85.645 101.715 85.935 101.945 ;
        RECT 15.270 101.560 15.560 101.605 ;
        RECT 17.130 101.560 17.420 101.605 ;
        RECT 19.910 101.560 20.200 101.605 ;
        RECT 15.270 101.420 20.200 101.560 ;
        RECT 15.270 101.375 15.560 101.420 ;
        RECT 17.130 101.375 17.420 101.420 ;
        RECT 19.910 101.375 20.200 101.420 ;
        RECT 64.025 101.375 64.315 101.605 ;
        RECT 64.950 101.560 65.240 101.605 ;
        RECT 66.810 101.560 67.100 101.605 ;
        RECT 69.590 101.560 69.880 101.605 ;
        RECT 64.950 101.420 69.880 101.560 ;
        RECT 85.720 101.560 85.860 101.715 ;
        RECT 86.090 101.700 86.410 101.960 ;
        RECT 86.550 101.700 86.870 101.960 ;
        RECT 89.310 101.900 89.630 101.960 ;
        RECT 89.785 101.900 90.075 101.945 ;
        RECT 97.130 101.900 97.450 101.960 ;
        RECT 102.280 101.900 102.420 102.380 ;
        RECT 105.885 102.240 106.175 102.285 ;
        RECT 106.330 102.240 106.650 102.300 ;
        RECT 105.885 102.100 106.650 102.240 ;
        RECT 105.885 102.055 106.175 102.100 ;
        RECT 106.330 102.040 106.650 102.100 ;
        RECT 89.310 101.760 90.075 101.900 ;
        RECT 89.310 101.700 89.630 101.760 ;
        RECT 89.785 101.715 90.075 101.760 ;
        RECT 90.320 101.760 102.420 101.900 ;
        RECT 90.320 101.560 90.460 101.760 ;
        RECT 97.130 101.700 97.450 101.760 ;
        RECT 110.025 101.715 110.315 101.945 ;
        RECT 85.720 101.420 90.460 101.560 ;
        RECT 93.930 101.560 94.220 101.605 ;
        RECT 95.790 101.560 96.080 101.605 ;
        RECT 98.570 101.560 98.860 101.605 ;
        RECT 93.930 101.420 98.860 101.560 ;
        RECT 110.100 101.560 110.240 101.715 ;
        RECT 110.470 101.700 110.790 101.960 ;
        RECT 110.930 101.560 111.250 101.620 ;
        RECT 110.100 101.420 111.250 101.560 ;
        RECT 64.950 101.375 65.240 101.420 ;
        RECT 66.810 101.375 67.100 101.420 ;
        RECT 69.590 101.375 69.880 101.420 ;
        RECT 93.930 101.375 94.220 101.420 ;
        RECT 95.790 101.375 96.080 101.420 ;
        RECT 98.570 101.375 98.860 101.420 ;
        RECT 110.930 101.360 111.250 101.420 ;
        RECT 11.570 101.020 11.890 101.280 ;
        RECT 13.870 101.020 14.190 101.280 ;
        RECT 72.290 101.220 72.610 101.280 ;
        RECT 73.455 101.220 73.745 101.265 ;
        RECT 72.290 101.080 73.745 101.220 ;
        RECT 72.290 101.020 72.610 101.080 ;
        RECT 73.455 101.035 73.745 101.080 ;
        RECT 75.510 101.020 75.830 101.280 ;
        RECT 98.050 101.220 98.370 101.280 ;
        RECT 102.435 101.220 102.725 101.265 ;
        RECT 98.050 101.080 102.725 101.220 ;
        RECT 98.050 101.020 98.370 101.080 ;
        RECT 102.435 101.035 102.725 101.080 ;
        RECT 5.520 100.400 118.680 100.880 ;
        RECT 12.490 100.200 12.810 100.260 ;
        RECT 18.945 100.200 19.235 100.245 ;
        RECT 12.490 100.060 19.235 100.200 ;
        RECT 12.490 100.000 12.810 100.060 ;
        RECT 18.945 100.015 19.235 100.060 ;
        RECT 64.930 100.200 65.250 100.260 ;
        RECT 65.405 100.200 65.695 100.245 ;
        RECT 64.930 100.060 65.695 100.200 ;
        RECT 64.930 100.000 65.250 100.060 ;
        RECT 65.405 100.015 65.695 100.060 ;
        RECT 96.210 100.000 96.530 100.260 ;
        RECT 106.330 100.000 106.650 100.260 ;
        RECT 8.830 99.860 9.120 99.905 ;
        RECT 10.690 99.860 10.980 99.905 ;
        RECT 13.470 99.860 13.760 99.905 ;
        RECT 8.830 99.720 13.760 99.860 ;
        RECT 8.830 99.675 9.120 99.720 ;
        RECT 10.690 99.675 10.980 99.720 ;
        RECT 13.470 99.675 13.760 99.720 ;
        RECT 71.390 99.860 71.680 99.905 ;
        RECT 73.250 99.860 73.540 99.905 ;
        RECT 76.030 99.860 76.320 99.905 ;
        RECT 71.390 99.720 76.320 99.860 ;
        RECT 71.390 99.675 71.680 99.720 ;
        RECT 73.250 99.675 73.540 99.720 ;
        RECT 76.030 99.675 76.320 99.720 ;
        RECT 86.090 99.860 86.410 99.920 ;
        RECT 87.010 99.860 87.330 99.920 ;
        RECT 89.310 99.860 89.630 99.920 ;
        RECT 86.090 99.720 99.660 99.860 ;
        RECT 86.090 99.660 86.410 99.720 ;
        RECT 87.010 99.660 87.330 99.720 ;
        RECT 89.310 99.660 89.630 99.720 ;
        RECT 10.205 99.520 10.495 99.565 ;
        RECT 11.570 99.520 11.890 99.580 ;
        RECT 10.205 99.380 11.890 99.520 ;
        RECT 10.205 99.335 10.495 99.380 ;
        RECT 11.570 99.320 11.890 99.380 ;
        RECT 19.390 99.520 19.710 99.580 ;
        RECT 22.165 99.520 22.455 99.565 ;
        RECT 27.670 99.520 27.990 99.580 ;
        RECT 19.390 99.380 27.990 99.520 ;
        RECT 19.390 99.320 19.710 99.380 ;
        RECT 22.165 99.335 22.455 99.380 ;
        RECT 27.670 99.320 27.990 99.380 ;
        RECT 68.150 99.320 68.470 99.580 ;
        RECT 91.150 99.520 91.470 99.580 ;
        RECT 96.210 99.520 96.530 99.580 ;
        RECT 99.520 99.565 99.660 99.720 ;
        RECT 98.525 99.520 98.815 99.565 ;
        RECT 91.150 99.380 98.815 99.520 ;
        RECT 91.150 99.320 91.470 99.380 ;
        RECT 96.210 99.320 96.530 99.380 ;
        RECT 98.525 99.335 98.815 99.380 ;
        RECT 99.445 99.520 99.735 99.565 ;
        RECT 109.565 99.520 109.855 99.565 ;
        RECT 110.930 99.520 111.250 99.580 ;
        RECT 99.445 99.380 111.250 99.520 ;
        RECT 99.445 99.335 99.735 99.380 ;
        RECT 109.565 99.335 109.855 99.380 ;
        RECT 110.930 99.320 111.250 99.380 ;
        RECT 8.350 98.980 8.670 99.240 ;
        RECT 13.470 99.180 13.760 99.225 ;
        RECT 11.225 99.040 13.760 99.180 ;
        RECT 11.225 98.885 11.440 99.040 ;
        RECT 13.470 98.995 13.760 99.040 ;
        RECT 17.335 99.180 17.625 99.225 ;
        RECT 20.310 99.180 20.630 99.240 ;
        RECT 20.785 99.180 21.075 99.225 ;
        RECT 17.335 99.040 21.075 99.180 ;
        RECT 17.335 98.995 17.625 99.040 ;
        RECT 20.310 98.980 20.630 99.040 ;
        RECT 20.785 98.995 21.075 99.040 ;
        RECT 32.730 99.180 33.050 99.240 ;
        RECT 40.105 99.180 40.395 99.225 ;
        RECT 41.930 99.180 42.250 99.240 ;
        RECT 32.730 99.040 42.250 99.180 ;
        RECT 32.730 98.980 33.050 99.040 ;
        RECT 40.105 98.995 40.395 99.040 ;
        RECT 41.930 98.980 42.250 99.040 ;
        RECT 49.290 98.980 49.610 99.240 ;
        RECT 49.750 99.180 50.070 99.240 ;
        RECT 50.225 99.180 50.515 99.225 ;
        RECT 59.870 99.180 60.190 99.240 ;
        RECT 49.750 99.040 60.190 99.180 ;
        RECT 49.750 98.980 50.070 99.040 ;
        RECT 50.225 98.995 50.515 99.040 ;
        RECT 59.870 98.980 60.190 99.040 ;
        RECT 67.705 99.180 67.995 99.225 ;
        RECT 68.610 99.180 68.930 99.240 ;
        RECT 67.705 99.040 68.930 99.180 ;
        RECT 67.705 98.995 67.995 99.040 ;
        RECT 68.610 98.980 68.930 99.040 ;
        RECT 69.070 99.180 69.390 99.240 ;
        RECT 70.925 99.180 71.215 99.225 ;
        RECT 69.070 99.040 71.215 99.180 ;
        RECT 69.070 98.980 69.390 99.040 ;
        RECT 70.925 98.995 71.215 99.040 ;
        RECT 72.750 98.980 73.070 99.240 ;
        RECT 76.030 99.180 76.320 99.225 ;
        RECT 73.785 99.040 76.320 99.180 ;
        RECT 9.290 98.840 9.580 98.885 ;
        RECT 11.150 98.840 11.440 98.885 ;
        RECT 9.290 98.700 11.440 98.840 ;
        RECT 9.290 98.655 9.580 98.700 ;
        RECT 11.150 98.655 11.440 98.700 ;
        RECT 12.070 98.840 12.360 98.885 ;
        RECT 13.870 98.840 14.190 98.900 ;
        RECT 15.330 98.840 15.620 98.885 ;
        RECT 12.070 98.700 15.620 98.840 ;
        RECT 12.070 98.655 12.360 98.700 ;
        RECT 13.870 98.640 14.190 98.700 ;
        RECT 15.330 98.655 15.620 98.700 ;
        RECT 19.850 98.840 20.170 98.900 ;
        RECT 73.785 98.885 74.000 99.040 ;
        RECT 76.030 98.995 76.320 99.040 ;
        RECT 98.050 98.980 98.370 99.240 ;
        RECT 21.245 98.840 21.535 98.885 ;
        RECT 19.850 98.700 21.535 98.840 ;
        RECT 19.850 98.640 20.170 98.700 ;
        RECT 21.245 98.655 21.535 98.700 ;
        RECT 71.850 98.840 72.140 98.885 ;
        RECT 73.710 98.840 74.000 98.885 ;
        RECT 71.850 98.700 74.000 98.840 ;
        RECT 71.850 98.655 72.140 98.700 ;
        RECT 73.710 98.655 74.000 98.700 ;
        RECT 74.630 98.840 74.920 98.885 ;
        RECT 75.510 98.840 75.830 98.900 ;
        RECT 77.890 98.840 78.180 98.885 ;
        RECT 74.630 98.700 78.180 98.840 ;
        RECT 74.630 98.655 74.920 98.700 ;
        RECT 75.510 98.640 75.830 98.700 ;
        RECT 77.890 98.655 78.180 98.700 ;
        RECT 108.260 98.700 110.470 98.840 ;
        RECT 39.630 98.300 39.950 98.560 ;
        RECT 47.450 98.500 47.770 98.560 ;
        RECT 48.385 98.500 48.675 98.545 ;
        RECT 47.450 98.360 48.675 98.500 ;
        RECT 47.450 98.300 47.770 98.360 ;
        RECT 48.385 98.315 48.675 98.360 ;
        RECT 50.210 98.500 50.530 98.560 ;
        RECT 50.685 98.500 50.975 98.545 ;
        RECT 50.210 98.360 50.975 98.500 ;
        RECT 50.210 98.300 50.530 98.360 ;
        RECT 50.685 98.315 50.975 98.360 ;
        RECT 67.245 98.500 67.535 98.545 ;
        RECT 72.290 98.500 72.610 98.560 ;
        RECT 67.245 98.360 72.610 98.500 ;
        RECT 67.245 98.315 67.535 98.360 ;
        RECT 72.290 98.300 72.610 98.360 ;
        RECT 77.350 98.500 77.670 98.560 ;
        RECT 79.895 98.500 80.185 98.545 ;
        RECT 77.350 98.360 80.185 98.500 ;
        RECT 77.350 98.300 77.670 98.360 ;
        RECT 79.895 98.315 80.185 98.360 ;
        RECT 90.230 98.500 90.550 98.560 ;
        RECT 108.260 98.545 108.400 98.700 ;
        RECT 110.330 98.560 110.470 98.700 ;
        RECT 108.185 98.500 108.475 98.545 ;
        RECT 90.230 98.360 108.475 98.500 ;
        RECT 90.230 98.300 90.550 98.360 ;
        RECT 108.185 98.315 108.475 98.360 ;
        RECT 108.645 98.500 108.935 98.545 ;
        RECT 109.550 98.500 109.870 98.560 ;
        RECT 108.645 98.360 109.870 98.500 ;
        RECT 110.330 98.360 110.790 98.560 ;
        RECT 108.645 98.315 108.935 98.360 ;
        RECT 109.550 98.300 109.870 98.360 ;
        RECT 110.470 98.300 110.790 98.360 ;
        RECT 5.520 97.680 118.680 98.160 ;
        RECT 17.335 97.480 17.625 97.525 ;
        RECT 19.850 97.480 20.170 97.540 ;
        RECT 17.335 97.340 20.170 97.480 ;
        RECT 17.335 97.295 17.625 97.340 ;
        RECT 19.850 97.280 20.170 97.340 ;
        RECT 63.090 97.480 63.410 97.540 ;
        RECT 70.005 97.480 70.295 97.525 ;
        RECT 63.090 97.340 70.295 97.480 ;
        RECT 63.090 97.280 63.410 97.340 ;
        RECT 70.005 97.295 70.295 97.340 ;
        RECT 72.750 97.480 73.070 97.540 ;
        RECT 74.145 97.480 74.435 97.525 ;
        RECT 72.750 97.340 74.435 97.480 ;
        RECT 72.750 97.280 73.070 97.340 ;
        RECT 74.145 97.295 74.435 97.340 ;
        RECT 85.185 97.480 85.475 97.525 ;
        RECT 87.010 97.480 87.330 97.540 ;
        RECT 85.185 97.340 87.330 97.480 ;
        RECT 85.185 97.295 85.475 97.340 ;
        RECT 87.010 97.280 87.330 97.340 ;
        RECT 9.290 97.140 9.580 97.185 ;
        RECT 11.150 97.140 11.440 97.185 ;
        RECT 9.290 97.000 11.440 97.140 ;
        RECT 9.290 96.955 9.580 97.000 ;
        RECT 11.150 96.955 11.440 97.000 ;
        RECT 12.070 97.140 12.360 97.185 ;
        RECT 14.330 97.140 14.650 97.200 ;
        RECT 39.630 97.185 39.950 97.200 ;
        RECT 15.330 97.140 15.620 97.185 ;
        RECT 12.070 97.000 15.620 97.140 ;
        RECT 12.070 96.955 12.360 97.000 ;
        RECT 8.350 96.600 8.670 96.860 ;
        RECT 11.225 96.800 11.440 96.955 ;
        RECT 14.330 96.940 14.650 97.000 ;
        RECT 15.330 96.955 15.620 97.000 ;
        RECT 36.360 97.140 36.650 97.185 ;
        RECT 39.620 97.140 39.950 97.185 ;
        RECT 36.360 97.000 39.950 97.140 ;
        RECT 36.360 96.955 36.650 97.000 ;
        RECT 39.620 96.955 39.950 97.000 ;
        RECT 39.630 96.940 39.950 96.955 ;
        RECT 40.540 97.140 40.830 97.185 ;
        RECT 42.400 97.140 42.690 97.185 ;
        RECT 40.540 97.000 42.690 97.140 ;
        RECT 40.540 96.955 40.830 97.000 ;
        RECT 42.400 96.955 42.690 97.000 ;
        RECT 46.550 97.140 46.840 97.185 ;
        RECT 48.410 97.140 48.700 97.185 ;
        RECT 46.550 97.000 48.700 97.140 ;
        RECT 46.550 96.955 46.840 97.000 ;
        RECT 48.410 96.955 48.700 97.000 ;
        RECT 49.330 97.140 49.620 97.185 ;
        RECT 50.210 97.140 50.530 97.200 ;
        RECT 52.590 97.140 52.880 97.185 ;
        RECT 83.805 97.140 84.095 97.185 ;
        RECT 49.330 97.000 52.880 97.140 ;
        RECT 49.330 96.955 49.620 97.000 ;
        RECT 13.470 96.800 13.760 96.845 ;
        RECT 11.225 96.660 13.760 96.800 ;
        RECT 13.470 96.615 13.760 96.660 ;
        RECT 20.325 96.800 20.615 96.845 ;
        RECT 27.670 96.800 27.990 96.860 ;
        RECT 20.325 96.660 27.990 96.800 ;
        RECT 20.325 96.615 20.615 96.660 ;
        RECT 27.670 96.600 27.990 96.660 ;
        RECT 31.810 96.600 32.130 96.860 ;
        RECT 32.730 96.600 33.050 96.860 ;
        RECT 33.650 96.600 33.970 96.860 ;
        RECT 38.220 96.800 38.510 96.845 ;
        RECT 40.540 96.800 40.755 96.955 ;
        RECT 43.325 96.800 43.615 96.845 ;
        RECT 45.625 96.800 45.915 96.845 ;
        RECT 38.220 96.660 40.755 96.800 ;
        RECT 41.100 96.660 45.915 96.800 ;
        RECT 38.220 96.615 38.510 96.660 ;
        RECT 10.205 96.460 10.495 96.505 ;
        RECT 12.490 96.460 12.810 96.520 ;
        RECT 10.205 96.320 12.810 96.460 ;
        RECT 10.205 96.275 10.495 96.320 ;
        RECT 12.490 96.260 12.810 96.320 ;
        RECT 19.390 96.460 19.710 96.520 ;
        RECT 20.785 96.460 21.075 96.505 ;
        RECT 19.390 96.320 21.075 96.460 ;
        RECT 19.390 96.260 19.710 96.320 ;
        RECT 20.785 96.275 21.075 96.320 ;
        RECT 34.570 96.460 34.890 96.520 ;
        RECT 41.100 96.460 41.240 96.660 ;
        RECT 43.325 96.615 43.615 96.660 ;
        RECT 45.625 96.615 45.915 96.660 ;
        RECT 47.450 96.600 47.770 96.860 ;
        RECT 48.485 96.800 48.700 96.955 ;
        RECT 50.210 96.940 50.530 97.000 ;
        RECT 52.590 96.955 52.880 97.000 ;
        RECT 62.030 97.000 84.095 97.140 ;
        RECT 50.730 96.800 51.020 96.845 ;
        RECT 48.485 96.660 51.020 96.800 ;
        RECT 50.730 96.615 51.020 96.660 ;
        RECT 59.885 96.800 60.175 96.845 ;
        RECT 61.250 96.800 61.570 96.860 ;
        RECT 62.030 96.800 62.170 97.000 ;
        RECT 83.805 96.955 84.095 97.000 ;
        RECT 87.945 97.140 88.235 97.185 ;
        RECT 89.770 97.140 90.090 97.200 ;
        RECT 92.990 97.140 93.310 97.200 ;
        RECT 87.945 97.000 90.090 97.140 ;
        RECT 87.945 96.955 88.235 97.000 ;
        RECT 89.770 96.940 90.090 97.000 ;
        RECT 90.320 97.000 91.840 97.140 ;
        RECT 59.885 96.660 62.170 96.800 ;
        RECT 59.885 96.615 60.175 96.660 ;
        RECT 61.250 96.600 61.570 96.660 ;
        RECT 62.630 96.600 62.950 96.860 ;
        RECT 63.090 96.800 63.410 96.860 ;
        RECT 63.565 96.800 63.855 96.845 ;
        RECT 63.090 96.660 63.855 96.800 ;
        RECT 63.090 96.600 63.410 96.660 ;
        RECT 63.565 96.615 63.855 96.660 ;
        RECT 64.025 96.800 64.315 96.845 ;
        RECT 64.470 96.800 64.790 96.860 ;
        RECT 64.025 96.660 64.790 96.800 ;
        RECT 64.025 96.615 64.315 96.660 ;
        RECT 64.470 96.600 64.790 96.660 ;
        RECT 71.845 96.615 72.135 96.845 ;
        RECT 34.570 96.320 41.240 96.460 ;
        RECT 41.485 96.460 41.775 96.505 ;
        RECT 44.690 96.460 45.010 96.520 ;
        RECT 41.485 96.320 45.010 96.460 ;
        RECT 34.570 96.260 34.890 96.320 ;
        RECT 41.485 96.275 41.775 96.320 ;
        RECT 44.690 96.260 45.010 96.320 ;
        RECT 48.370 96.460 48.690 96.520 ;
        RECT 53.430 96.460 53.750 96.520 ;
        RECT 58.505 96.460 58.795 96.505 ;
        RECT 48.370 96.320 58.795 96.460 ;
        RECT 71.920 96.460 72.060 96.615 ;
        RECT 72.290 96.600 72.610 96.860 ;
        RECT 75.050 96.600 75.370 96.860 ;
        RECT 86.550 96.600 86.870 96.860 ;
        RECT 87.010 96.600 87.330 96.860 ;
        RECT 88.390 96.600 88.710 96.860 ;
        RECT 89.325 96.800 89.615 96.845 ;
        RECT 90.320 96.800 90.460 97.000 ;
        RECT 89.325 96.660 90.460 96.800 ;
        RECT 89.325 96.615 89.615 96.660 ;
        RECT 73.225 96.460 73.515 96.505 ;
        RECT 78.270 96.460 78.590 96.520 ;
        RECT 71.920 96.320 72.520 96.460 ;
        RECT 48.370 96.260 48.690 96.320 ;
        RECT 53.430 96.260 53.750 96.320 ;
        RECT 58.505 96.275 58.795 96.320 ;
        RECT 8.830 96.120 9.120 96.165 ;
        RECT 10.690 96.120 10.980 96.165 ;
        RECT 13.470 96.120 13.760 96.165 ;
        RECT 8.830 95.980 13.760 96.120 ;
        RECT 8.830 95.935 9.120 95.980 ;
        RECT 10.690 95.935 10.980 95.980 ;
        RECT 13.470 95.935 13.760 95.980 ;
        RECT 38.220 96.120 38.510 96.165 ;
        RECT 41.000 96.120 41.290 96.165 ;
        RECT 42.860 96.120 43.150 96.165 ;
        RECT 38.220 95.980 43.150 96.120 ;
        RECT 38.220 95.935 38.510 95.980 ;
        RECT 41.000 95.935 41.290 95.980 ;
        RECT 42.860 95.935 43.150 95.980 ;
        RECT 46.090 96.120 46.380 96.165 ;
        RECT 47.950 96.120 48.240 96.165 ;
        RECT 50.730 96.120 51.020 96.165 ;
        RECT 46.090 95.980 51.020 96.120 ;
        RECT 72.380 96.120 72.520 96.320 ;
        RECT 73.225 96.320 78.590 96.460 ;
        RECT 87.100 96.460 87.240 96.600 ;
        RECT 89.400 96.460 89.540 96.615 ;
        RECT 90.690 96.600 91.010 96.860 ;
        RECT 91.700 96.845 91.840 97.000 ;
        RECT 92.990 97.000 95.520 97.140 ;
        RECT 92.990 96.940 93.310 97.000 ;
        RECT 91.625 96.615 91.915 96.845 ;
        RECT 92.530 96.600 92.850 96.860 ;
        RECT 94.385 96.800 94.675 96.845 ;
        RECT 94.830 96.800 95.150 96.860 ;
        RECT 95.380 96.845 95.520 97.000 ;
        RECT 94.385 96.660 95.150 96.800 ;
        RECT 94.385 96.615 94.675 96.660 ;
        RECT 94.830 96.600 95.150 96.660 ;
        RECT 95.305 96.615 95.595 96.845 ;
        RECT 96.210 96.600 96.530 96.860 ;
        RECT 110.010 96.600 110.330 96.860 ;
        RECT 110.945 96.615 111.235 96.845 ;
        RECT 111.405 96.800 111.695 96.845 ;
        RECT 111.850 96.800 112.170 96.860 ;
        RECT 111.405 96.660 112.170 96.800 ;
        RECT 111.405 96.615 111.695 96.660 ;
        RECT 87.100 96.320 89.540 96.460 ;
        RECT 90.245 96.460 90.535 96.505 ;
        RECT 97.130 96.460 97.450 96.520 ;
        RECT 90.245 96.320 97.450 96.460 ;
        RECT 73.225 96.275 73.515 96.320 ;
        RECT 78.270 96.260 78.590 96.320 ;
        RECT 90.245 96.275 90.535 96.320 ;
        RECT 97.130 96.260 97.450 96.320 ;
        RECT 102.650 96.460 102.970 96.520 ;
        RECT 111.020 96.460 111.160 96.615 ;
        RECT 111.850 96.600 112.170 96.660 ;
        RECT 113.230 96.460 113.550 96.520 ;
        RECT 102.650 96.320 113.550 96.460 ;
        RECT 102.650 96.260 102.970 96.320 ;
        RECT 113.230 96.260 113.550 96.320 ;
        RECT 77.350 96.120 77.670 96.180 ;
        RECT 72.380 95.980 77.670 96.120 ;
        RECT 46.090 95.935 46.380 95.980 ;
        RECT 47.950 95.935 48.240 95.980 ;
        RECT 50.730 95.935 51.020 95.980 ;
        RECT 77.350 95.920 77.670 95.980 ;
        RECT 18.010 95.580 18.330 95.840 ;
        RECT 34.110 95.825 34.430 95.840 ;
        RECT 34.110 95.595 34.645 95.825 ;
        RECT 52.510 95.780 52.830 95.840 ;
        RECT 53.890 95.780 54.210 95.840 ;
        RECT 52.510 95.640 54.210 95.780 ;
        RECT 34.110 95.580 34.430 95.595 ;
        RECT 52.510 95.580 52.830 95.640 ;
        RECT 53.890 95.580 54.210 95.640 ;
        RECT 54.350 95.825 54.670 95.840 ;
        RECT 54.350 95.595 54.885 95.825 ;
        RECT 60.790 95.780 61.110 95.840 ;
        RECT 61.725 95.780 62.015 95.825 ;
        RECT 60.790 95.640 62.015 95.780 ;
        RECT 54.350 95.580 54.670 95.595 ;
        RECT 60.790 95.580 61.110 95.640 ;
        RECT 61.725 95.595 62.015 95.640 ;
        RECT 109.090 95.580 109.410 95.840 ;
        RECT 5.520 94.960 118.680 95.440 ;
        RECT 12.490 94.560 12.810 94.820 ;
        RECT 14.330 94.560 14.650 94.820 ;
        RECT 48.370 94.760 48.690 94.820 ;
        RECT 40.640 94.620 48.690 94.760 ;
        RECT 21.245 94.420 21.535 94.465 ;
        RECT 29.970 94.420 30.290 94.480 ;
        RECT 21.245 94.280 30.290 94.420 ;
        RECT 21.245 94.235 21.535 94.280 ;
        RECT 29.970 94.220 30.290 94.280 ;
        RECT 18.010 94.080 18.330 94.140 ;
        RECT 13.500 93.940 18.330 94.080 ;
        RECT 13.500 93.785 13.640 93.940 ;
        RECT 18.010 93.880 18.330 93.940 ;
        RECT 23.530 93.880 23.850 94.140 ;
        RECT 24.005 94.080 24.295 94.125 ;
        RECT 27.670 94.080 27.990 94.140 ;
        RECT 34.110 94.080 34.430 94.140 ;
        RECT 40.640 94.125 40.780 94.620 ;
        RECT 48.370 94.560 48.690 94.620 ;
        RECT 49.290 94.760 49.610 94.820 ;
        RECT 50.225 94.760 50.515 94.805 ;
        RECT 49.290 94.620 50.515 94.760 ;
        RECT 49.290 94.560 49.610 94.620 ;
        RECT 50.225 94.575 50.515 94.620 ;
        RECT 51.130 94.760 51.450 94.820 ;
        RECT 56.665 94.760 56.955 94.805 ;
        RECT 51.130 94.620 56.955 94.760 ;
        RECT 51.130 94.560 51.450 94.620 ;
        RECT 56.665 94.575 56.955 94.620 ;
        RECT 74.605 94.760 74.895 94.805 ;
        RECT 75.050 94.760 75.370 94.820 ;
        RECT 110.470 94.760 110.790 94.820 ;
        RECT 74.605 94.620 75.370 94.760 ;
        RECT 74.605 94.575 74.895 94.620 ;
        RECT 75.050 94.560 75.370 94.620 ;
        RECT 90.780 94.620 110.790 94.760 ;
        RECT 41.470 94.420 41.790 94.480 ;
        RECT 48.460 94.420 48.600 94.560 ;
        RECT 53.890 94.420 54.210 94.480 ;
        RECT 59.430 94.420 59.720 94.465 ;
        RECT 61.290 94.420 61.580 94.465 ;
        RECT 64.070 94.420 64.360 94.465 ;
        RECT 41.470 94.280 48.140 94.420 ;
        RECT 48.460 94.280 53.200 94.420 ;
        RECT 41.470 94.220 41.790 94.280 ;
        RECT 24.005 93.940 39.860 94.080 ;
        RECT 24.005 93.895 24.295 93.940 ;
        RECT 27.670 93.880 27.990 93.940 ;
        RECT 34.110 93.880 34.430 93.940 ;
        RECT 13.425 93.555 13.715 93.785 ;
        RECT 14.790 93.540 15.110 93.800 ;
        RECT 19.850 93.540 20.170 93.800 ;
        RECT 20.325 93.740 20.615 93.785 ;
        RECT 22.150 93.740 22.470 93.800 ;
        RECT 22.625 93.740 22.915 93.785 ;
        RECT 24.925 93.740 25.215 93.785 ;
        RECT 20.325 93.600 25.215 93.740 ;
        RECT 20.325 93.555 20.615 93.600 ;
        RECT 22.150 93.540 22.470 93.600 ;
        RECT 22.625 93.555 22.915 93.600 ;
        RECT 24.925 93.555 25.215 93.600 ;
        RECT 25.000 93.400 25.140 93.555 ;
        RECT 26.750 93.540 27.070 93.800 ;
        RECT 27.225 93.740 27.515 93.785 ;
        RECT 32.730 93.740 33.050 93.800 ;
        RECT 27.225 93.600 33.050 93.740 ;
        RECT 27.225 93.555 27.515 93.600 ;
        RECT 27.300 93.400 27.440 93.555 ;
        RECT 32.730 93.540 33.050 93.600 ;
        RECT 38.725 93.740 39.015 93.785 ;
        RECT 39.170 93.740 39.490 93.800 ;
        RECT 38.725 93.600 39.490 93.740 ;
        RECT 39.720 93.740 39.860 93.940 ;
        RECT 40.565 93.895 40.855 94.125 ;
        RECT 41.025 94.080 41.315 94.125 ;
        RECT 41.025 93.940 47.680 94.080 ;
        RECT 41.025 93.895 41.315 93.940 ;
        RECT 41.485 93.740 41.775 93.785 ;
        RECT 45.625 93.740 45.915 93.785 ;
        RECT 39.720 93.600 41.775 93.740 ;
        RECT 38.725 93.555 39.015 93.600 ;
        RECT 39.170 93.540 39.490 93.600 ;
        RECT 41.485 93.555 41.775 93.600 ;
        RECT 43.400 93.600 45.915 93.740 ;
        RECT 25.000 93.260 27.440 93.400 ;
        RECT 37.330 93.200 37.650 93.460 ;
        RECT 21.690 92.860 22.010 93.120 ;
        RECT 25.845 93.060 26.135 93.105 ;
        RECT 26.750 93.060 27.070 93.120 ;
        RECT 25.845 92.920 27.070 93.060 ;
        RECT 25.845 92.875 26.135 92.920 ;
        RECT 26.750 92.860 27.070 92.920 ;
        RECT 28.130 92.860 28.450 93.120 ;
        RECT 30.905 93.060 31.195 93.105 ;
        RECT 34.570 93.060 34.890 93.120 ;
        RECT 30.905 92.920 34.890 93.060 ;
        RECT 30.905 92.875 31.195 92.920 ;
        RECT 34.570 92.860 34.890 92.920 ;
        RECT 37.790 92.860 38.110 93.120 ;
        RECT 43.400 93.105 43.540 93.600 ;
        RECT 45.625 93.555 45.915 93.600 ;
        RECT 47.540 93.400 47.680 93.940 ;
        RECT 48.000 93.785 48.140 94.280 ;
        RECT 48.460 93.940 52.280 94.080 ;
        RECT 47.925 93.555 48.215 93.785 ;
        RECT 48.460 93.400 48.600 93.940 ;
        RECT 52.140 93.785 52.280 93.940 ;
        RECT 52.510 93.880 52.830 94.140 ;
        RECT 53.060 94.125 53.200 94.280 ;
        RECT 53.890 94.280 58.720 94.420 ;
        RECT 53.890 94.220 54.210 94.280 ;
        RECT 52.985 93.895 53.275 94.125 ;
        RECT 54.350 94.080 54.670 94.140 ;
        RECT 58.580 94.125 58.720 94.280 ;
        RECT 59.430 94.280 64.360 94.420 ;
        RECT 59.430 94.235 59.720 94.280 ;
        RECT 61.290 94.235 61.580 94.280 ;
        RECT 64.070 94.235 64.360 94.280 ;
        RECT 56.205 94.080 56.495 94.125 ;
        RECT 53.980 93.940 56.495 94.080 ;
        RECT 48.845 93.555 49.135 93.785 ;
        RECT 52.065 93.740 52.355 93.785 ;
        RECT 53.980 93.740 54.120 93.940 ;
        RECT 54.350 93.880 54.670 93.940 ;
        RECT 56.205 93.895 56.495 93.940 ;
        RECT 58.505 93.895 58.795 94.125 ;
        RECT 58.965 94.080 59.255 94.125 ;
        RECT 69.070 94.080 69.390 94.140 ;
        RECT 58.965 93.940 69.390 94.080 ;
        RECT 58.965 93.895 59.255 93.940 ;
        RECT 69.070 93.880 69.390 93.940 ;
        RECT 77.825 94.080 78.115 94.125 ;
        RECT 78.270 94.080 78.590 94.140 ;
        RECT 77.825 93.940 78.590 94.080 ;
        RECT 77.825 93.895 78.115 93.940 ;
        RECT 78.270 93.880 78.590 93.940 ;
        RECT 85.645 94.080 85.935 94.125 ;
        RECT 90.230 94.080 90.550 94.140 ;
        RECT 90.780 94.125 90.920 94.620 ;
        RECT 110.470 94.560 110.790 94.620 ;
        RECT 106.810 94.420 107.100 94.465 ;
        RECT 108.670 94.420 108.960 94.465 ;
        RECT 111.450 94.420 111.740 94.465 ;
        RECT 106.810 94.280 111.740 94.420 ;
        RECT 106.810 94.235 107.100 94.280 ;
        RECT 108.670 94.235 108.960 94.280 ;
        RECT 111.450 94.235 111.740 94.280 ;
        RECT 85.645 93.940 90.550 94.080 ;
        RECT 85.645 93.895 85.935 93.940 ;
        RECT 90.230 93.880 90.550 93.940 ;
        RECT 90.705 93.895 90.995 94.125 ;
        RECT 108.185 94.080 108.475 94.125 ;
        RECT 109.090 94.080 109.410 94.140 ;
        RECT 108.185 93.940 109.410 94.080 ;
        RECT 108.185 93.895 108.475 93.940 ;
        RECT 109.090 93.880 109.410 93.940 ;
        RECT 52.065 93.600 54.120 93.740 ;
        RECT 55.285 93.740 55.575 93.785 ;
        RECT 57.585 93.740 57.875 93.785 ;
        RECT 58.030 93.740 58.350 93.800 ;
        RECT 55.285 93.600 58.350 93.740 ;
        RECT 52.065 93.555 52.355 93.600 ;
        RECT 55.285 93.555 55.575 93.600 ;
        RECT 57.585 93.555 57.875 93.600 ;
        RECT 47.540 93.260 48.600 93.400 ;
        RECT 48.920 93.400 49.060 93.555 ;
        RECT 52.510 93.400 52.830 93.460 ;
        RECT 54.365 93.400 54.655 93.445 ;
        RECT 48.920 93.260 51.820 93.400 ;
        RECT 43.325 92.875 43.615 93.105 ;
        RECT 44.690 92.860 45.010 93.120 ;
        RECT 49.750 92.860 50.070 93.120 ;
        RECT 51.680 93.060 51.820 93.260 ;
        RECT 52.510 93.260 54.655 93.400 ;
        RECT 52.510 93.200 52.830 93.260 ;
        RECT 54.365 93.215 54.655 93.260 ;
        RECT 55.360 93.060 55.500 93.555 ;
        RECT 58.030 93.540 58.350 93.600 ;
        RECT 60.790 93.540 61.110 93.800 ;
        RECT 64.070 93.740 64.360 93.785 ;
        RECT 61.825 93.600 64.360 93.740 ;
        RECT 61.825 93.445 62.040 93.600 ;
        RECT 64.070 93.555 64.360 93.600 ;
        RECT 64.930 93.740 65.250 93.800 ;
        RECT 84.725 93.740 85.015 93.785 ;
        RECT 87.010 93.740 87.330 93.800 ;
        RECT 89.785 93.740 90.075 93.785 ;
        RECT 92.085 93.740 92.375 93.785 ;
        RECT 64.930 93.600 92.375 93.740 ;
        RECT 64.930 93.540 65.250 93.600 ;
        RECT 84.725 93.555 85.015 93.600 ;
        RECT 87.010 93.540 87.330 93.600 ;
        RECT 89.785 93.555 90.075 93.600 ;
        RECT 92.085 93.555 92.375 93.600 ;
        RECT 93.005 93.555 93.295 93.785 ;
        RECT 59.890 93.400 60.180 93.445 ;
        RECT 61.750 93.400 62.040 93.445 ;
        RECT 59.890 93.260 62.040 93.400 ;
        RECT 59.890 93.215 60.180 93.260 ;
        RECT 61.750 93.215 62.040 93.260 ;
        RECT 62.670 93.400 62.960 93.445 ;
        RECT 64.470 93.400 64.790 93.460 ;
        RECT 65.930 93.400 66.220 93.445 ;
        RECT 62.670 93.260 66.220 93.400 ;
        RECT 62.670 93.215 62.960 93.260 ;
        RECT 64.470 93.200 64.790 93.260 ;
        RECT 65.930 93.215 66.220 93.260 ;
        RECT 69.070 93.400 69.390 93.460 ;
        RECT 86.105 93.400 86.395 93.445 ;
        RECT 90.230 93.400 90.550 93.460 ;
        RECT 69.070 93.260 90.550 93.400 ;
        RECT 93.080 93.400 93.220 93.555 ;
        RECT 93.450 93.540 93.770 93.800 ;
        RECT 99.445 93.740 99.735 93.785 ;
        RECT 102.650 93.740 102.970 93.800 ;
        RECT 99.445 93.600 102.970 93.740 ;
        RECT 99.445 93.555 99.735 93.600 ;
        RECT 102.650 93.540 102.970 93.600 ;
        RECT 103.110 93.740 103.430 93.800 ;
        RECT 106.345 93.740 106.635 93.785 ;
        RECT 111.450 93.740 111.740 93.785 ;
        RECT 103.110 93.600 106.635 93.740 ;
        RECT 103.110 93.540 103.430 93.600 ;
        RECT 106.345 93.555 106.635 93.600 ;
        RECT 109.205 93.600 111.740 93.740 ;
        RECT 109.205 93.445 109.420 93.600 ;
        RECT 111.450 93.555 111.740 93.600 ;
        RECT 107.270 93.400 107.560 93.445 ;
        RECT 109.130 93.400 109.420 93.445 ;
        RECT 93.080 93.260 105.640 93.400 ;
        RECT 69.070 93.200 69.390 93.260 ;
        RECT 86.105 93.215 86.395 93.260 ;
        RECT 90.230 93.200 90.550 93.260 ;
        RECT 51.680 92.920 55.500 93.060 ;
        RECT 66.770 93.060 67.090 93.120 ;
        RECT 67.935 93.060 68.225 93.105 ;
        RECT 66.770 92.920 68.225 93.060 ;
        RECT 66.770 92.860 67.090 92.920 ;
        RECT 67.935 92.875 68.225 92.920 ;
        RECT 76.430 92.860 76.750 93.120 ;
        RECT 76.905 93.060 77.195 93.105 ;
        RECT 77.350 93.060 77.670 93.120 ;
        RECT 76.905 92.920 77.670 93.060 ;
        RECT 76.905 92.875 77.195 92.920 ;
        RECT 77.350 92.860 77.670 92.920 ;
        RECT 83.330 93.060 83.650 93.120 ;
        RECT 83.805 93.060 84.095 93.105 ;
        RECT 83.330 92.920 84.095 93.060 ;
        RECT 83.330 92.860 83.650 92.920 ;
        RECT 83.805 92.875 84.095 92.920 ;
        RECT 87.930 93.060 88.250 93.120 ;
        RECT 88.865 93.060 89.155 93.105 ;
        RECT 87.930 92.920 89.155 93.060 ;
        RECT 87.930 92.860 88.250 92.920 ;
        RECT 88.865 92.875 89.155 92.920 ;
        RECT 89.310 93.060 89.630 93.120 ;
        RECT 91.165 93.060 91.455 93.105 ;
        RECT 89.310 92.920 91.455 93.060 ;
        RECT 89.310 92.860 89.630 92.920 ;
        RECT 91.165 92.875 91.455 92.920 ;
        RECT 94.385 93.060 94.675 93.105 ;
        RECT 95.290 93.060 95.610 93.120 ;
        RECT 94.385 92.920 95.610 93.060 ;
        RECT 94.385 92.875 94.675 92.920 ;
        RECT 95.290 92.860 95.610 92.920 ;
        RECT 98.970 92.860 99.290 93.120 ;
        RECT 105.500 93.060 105.640 93.260 ;
        RECT 107.270 93.260 109.420 93.400 ;
        RECT 107.270 93.215 107.560 93.260 ;
        RECT 109.130 93.215 109.420 93.260 ;
        RECT 110.050 93.400 110.340 93.445 ;
        RECT 111.850 93.400 112.170 93.460 ;
        RECT 113.310 93.400 113.600 93.445 ;
        RECT 110.050 93.260 113.600 93.400 ;
        RECT 110.050 93.215 110.340 93.260 ;
        RECT 111.850 93.200 112.170 93.260 ;
        RECT 113.310 93.215 113.600 93.260 ;
        RECT 109.550 93.060 109.870 93.120 ;
        RECT 115.315 93.060 115.605 93.105 ;
        RECT 105.500 92.920 115.605 93.060 ;
        RECT 109.550 92.860 109.870 92.920 ;
        RECT 115.315 92.875 115.605 92.920 ;
        RECT 5.520 92.240 118.680 92.720 ;
        RECT 58.030 91.840 58.350 92.100 ;
        RECT 61.250 91.840 61.570 92.100 ;
        RECT 62.630 92.040 62.950 92.100 ;
        RECT 63.565 92.040 63.855 92.085 ;
        RECT 62.630 91.900 63.855 92.040 ;
        RECT 62.630 91.840 62.950 91.900 ;
        RECT 63.565 91.855 63.855 91.900 ;
        RECT 65.865 92.040 66.155 92.085 ;
        RECT 66.770 92.040 67.090 92.100 ;
        RECT 65.865 91.900 67.090 92.040 ;
        RECT 65.865 91.855 66.155 91.900 ;
        RECT 66.770 91.840 67.090 91.900 ;
        RECT 90.230 92.040 90.550 92.100 ;
        RECT 90.705 92.040 90.995 92.085 ;
        RECT 90.230 91.900 90.995 92.040 ;
        RECT 90.230 91.840 90.550 91.900 ;
        RECT 90.705 91.855 90.995 91.900 ;
        RECT 109.105 92.040 109.395 92.085 ;
        RECT 110.010 92.040 110.330 92.100 ;
        RECT 109.105 91.900 110.330 92.040 ;
        RECT 109.105 91.855 109.395 91.900 ;
        RECT 58.120 91.700 58.260 91.840 ;
        RECT 64.930 91.700 65.250 91.760 ;
        RECT 58.120 91.560 65.250 91.700 ;
        RECT 20.770 91.360 21.090 91.420 ;
        RECT 21.245 91.360 21.535 91.405 ;
        RECT 20.770 91.220 21.535 91.360 ;
        RECT 20.770 91.160 21.090 91.220 ;
        RECT 21.245 91.175 21.535 91.220 ;
        RECT 22.150 91.160 22.470 91.420 ;
        RECT 32.745 91.360 33.035 91.405 ;
        RECT 34.570 91.360 34.890 91.420 ;
        RECT 32.745 91.220 34.890 91.360 ;
        RECT 32.745 91.175 33.035 91.220 ;
        RECT 34.570 91.160 34.890 91.220 ;
        RECT 41.930 91.360 42.250 91.420 ;
        RECT 43.785 91.360 44.075 91.405 ;
        RECT 44.690 91.360 45.010 91.420 ;
        RECT 41.930 91.220 45.010 91.360 ;
        RECT 41.930 91.160 42.250 91.220 ;
        RECT 43.785 91.175 44.075 91.220 ;
        RECT 44.690 91.160 45.010 91.220 ;
        RECT 52.970 91.160 53.290 91.420 ;
        RECT 53.445 91.360 53.735 91.405 ;
        RECT 58.120 91.360 58.260 91.560 ;
        RECT 64.930 91.500 65.250 91.560 ;
        RECT 65.405 91.700 65.695 91.745 ;
        RECT 67.230 91.700 67.550 91.760 ;
        RECT 68.610 91.700 68.930 91.760 ;
        RECT 65.405 91.560 68.930 91.700 ;
        RECT 65.405 91.515 65.695 91.560 ;
        RECT 67.230 91.500 67.550 91.560 ;
        RECT 68.610 91.500 68.930 91.560 ;
        RECT 83.790 91.700 84.110 91.760 ;
        RECT 84.265 91.700 84.555 91.745 ;
        RECT 83.790 91.560 84.555 91.700 ;
        RECT 83.790 91.500 84.110 91.560 ;
        RECT 84.265 91.515 84.555 91.560 ;
        RECT 53.445 91.220 58.260 91.360 ;
        RECT 58.505 91.360 58.795 91.405 ;
        RECT 60.330 91.360 60.650 91.420 ;
        RECT 62.185 91.360 62.475 91.405 ;
        RECT 58.505 91.220 62.475 91.360 ;
        RECT 90.780 91.360 90.920 91.855 ;
        RECT 110.010 91.840 110.330 91.900 ;
        RECT 110.470 92.040 110.790 92.100 ;
        RECT 111.405 92.040 111.695 92.085 ;
        RECT 110.470 91.900 111.695 92.040 ;
        RECT 110.470 91.840 110.790 91.900 ;
        RECT 111.405 91.855 111.695 91.900 ;
        RECT 94.390 91.700 94.680 91.745 ;
        RECT 96.250 91.700 96.540 91.745 ;
        RECT 94.390 91.560 96.540 91.700 ;
        RECT 94.390 91.515 94.680 91.560 ;
        RECT 96.250 91.515 96.540 91.560 ;
        RECT 97.170 91.700 97.460 91.745 ;
        RECT 98.970 91.700 99.290 91.760 ;
        RECT 100.430 91.700 100.720 91.745 ;
        RECT 97.170 91.560 100.720 91.700 ;
        RECT 97.170 91.515 97.460 91.560 ;
        RECT 93.465 91.360 93.755 91.405 ;
        RECT 96.325 91.360 96.540 91.515 ;
        RECT 98.970 91.500 99.290 91.560 ;
        RECT 100.430 91.515 100.720 91.560 ;
        RECT 109.550 91.700 109.870 91.760 ;
        RECT 110.945 91.700 111.235 91.745 ;
        RECT 109.550 91.560 111.235 91.700 ;
        RECT 109.550 91.500 109.870 91.560 ;
        RECT 110.945 91.515 111.235 91.560 ;
        RECT 98.570 91.360 98.860 91.405 ;
        RECT 90.780 91.220 95.980 91.360 ;
        RECT 96.325 91.220 98.860 91.360 ;
        RECT 53.445 91.175 53.735 91.220 ;
        RECT 58.505 91.175 58.795 91.220 ;
        RECT 60.330 91.160 60.650 91.220 ;
        RECT 62.185 91.175 62.475 91.220 ;
        RECT 93.465 91.175 93.755 91.220 ;
        RECT 58.950 91.020 59.270 91.080 ;
        RECT 59.425 91.020 59.715 91.065 ;
        RECT 58.950 90.880 59.715 91.020 ;
        RECT 58.950 90.820 59.270 90.880 ;
        RECT 59.425 90.835 59.715 90.880 ;
        RECT 63.550 91.020 63.870 91.080 ;
        RECT 66.325 91.020 66.615 91.065 ;
        RECT 68.150 91.020 68.470 91.080 ;
        RECT 63.550 90.880 68.470 91.020 ;
        RECT 63.550 90.820 63.870 90.880 ;
        RECT 66.325 90.835 66.615 90.880 ;
        RECT 68.150 90.820 68.470 90.880 ;
        RECT 95.290 90.820 95.610 91.080 ;
        RECT 95.840 91.020 95.980 91.220 ;
        RECT 98.570 91.175 98.860 91.220 ;
        RECT 103.125 91.360 103.415 91.405 ;
        RECT 104.490 91.360 104.810 91.420 ;
        RECT 103.125 91.220 104.810 91.360 ;
        RECT 103.125 91.175 103.415 91.220 ;
        RECT 104.490 91.160 104.810 91.220 ;
        RECT 96.670 91.020 96.990 91.080 ;
        RECT 95.840 90.880 96.990 91.020 ;
        RECT 96.670 90.820 96.990 90.880 ;
        RECT 110.930 91.020 111.250 91.080 ;
        RECT 111.865 91.020 112.155 91.065 ;
        RECT 110.930 90.880 112.155 91.020 ;
        RECT 110.930 90.820 111.250 90.880 ;
        RECT 111.865 90.835 112.155 90.880 ;
        RECT 14.790 90.680 15.110 90.740 ;
        RECT 30.430 90.680 30.750 90.740 ;
        RECT 14.790 90.540 30.750 90.680 ;
        RECT 14.790 90.480 15.110 90.540 ;
        RECT 30.430 90.480 30.750 90.540 ;
        RECT 32.730 90.680 33.050 90.740 ;
        RECT 63.105 90.680 63.395 90.725 ;
        RECT 92.990 90.680 93.310 90.740 ;
        RECT 32.730 90.540 93.310 90.680 ;
        RECT 32.730 90.480 33.050 90.540 ;
        RECT 63.105 90.495 63.395 90.540 ;
        RECT 92.990 90.480 93.310 90.540 ;
        RECT 93.930 90.680 94.220 90.725 ;
        RECT 95.790 90.680 96.080 90.725 ;
        RECT 98.570 90.680 98.860 90.725 ;
        RECT 93.930 90.540 98.860 90.680 ;
        RECT 93.930 90.495 94.220 90.540 ;
        RECT 95.790 90.495 96.080 90.540 ;
        RECT 98.570 90.495 98.860 90.540 ;
        RECT 23.070 90.140 23.390 90.400 ;
        RECT 42.390 90.340 42.710 90.400 ;
        RECT 43.325 90.340 43.615 90.385 ;
        RECT 42.390 90.200 43.615 90.340 ;
        RECT 42.390 90.140 42.710 90.200 ;
        RECT 43.325 90.155 43.615 90.200 ;
        RECT 52.970 90.340 53.290 90.400 ;
        RECT 54.365 90.340 54.655 90.385 ;
        RECT 52.970 90.200 54.655 90.340 ;
        RECT 93.080 90.340 93.220 90.480 ;
        RECT 98.970 90.340 99.290 90.400 ;
        RECT 93.080 90.200 99.290 90.340 ;
        RECT 52.970 90.140 53.290 90.200 ;
        RECT 54.365 90.155 54.655 90.200 ;
        RECT 98.970 90.140 99.290 90.200 ;
        RECT 102.190 90.385 102.510 90.400 ;
        RECT 102.190 90.155 102.725 90.385 ;
        RECT 102.190 90.140 102.510 90.155 ;
        RECT 104.030 90.140 104.350 90.400 ;
        RECT 5.520 89.520 118.680 90.000 ;
        RECT 21.690 89.120 22.010 89.380 ;
        RECT 22.610 89.320 22.930 89.380 ;
        RECT 23.085 89.320 23.375 89.365 ;
        RECT 22.610 89.180 23.375 89.320 ;
        RECT 22.610 89.120 22.930 89.180 ;
        RECT 23.085 89.135 23.375 89.180 ;
        RECT 28.130 89.120 28.450 89.380 ;
        RECT 29.510 89.120 29.830 89.380 ;
        RECT 31.810 89.120 32.130 89.380 ;
        RECT 33.190 89.320 33.510 89.380 ;
        RECT 34.125 89.320 34.415 89.365 ;
        RECT 33.190 89.180 34.415 89.320 ;
        RECT 33.190 89.120 33.510 89.180 ;
        RECT 34.125 89.135 34.415 89.180 ;
        RECT 38.250 89.320 38.570 89.380 ;
        RECT 49.750 89.320 50.070 89.380 ;
        RECT 52.525 89.320 52.815 89.365 ;
        RECT 38.250 89.180 45.380 89.320 ;
        RECT 38.250 89.120 38.570 89.180 ;
        RECT 35.050 88.980 35.340 89.025 ;
        RECT 36.910 88.980 37.200 89.025 ;
        RECT 39.690 88.980 39.980 89.025 ;
        RECT 23.620 88.840 32.960 88.980 ;
        RECT 23.620 88.360 23.760 88.840 ;
        RECT 28.145 88.640 28.435 88.685 ;
        RECT 30.890 88.640 31.210 88.700 ;
        RECT 28.145 88.500 31.210 88.640 ;
        RECT 28.145 88.455 28.435 88.500 ;
        RECT 30.890 88.440 31.210 88.500 ;
        RECT 32.270 88.440 32.590 88.700 ;
        RECT 32.820 88.640 32.960 88.840 ;
        RECT 35.050 88.840 39.980 88.980 ;
        RECT 45.240 88.980 45.380 89.180 ;
        RECT 49.750 89.180 52.815 89.320 ;
        RECT 49.750 89.120 50.070 89.180 ;
        RECT 52.525 89.135 52.815 89.180 ;
        RECT 82.410 89.320 82.730 89.380 ;
        RECT 88.405 89.320 88.695 89.365 ;
        RECT 88.850 89.320 89.170 89.380 ;
        RECT 82.410 89.180 86.320 89.320 ;
        RECT 82.410 89.120 82.730 89.180 ;
        RECT 51.605 88.980 51.895 89.025 ;
        RECT 45.240 88.840 51.895 88.980 ;
        RECT 35.050 88.795 35.340 88.840 ;
        RECT 36.910 88.795 37.200 88.840 ;
        RECT 39.690 88.795 39.980 88.840 ;
        RECT 51.605 88.795 51.895 88.840 ;
        RECT 71.850 88.980 72.140 89.025 ;
        RECT 73.710 88.980 74.000 89.025 ;
        RECT 76.490 88.980 76.780 89.025 ;
        RECT 71.850 88.840 76.780 88.980 ;
        RECT 71.850 88.795 72.140 88.840 ;
        RECT 73.710 88.795 74.000 88.840 ;
        RECT 76.490 88.795 76.780 88.840 ;
        RECT 77.350 88.980 77.670 89.040 ;
        RECT 77.350 88.840 85.860 88.980 ;
        RECT 77.350 88.780 77.670 88.840 ;
        RECT 36.425 88.640 36.715 88.685 ;
        RECT 37.790 88.640 38.110 88.700 ;
        RECT 32.820 88.500 35.260 88.640 ;
        RECT 35.120 88.360 35.260 88.500 ;
        RECT 36.425 88.500 38.110 88.640 ;
        RECT 36.425 88.455 36.715 88.500 ;
        RECT 37.790 88.440 38.110 88.500 ;
        RECT 41.470 88.640 41.790 88.700 ;
        RECT 43.555 88.640 43.845 88.685 ;
        RECT 46.530 88.640 46.850 88.700 ;
        RECT 41.470 88.500 46.850 88.640 ;
        RECT 41.470 88.440 41.790 88.500 ;
        RECT 43.555 88.455 43.845 88.500 ;
        RECT 46.530 88.440 46.850 88.500 ;
        RECT 49.290 88.640 49.610 88.700 ;
        RECT 52.985 88.640 53.275 88.685 ;
        RECT 49.290 88.500 53.275 88.640 ;
        RECT 49.290 88.440 49.610 88.500 ;
        RECT 52.985 88.455 53.275 88.500 ;
        RECT 69.545 88.640 69.835 88.685 ;
        RECT 83.790 88.640 84.110 88.700 ;
        RECT 69.545 88.500 84.110 88.640 ;
        RECT 69.545 88.455 69.835 88.500 ;
        RECT 83.790 88.440 84.110 88.500 ;
        RECT 13.885 88.300 14.175 88.345 ;
        RECT 19.850 88.300 20.170 88.360 ;
        RECT 13.885 88.160 20.170 88.300 ;
        RECT 13.885 88.115 14.175 88.160 ;
        RECT 19.850 88.100 20.170 88.160 ;
        RECT 21.690 88.100 22.010 88.360 ;
        RECT 22.150 88.100 22.470 88.360 ;
        RECT 23.530 88.100 23.850 88.360 ;
        RECT 23.990 88.300 24.310 88.360 ;
        RECT 24.465 88.300 24.755 88.345 ;
        RECT 23.990 88.160 24.755 88.300 ;
        RECT 23.990 88.100 24.310 88.160 ;
        RECT 24.465 88.115 24.755 88.160 ;
        RECT 24.910 88.100 25.230 88.360 ;
        RECT 25.385 88.300 25.675 88.345 ;
        RECT 28.605 88.300 28.895 88.345 ;
        RECT 29.050 88.300 29.370 88.360 ;
        RECT 25.385 88.160 28.460 88.300 ;
        RECT 25.385 88.115 25.675 88.160 ;
        RECT 20.770 87.760 21.090 88.020 ;
        RECT 22.610 87.960 22.930 88.020 ;
        RECT 25.460 87.960 25.600 88.115 ;
        RECT 22.610 87.820 25.600 87.960 ;
        RECT 26.765 87.960 27.055 88.005 ;
        RECT 27.225 87.960 27.515 88.005 ;
        RECT 26.765 87.820 27.515 87.960 ;
        RECT 28.320 87.960 28.460 88.160 ;
        RECT 28.605 88.160 29.370 88.300 ;
        RECT 28.605 88.115 28.895 88.160 ;
        RECT 29.050 88.100 29.370 88.160 ;
        RECT 30.430 88.100 30.750 88.360 ;
        RECT 33.190 88.100 33.510 88.360 ;
        RECT 34.570 88.100 34.890 88.360 ;
        RECT 35.030 88.100 35.350 88.360 ;
        RECT 39.690 88.300 39.980 88.345 ;
        RECT 37.445 88.160 39.980 88.300 ;
        RECT 28.320 87.820 31.580 87.960 ;
        RECT 22.610 87.760 22.930 87.820 ;
        RECT 26.765 87.775 27.055 87.820 ;
        RECT 27.225 87.775 27.515 87.820 ;
        RECT 12.030 87.620 12.350 87.680 ;
        RECT 12.965 87.620 13.255 87.665 ;
        RECT 12.030 87.480 13.255 87.620 ;
        RECT 12.030 87.420 12.350 87.480 ;
        RECT 12.965 87.435 13.255 87.480 ;
        RECT 30.430 87.620 30.750 87.680 ;
        RECT 30.905 87.620 31.195 87.665 ;
        RECT 30.430 87.480 31.195 87.620 ;
        RECT 31.440 87.620 31.580 87.820 ;
        RECT 31.810 87.760 32.130 88.020 ;
        RECT 37.445 88.005 37.660 88.160 ;
        RECT 39.690 88.115 39.980 88.160 ;
        RECT 44.690 88.100 45.010 88.360 ;
        RECT 52.510 88.100 52.830 88.360 ;
        RECT 66.325 88.300 66.615 88.345 ;
        RECT 53.060 88.160 66.615 88.300 ;
        RECT 35.510 87.960 35.800 88.005 ;
        RECT 37.370 87.960 37.660 88.005 ;
        RECT 35.510 87.820 37.660 87.960 ;
        RECT 35.510 87.775 35.800 87.820 ;
        RECT 37.370 87.775 37.660 87.820 ;
        RECT 38.290 87.960 38.580 88.005 ;
        RECT 41.550 87.960 41.840 88.005 ;
        RECT 42.390 87.960 42.710 88.020 ;
        RECT 47.910 87.960 48.230 88.020 ;
        RECT 53.060 87.960 53.200 88.160 ;
        RECT 66.325 88.115 66.615 88.160 ;
        RECT 38.290 87.820 42.710 87.960 ;
        RECT 38.290 87.775 38.580 87.820 ;
        RECT 41.550 87.775 41.840 87.820 ;
        RECT 42.390 87.760 42.710 87.820 ;
        RECT 42.940 87.820 45.840 87.960 ;
        RECT 32.730 87.620 33.050 87.680 ;
        RECT 42.940 87.620 43.080 87.820 ;
        RECT 31.440 87.480 43.080 87.620 ;
        RECT 44.690 87.620 45.010 87.680 ;
        RECT 45.165 87.620 45.455 87.665 ;
        RECT 44.690 87.480 45.455 87.620 ;
        RECT 45.700 87.620 45.840 87.820 ;
        RECT 47.910 87.820 53.200 87.960 ;
        RECT 47.910 87.760 48.230 87.820 ;
        RECT 53.890 87.760 54.210 88.020 ;
        RECT 66.400 87.960 66.540 88.115 ;
        RECT 67.230 88.100 67.550 88.360 ;
        RECT 67.690 88.100 68.010 88.360 ;
        RECT 68.150 88.100 68.470 88.360 ;
        RECT 69.070 88.300 69.390 88.360 ;
        RECT 71.385 88.300 71.675 88.345 ;
        RECT 69.070 88.160 71.675 88.300 ;
        RECT 69.070 88.100 69.390 88.160 ;
        RECT 71.385 88.115 71.675 88.160 ;
        RECT 73.210 88.100 73.530 88.360 ;
        RECT 76.490 88.300 76.780 88.345 ;
        RECT 74.245 88.160 76.780 88.300 ;
        RECT 68.610 87.960 68.930 88.020 ;
        RECT 74.245 88.005 74.460 88.160 ;
        RECT 76.490 88.115 76.780 88.160 ;
        RECT 80.570 88.300 80.890 88.360 ;
        RECT 81.045 88.300 81.335 88.345 ;
        RECT 80.570 88.160 81.335 88.300 ;
        RECT 80.570 88.100 80.890 88.160 ;
        RECT 81.045 88.115 81.335 88.160 ;
        RECT 81.965 88.115 82.255 88.345 ;
        RECT 66.400 87.820 68.930 87.960 ;
        RECT 68.610 87.760 68.930 87.820 ;
        RECT 72.310 87.960 72.600 88.005 ;
        RECT 74.170 87.960 74.460 88.005 ;
        RECT 72.310 87.820 74.460 87.960 ;
        RECT 72.310 87.775 72.600 87.820 ;
        RECT 74.170 87.775 74.460 87.820 ;
        RECT 75.090 87.960 75.380 88.005 ;
        RECT 76.890 87.960 77.210 88.020 ;
        RECT 78.350 87.960 78.640 88.005 ;
        RECT 75.090 87.820 78.640 87.960 ;
        RECT 75.090 87.775 75.380 87.820 ;
        RECT 76.890 87.760 77.210 87.820 ;
        RECT 78.350 87.775 78.640 87.820 ;
        RECT 58.490 87.620 58.810 87.680 ;
        RECT 45.700 87.480 58.810 87.620 ;
        RECT 30.430 87.420 30.750 87.480 ;
        RECT 30.905 87.435 31.195 87.480 ;
        RECT 32.730 87.420 33.050 87.480 ;
        RECT 44.690 87.420 45.010 87.480 ;
        RECT 45.165 87.435 45.455 87.480 ;
        RECT 58.490 87.420 58.810 87.480 ;
        RECT 76.430 87.620 76.750 87.680 ;
        RECT 80.355 87.620 80.645 87.665 ;
        RECT 82.040 87.620 82.180 88.115 ;
        RECT 82.410 88.100 82.730 88.360 ;
        RECT 82.870 88.100 83.190 88.360 ;
        RECT 85.720 88.345 85.860 88.840 ;
        RECT 86.180 88.345 86.320 89.180 ;
        RECT 88.405 89.180 89.170 89.320 ;
        RECT 88.405 89.135 88.695 89.180 ;
        RECT 88.850 89.120 89.170 89.180 ;
        RECT 89.770 89.120 90.090 89.380 ;
        RECT 91.165 89.320 91.455 89.365 ;
        RECT 91.610 89.320 91.930 89.380 ;
        RECT 91.165 89.180 91.930 89.320 ;
        RECT 91.165 89.135 91.455 89.180 ;
        RECT 91.610 89.120 91.930 89.180 ;
        RECT 92.530 89.120 92.850 89.380 ;
        RECT 93.450 89.320 93.770 89.380 ;
        RECT 96.225 89.320 96.515 89.365 ;
        RECT 93.450 89.180 96.515 89.320 ;
        RECT 93.450 89.120 93.770 89.180 ;
        RECT 96.225 89.135 96.515 89.180 ;
        RECT 97.130 89.320 97.450 89.380 ;
        RECT 101.730 89.320 102.050 89.380 ;
        RECT 97.130 89.180 102.050 89.320 ;
        RECT 97.130 89.120 97.450 89.180 ;
        RECT 101.730 89.120 102.050 89.180 ;
        RECT 98.050 88.980 98.370 89.040 ;
        RECT 103.590 88.980 103.880 89.025 ;
        RECT 105.450 88.980 105.740 89.025 ;
        RECT 108.230 88.980 108.520 89.025 ;
        RECT 98.050 88.840 102.420 88.980 ;
        RECT 98.050 88.780 98.370 88.840 ;
        RECT 98.600 88.685 98.740 88.840 ;
        RECT 102.280 88.685 102.420 88.840 ;
        RECT 103.590 88.840 108.520 88.980 ;
        RECT 103.590 88.795 103.880 88.840 ;
        RECT 105.450 88.795 105.740 88.840 ;
        RECT 108.230 88.795 108.520 88.840 ;
        RECT 109.550 88.980 109.870 89.040 ;
        RECT 114.165 88.980 114.455 89.025 ;
        RECT 109.550 88.840 114.455 88.980 ;
        RECT 109.550 88.780 109.870 88.840 ;
        RECT 114.165 88.795 114.455 88.840 ;
        RECT 87.945 88.640 88.235 88.685 ;
        RECT 87.945 88.500 93.680 88.640 ;
        RECT 87.945 88.455 88.235 88.500 ;
        RECT 84.725 88.300 85.015 88.345 ;
        RECT 83.420 88.160 85.015 88.300 ;
        RECT 83.420 87.960 83.560 88.160 ;
        RECT 84.725 88.115 85.015 88.160 ;
        RECT 85.645 88.115 85.935 88.345 ;
        RECT 86.105 88.115 86.395 88.345 ;
        RECT 86.550 88.100 86.870 88.360 ;
        RECT 89.310 88.100 89.630 88.360 ;
        RECT 89.785 88.300 90.075 88.345 ;
        RECT 90.230 88.300 90.550 88.360 ;
        RECT 89.785 88.160 90.550 88.300 ;
        RECT 89.785 88.115 90.075 88.160 ;
        RECT 90.230 88.100 90.550 88.160 ;
        RECT 92.070 88.100 92.390 88.360 ;
        RECT 92.530 88.100 92.850 88.360 ;
        RECT 93.540 88.345 93.680 88.500 ;
        RECT 98.525 88.455 98.815 88.685 ;
        RECT 99.445 88.640 99.735 88.685 ;
        RECT 99.445 88.500 101.960 88.640 ;
        RECT 99.445 88.455 99.735 88.500 ;
        RECT 101.820 88.360 101.960 88.500 ;
        RECT 102.205 88.455 102.495 88.685 ;
        RECT 104.030 88.640 104.350 88.700 ;
        RECT 104.965 88.640 105.255 88.685 ;
        RECT 110.930 88.640 111.250 88.700 ;
        RECT 102.740 88.500 103.800 88.640 ;
        RECT 93.465 88.115 93.755 88.345 ;
        RECT 98.065 88.300 98.355 88.345 ;
        RECT 100.350 88.300 100.670 88.360 ;
        RECT 98.065 88.160 100.670 88.300 ;
        RECT 98.065 88.115 98.355 88.160 ;
        RECT 100.350 88.100 100.670 88.160 ;
        RECT 100.810 88.300 101.130 88.360 ;
        RECT 101.285 88.300 101.575 88.345 ;
        RECT 100.810 88.160 101.575 88.300 ;
        RECT 100.810 88.100 101.130 88.160 ;
        RECT 101.285 88.115 101.575 88.160 ;
        RECT 101.730 88.300 102.050 88.360 ;
        RECT 102.740 88.300 102.880 88.500 ;
        RECT 101.730 88.160 102.880 88.300 ;
        RECT 101.730 88.100 102.050 88.160 ;
        RECT 103.110 88.100 103.430 88.360 ;
        RECT 103.660 88.300 103.800 88.500 ;
        RECT 104.030 88.500 105.255 88.640 ;
        RECT 104.030 88.440 104.350 88.500 ;
        RECT 104.965 88.455 105.255 88.500 ;
        RECT 105.500 88.500 111.250 88.640 ;
        RECT 105.500 88.300 105.640 88.500 ;
        RECT 110.930 88.440 111.250 88.500 ;
        RECT 113.230 88.640 113.550 88.700 ;
        RECT 113.230 88.500 115.760 88.640 ;
        RECT 113.230 88.440 113.550 88.500 ;
        RECT 108.230 88.300 108.520 88.345 ;
        RECT 103.660 88.160 105.640 88.300 ;
        RECT 105.985 88.160 108.520 88.300 ;
        RECT 113.320 88.300 113.460 88.440 ;
        RECT 113.705 88.300 113.995 88.345 ;
        RECT 113.320 88.160 113.995 88.300 ;
        RECT 82.500 87.820 83.560 87.960 ;
        RECT 84.265 87.960 84.555 88.005 ;
        RECT 90.705 87.960 90.995 88.005 ;
        RECT 84.265 87.820 90.995 87.960 ;
        RECT 82.500 87.680 82.640 87.820 ;
        RECT 84.265 87.775 84.555 87.820 ;
        RECT 90.705 87.775 90.995 87.820 ;
        RECT 96.670 87.960 96.990 88.020 ;
        RECT 103.200 87.960 103.340 88.100 ;
        RECT 105.985 88.005 106.200 88.160 ;
        RECT 108.230 88.115 108.520 88.160 ;
        RECT 113.705 88.115 113.995 88.160 ;
        RECT 114.150 88.300 114.470 88.360 ;
        RECT 115.620 88.345 115.760 88.500 ;
        RECT 115.085 88.300 115.375 88.345 ;
        RECT 114.150 88.160 115.375 88.300 ;
        RECT 114.150 88.100 114.470 88.160 ;
        RECT 115.085 88.115 115.375 88.160 ;
        RECT 115.545 88.115 115.835 88.345 ;
        RECT 96.670 87.820 103.340 87.960 ;
        RECT 104.050 87.960 104.340 88.005 ;
        RECT 105.910 87.960 106.200 88.005 ;
        RECT 104.050 87.820 106.200 87.960 ;
        RECT 96.670 87.760 96.990 87.820 ;
        RECT 104.050 87.775 104.340 87.820 ;
        RECT 105.910 87.775 106.200 87.820 ;
        RECT 106.830 87.960 107.120 88.005 ;
        RECT 110.090 87.960 110.380 88.005 ;
        RECT 113.245 87.960 113.535 88.005 ;
        RECT 116.005 87.960 116.295 88.005 ;
        RECT 106.830 87.820 113.535 87.960 ;
        RECT 106.830 87.775 107.120 87.820 ;
        RECT 110.090 87.775 110.380 87.820 ;
        RECT 113.245 87.775 113.535 87.820 ;
        RECT 113.780 87.820 116.295 87.960 ;
        RECT 113.780 87.680 113.920 87.820 ;
        RECT 116.005 87.775 116.295 87.820 ;
        RECT 76.430 87.480 82.180 87.620 ;
        RECT 76.430 87.420 76.750 87.480 ;
        RECT 80.355 87.435 80.645 87.480 ;
        RECT 82.410 87.420 82.730 87.680 ;
        RECT 98.970 87.620 99.290 87.680 ;
        RECT 100.365 87.620 100.655 87.665 ;
        RECT 98.970 87.480 100.655 87.620 ;
        RECT 98.970 87.420 99.290 87.480 ;
        RECT 100.365 87.435 100.655 87.480 ;
        RECT 110.930 87.620 111.250 87.680 ;
        RECT 112.095 87.620 112.385 87.665 ;
        RECT 110.930 87.480 112.385 87.620 ;
        RECT 110.930 87.420 111.250 87.480 ;
        RECT 112.095 87.435 112.385 87.480 ;
        RECT 113.690 87.420 114.010 87.680 ;
        RECT 5.520 86.800 118.680 87.280 ;
        RECT 19.850 86.400 20.170 86.660 ;
        RECT 26.305 86.415 26.595 86.645 ;
        RECT 17.090 86.305 17.410 86.320 ;
        RECT 11.130 86.260 11.420 86.305 ;
        RECT 12.990 86.260 13.280 86.305 ;
        RECT 11.130 86.120 13.280 86.260 ;
        RECT 11.130 86.075 11.420 86.120 ;
        RECT 12.990 86.075 13.280 86.120 ;
        RECT 13.910 86.260 14.200 86.305 ;
        RECT 17.090 86.260 17.460 86.305 ;
        RECT 13.910 86.120 17.460 86.260 ;
        RECT 13.910 86.075 14.200 86.120 ;
        RECT 17.090 86.075 17.460 86.120 ;
        RECT 19.175 86.260 19.465 86.305 ;
        RECT 22.165 86.260 22.455 86.305 ;
        RECT 23.990 86.260 24.310 86.320 ;
        RECT 19.175 86.120 24.310 86.260 ;
        RECT 19.175 86.075 19.465 86.120 ;
        RECT 22.165 86.075 22.455 86.120 ;
        RECT 9.745 85.735 10.035 85.965 ;
        RECT 8.810 84.700 9.130 84.960 ;
        RECT 9.820 84.900 9.960 85.735 ;
        RECT 12.030 85.720 12.350 85.980 ;
        RECT 13.065 85.920 13.280 86.075 ;
        RECT 17.090 86.060 17.410 86.075 ;
        RECT 23.990 86.060 24.310 86.120 ;
        RECT 15.310 85.920 15.600 85.965 ;
        RECT 13.065 85.780 15.600 85.920 ;
        RECT 15.310 85.735 15.600 85.780 ;
        RECT 20.310 85.920 20.630 85.980 ;
        RECT 21.705 85.920 21.995 85.965 ;
        RECT 20.310 85.780 21.995 85.920 ;
        RECT 20.310 85.720 20.630 85.780 ;
        RECT 21.705 85.735 21.995 85.780 ;
        RECT 10.205 85.580 10.495 85.625 ;
        RECT 11.570 85.580 11.890 85.640 ;
        RECT 10.205 85.440 11.890 85.580 ;
        RECT 10.205 85.395 10.495 85.440 ;
        RECT 11.570 85.380 11.890 85.440 ;
        RECT 23.085 85.395 23.375 85.625 ;
        RECT 24.080 85.580 24.220 86.060 ;
        RECT 24.925 85.920 25.215 85.965 ;
        RECT 26.380 85.920 26.520 86.415 ;
        RECT 31.810 86.400 32.130 86.660 ;
        RECT 37.805 86.600 38.095 86.645 ;
        RECT 34.200 86.460 38.095 86.600 ;
        RECT 34.200 86.260 34.340 86.460 ;
        RECT 37.805 86.415 38.095 86.460 ;
        RECT 39.170 86.600 39.490 86.660 ;
        RECT 39.645 86.600 39.935 86.645 ;
        RECT 39.170 86.460 39.935 86.600 ;
        RECT 39.170 86.400 39.490 86.460 ;
        RECT 39.645 86.415 39.935 86.460 ;
        RECT 40.090 86.600 40.410 86.660 ;
        RECT 47.910 86.600 48.230 86.660 ;
        RECT 40.090 86.460 48.230 86.600 ;
        RECT 40.090 86.400 40.410 86.460 ;
        RECT 47.910 86.400 48.230 86.460 ;
        RECT 52.985 86.600 53.275 86.645 ;
        RECT 53.890 86.600 54.210 86.660 ;
        RECT 71.830 86.600 72.150 86.660 ;
        RECT 52.985 86.460 54.210 86.600 ;
        RECT 52.985 86.415 53.275 86.460 ;
        RECT 53.890 86.400 54.210 86.460 ;
        RECT 63.180 86.460 72.150 86.600 ;
        RECT 32.360 86.120 34.340 86.260 ;
        RECT 24.925 85.780 26.520 85.920 ;
        RECT 24.925 85.735 25.215 85.780 ;
        RECT 28.145 85.735 28.435 85.965 ;
        RECT 28.605 85.920 28.895 85.965 ;
        RECT 32.360 85.920 32.500 86.120 ;
        RECT 34.200 85.980 34.340 86.120 ;
        RECT 34.570 86.260 34.890 86.320 ;
        RECT 38.710 86.260 39.030 86.320 ;
        RECT 41.030 86.260 41.320 86.305 ;
        RECT 42.890 86.260 43.180 86.305 ;
        RECT 34.570 86.120 40.320 86.260 ;
        RECT 34.570 86.060 34.890 86.120 ;
        RECT 38.710 86.060 39.030 86.120 ;
        RECT 28.605 85.780 32.500 85.920 ;
        RECT 32.730 85.920 33.050 85.980 ;
        RECT 33.205 85.920 33.495 85.965 ;
        RECT 32.730 85.780 33.495 85.920 ;
        RECT 28.605 85.735 28.895 85.780 ;
        RECT 28.220 85.580 28.360 85.735 ;
        RECT 32.730 85.720 33.050 85.780 ;
        RECT 33.205 85.735 33.495 85.780 ;
        RECT 33.650 85.720 33.970 85.980 ;
        RECT 34.110 85.720 34.430 85.980 ;
        RECT 35.030 85.920 35.350 85.980 ;
        RECT 39.630 85.920 39.950 85.980 ;
        RECT 40.180 85.965 40.320 86.120 ;
        RECT 41.030 86.120 43.180 86.260 ;
        RECT 41.030 86.075 41.320 86.120 ;
        RECT 42.890 86.075 43.180 86.120 ;
        RECT 43.810 86.260 44.100 86.305 ;
        RECT 44.690 86.260 45.010 86.320 ;
        RECT 47.070 86.260 47.360 86.305 ;
        RECT 43.810 86.120 47.360 86.260 ;
        RECT 43.810 86.075 44.100 86.120 ;
        RECT 35.030 85.780 39.950 85.920 ;
        RECT 35.030 85.720 35.350 85.780 ;
        RECT 39.630 85.720 39.950 85.780 ;
        RECT 40.105 85.735 40.395 85.965 ;
        RECT 42.965 85.920 43.180 86.075 ;
        RECT 44.690 86.060 45.010 86.120 ;
        RECT 47.070 86.075 47.360 86.120 ;
        RECT 48.830 86.260 49.150 86.320 ;
        RECT 63.180 86.260 63.320 86.460 ;
        RECT 71.830 86.400 72.150 86.460 ;
        RECT 73.210 86.600 73.530 86.660 ;
        RECT 74.145 86.600 74.435 86.645 ;
        RECT 73.210 86.460 74.435 86.600 ;
        RECT 73.210 86.400 73.530 86.460 ;
        RECT 74.145 86.415 74.435 86.460 ;
        RECT 75.985 86.415 76.275 86.645 ;
        RECT 76.430 86.600 76.750 86.660 ;
        RECT 78.285 86.600 78.575 86.645 ;
        RECT 76.430 86.460 78.575 86.600 ;
        RECT 48.830 86.120 54.580 86.260 ;
        RECT 48.830 86.060 49.150 86.120 ;
        RECT 45.210 85.920 45.500 85.965 ;
        RECT 42.965 85.780 45.500 85.920 ;
        RECT 45.210 85.735 45.500 85.780 ;
        RECT 49.750 85.720 50.070 85.980 ;
        RECT 50.685 85.735 50.975 85.965 ;
        RECT 51.145 85.735 51.435 85.965 ;
        RECT 24.080 85.440 28.360 85.580 ;
        RECT 29.525 85.580 29.815 85.625 ;
        RECT 36.885 85.580 37.175 85.625 ;
        RECT 29.525 85.440 37.175 85.580 ;
        RECT 29.525 85.395 29.815 85.440 ;
        RECT 36.885 85.395 37.175 85.440 ;
        RECT 37.345 85.580 37.635 85.625 ;
        RECT 41.470 85.580 41.790 85.640 ;
        RECT 37.345 85.440 41.790 85.580 ;
        RECT 37.345 85.395 37.635 85.440 ;
        RECT 10.670 85.240 10.960 85.285 ;
        RECT 12.530 85.240 12.820 85.285 ;
        RECT 15.310 85.240 15.600 85.285 ;
        RECT 10.670 85.100 15.600 85.240 ;
        RECT 10.670 85.055 10.960 85.100 ;
        RECT 12.530 85.055 12.820 85.100 ;
        RECT 15.310 85.055 15.600 85.100 ;
        RECT 19.850 85.240 20.170 85.300 ;
        RECT 23.160 85.240 23.300 85.395 ;
        RECT 29.600 85.240 29.740 85.395 ;
        RECT 19.850 85.100 29.740 85.240 ;
        RECT 36.960 85.240 37.100 85.395 ;
        RECT 41.470 85.380 41.790 85.440 ;
        RECT 41.930 85.380 42.250 85.640 ;
        RECT 46.530 85.580 46.850 85.640 ;
        RECT 50.760 85.580 50.900 85.735 ;
        RECT 46.530 85.440 50.900 85.580 ;
        RECT 46.530 85.380 46.850 85.440 ;
        RECT 40.570 85.240 40.860 85.285 ;
        RECT 42.430 85.240 42.720 85.285 ;
        RECT 45.210 85.240 45.500 85.285 ;
        RECT 36.960 85.100 37.560 85.240 ;
        RECT 19.850 85.040 20.170 85.100 ;
        RECT 13.410 84.900 13.730 84.960 ;
        RECT 9.820 84.760 13.730 84.900 ;
        RECT 13.410 84.700 13.730 84.760 ;
        RECT 25.845 84.900 26.135 84.945 ;
        RECT 27.670 84.900 27.990 84.960 ;
        RECT 25.845 84.760 27.990 84.900 ;
        RECT 37.420 84.900 37.560 85.100 ;
        RECT 40.570 85.100 45.500 85.240 ;
        RECT 40.570 85.055 40.860 85.100 ;
        RECT 42.430 85.055 42.720 85.100 ;
        RECT 45.210 85.055 45.500 85.100 ;
        RECT 46.070 85.240 46.390 85.300 ;
        RECT 50.670 85.240 50.990 85.300 ;
        RECT 51.220 85.240 51.360 85.735 ;
        RECT 51.590 85.720 51.910 85.980 ;
        RECT 53.430 85.720 53.750 85.980 ;
        RECT 54.440 85.965 54.580 86.120 ;
        RECT 62.720 86.120 63.320 86.260 ;
        RECT 66.310 86.260 66.630 86.320 ;
        RECT 67.690 86.260 68.010 86.320 ;
        RECT 72.290 86.260 72.610 86.320 ;
        RECT 66.310 86.120 69.300 86.260 ;
        RECT 54.365 85.735 54.655 85.965 ;
        RECT 54.825 85.920 55.115 85.965 ;
        RECT 56.650 85.920 56.970 85.980 ;
        RECT 62.720 85.965 62.860 86.120 ;
        RECT 66.310 86.060 66.630 86.120 ;
        RECT 67.690 86.060 68.010 86.120 ;
        RECT 54.825 85.780 56.970 85.920 ;
        RECT 54.825 85.735 55.115 85.780 ;
        RECT 56.650 85.720 56.970 85.780 ;
        RECT 62.645 85.735 62.935 85.965 ;
        RECT 63.105 85.735 63.395 85.965 ;
        RECT 58.950 85.580 59.270 85.640 ;
        RECT 63.180 85.580 63.320 85.735 ;
        RECT 63.550 85.720 63.870 85.980 ;
        RECT 64.485 85.920 64.775 85.965 ;
        RECT 64.945 85.920 65.235 85.965 ;
        RECT 64.485 85.780 65.235 85.920 ;
        RECT 64.485 85.735 64.775 85.780 ;
        RECT 64.945 85.735 65.235 85.780 ;
        RECT 68.610 85.720 68.930 85.980 ;
        RECT 58.950 85.440 63.320 85.580 ;
        RECT 67.230 85.580 67.550 85.640 ;
        RECT 67.705 85.580 67.995 85.625 ;
        RECT 67.230 85.440 67.995 85.580 ;
        RECT 69.160 85.580 69.300 86.120 ;
        RECT 69.620 86.120 72.610 86.260 ;
        RECT 69.620 85.965 69.760 86.120 ;
        RECT 72.290 86.060 72.610 86.120 ;
        RECT 69.545 85.735 69.835 85.965 ;
        RECT 70.005 85.735 70.295 85.965 ;
        RECT 70.465 85.735 70.755 85.965 ;
        RECT 75.065 85.920 75.355 85.965 ;
        RECT 76.060 85.920 76.200 86.415 ;
        RECT 76.430 86.400 76.750 86.460 ;
        RECT 78.285 86.415 78.575 86.460 ;
        RECT 81.030 86.600 81.350 86.660 ;
        RECT 89.325 86.600 89.615 86.645 ;
        RECT 81.030 86.460 89.615 86.600 ;
        RECT 81.030 86.400 81.350 86.460 ;
        RECT 89.325 86.415 89.615 86.460 ;
        RECT 94.370 86.600 94.690 86.660 ;
        RECT 95.305 86.600 95.595 86.645 ;
        RECT 94.370 86.460 95.595 86.600 ;
        RECT 94.370 86.400 94.690 86.460 ;
        RECT 95.305 86.415 95.595 86.460 ;
        RECT 98.065 86.600 98.355 86.645 ;
        RECT 98.510 86.600 98.830 86.660 ;
        RECT 98.065 86.460 98.830 86.600 ;
        RECT 98.065 86.415 98.355 86.460 ;
        RECT 98.510 86.400 98.830 86.460 ;
        RECT 100.350 86.600 100.670 86.660 ;
        RECT 102.190 86.600 102.510 86.660 ;
        RECT 100.350 86.460 102.510 86.600 ;
        RECT 100.350 86.400 100.670 86.460 ;
        RECT 102.190 86.400 102.510 86.460 ;
        RECT 104.490 86.400 104.810 86.660 ;
        RECT 110.485 86.600 110.775 86.645 ;
        RECT 110.930 86.600 111.250 86.660 ;
        RECT 110.485 86.460 111.250 86.600 ;
        RECT 110.485 86.415 110.775 86.460 ;
        RECT 77.350 86.260 77.670 86.320 ;
        RECT 80.570 86.260 80.890 86.320 ;
        RECT 82.410 86.260 82.730 86.320 ;
        RECT 83.790 86.260 84.110 86.320 ;
        RECT 86.565 86.260 86.855 86.305 ;
        RECT 87.025 86.260 87.315 86.305 ;
        RECT 95.765 86.260 96.055 86.305 ;
        RECT 77.350 86.120 83.560 86.260 ;
        RECT 77.350 86.060 77.670 86.120 ;
        RECT 80.570 86.060 80.890 86.120 ;
        RECT 82.410 86.060 82.730 86.120 ;
        RECT 83.420 85.965 83.560 86.120 ;
        RECT 83.790 86.120 85.860 86.260 ;
        RECT 83.790 86.060 84.110 86.120 ;
        RECT 75.065 85.780 76.200 85.920 ;
        RECT 77.825 85.920 78.115 85.965 ;
        RECT 77.825 85.780 82.640 85.920 ;
        RECT 75.065 85.735 75.355 85.780 ;
        RECT 77.825 85.735 78.115 85.780 ;
        RECT 70.080 85.580 70.220 85.735 ;
        RECT 69.160 85.440 70.220 85.580 ;
        RECT 58.950 85.380 59.270 85.440 ;
        RECT 67.230 85.380 67.550 85.440 ;
        RECT 67.705 85.395 67.995 85.440 ;
        RECT 55.745 85.240 56.035 85.285 ;
        RECT 46.070 85.100 50.440 85.240 ;
        RECT 46.070 85.040 46.390 85.100 ;
        RECT 47.910 84.900 48.230 84.960 ;
        RECT 37.420 84.760 48.230 84.900 ;
        RECT 25.845 84.715 26.135 84.760 ;
        RECT 27.670 84.700 27.990 84.760 ;
        RECT 47.910 84.700 48.230 84.760 ;
        RECT 48.370 84.900 48.690 84.960 ;
        RECT 49.075 84.900 49.365 84.945 ;
        RECT 48.370 84.760 49.365 84.900 ;
        RECT 50.300 84.900 50.440 85.100 ;
        RECT 50.670 85.100 51.360 85.240 ;
        RECT 51.680 85.100 56.035 85.240 ;
        RECT 50.670 85.040 50.990 85.100 ;
        RECT 51.680 84.900 51.820 85.100 ;
        RECT 55.745 85.055 56.035 85.100 ;
        RECT 58.490 85.240 58.810 85.300 ;
        RECT 70.540 85.240 70.680 85.735 ;
        RECT 82.500 85.640 82.640 85.780 ;
        RECT 83.345 85.735 83.635 85.965 ;
        RECT 84.265 85.735 84.555 85.965 ;
        RECT 78.270 85.580 78.590 85.640 ;
        RECT 78.745 85.580 79.035 85.625 ;
        RECT 78.270 85.440 79.035 85.580 ;
        RECT 78.270 85.380 78.590 85.440 ;
        RECT 78.745 85.395 79.035 85.440 ;
        RECT 82.410 85.580 82.730 85.640 ;
        RECT 84.340 85.580 84.480 85.735 ;
        RECT 84.710 85.720 85.030 85.980 ;
        RECT 85.170 85.720 85.490 85.980 ;
        RECT 85.720 85.920 85.860 86.120 ;
        RECT 86.565 86.120 87.315 86.260 ;
        RECT 86.565 86.075 86.855 86.120 ;
        RECT 87.025 86.075 87.315 86.120 ;
        RECT 87.560 86.120 96.055 86.260 ;
        RECT 87.560 85.920 87.700 86.120 ;
        RECT 95.765 86.075 96.055 86.120 ;
        RECT 85.720 85.780 87.700 85.920 ;
        RECT 88.405 85.920 88.695 85.965 ;
        RECT 90.690 85.920 91.010 85.980 ;
        RECT 88.405 85.780 91.010 85.920 ;
        RECT 88.405 85.735 88.695 85.780 ;
        RECT 90.690 85.720 91.010 85.780 ;
        RECT 93.005 85.735 93.295 85.965 ;
        RECT 82.410 85.440 84.480 85.580 ;
        RECT 82.410 85.380 82.730 85.440 ;
        RECT 87.470 85.380 87.790 85.640 ;
        RECT 58.490 85.100 70.680 85.240 ;
        RECT 58.490 85.040 58.810 85.100 ;
        RECT 67.780 84.960 67.920 85.100 ;
        RECT 50.300 84.760 51.820 84.900 ;
        RECT 52.970 84.900 53.290 84.960 ;
        RECT 53.445 84.900 53.735 84.945 ;
        RECT 52.970 84.760 53.735 84.900 ;
        RECT 48.370 84.700 48.690 84.760 ;
        RECT 49.075 84.715 49.365 84.760 ;
        RECT 52.970 84.700 53.290 84.760 ;
        RECT 53.445 84.715 53.735 84.760 ;
        RECT 58.030 84.900 58.350 84.960 ;
        RECT 61.725 84.900 62.015 84.945 ;
        RECT 58.030 84.760 62.015 84.900 ;
        RECT 58.030 84.700 58.350 84.760 ;
        RECT 61.725 84.715 62.015 84.760 ;
        RECT 67.690 84.700 68.010 84.960 ;
        RECT 70.540 84.900 70.680 85.100 ;
        RECT 71.845 85.240 72.135 85.285 ;
        RECT 93.080 85.240 93.220 85.735 ;
        RECT 94.370 85.720 94.690 85.980 ;
        RECT 96.210 85.920 96.530 85.980 ;
        RECT 97.145 85.920 97.435 85.965 ;
        RECT 96.210 85.780 97.435 85.920 ;
        RECT 96.210 85.720 96.530 85.780 ;
        RECT 97.145 85.735 97.435 85.780 ;
        RECT 98.050 85.920 98.370 85.980 ;
        RECT 99.430 85.920 99.750 85.980 ;
        RECT 100.440 85.965 100.580 86.400 ;
        RECT 102.650 86.260 102.970 86.320 ;
        RECT 110.560 86.260 110.700 86.415 ;
        RECT 110.930 86.400 111.250 86.460 ;
        RECT 112.785 86.600 113.075 86.645 ;
        RECT 114.150 86.600 114.470 86.660 ;
        RECT 112.785 86.460 114.470 86.600 ;
        RECT 112.785 86.415 113.075 86.460 ;
        RECT 114.150 86.400 114.470 86.460 ;
        RECT 102.650 86.120 110.700 86.260 ;
        RECT 102.650 86.060 102.970 86.120 ;
        RECT 98.050 85.780 99.750 85.920 ;
        RECT 98.050 85.720 98.370 85.780 ;
        RECT 99.430 85.720 99.750 85.780 ;
        RECT 100.365 85.735 100.655 85.965 ;
        RECT 110.470 85.920 110.790 85.980 ;
        RECT 110.945 85.920 111.235 85.965 ;
        RECT 110.470 85.780 111.235 85.920 ;
        RECT 110.470 85.720 110.790 85.780 ;
        RECT 110.945 85.735 111.235 85.780 ;
        RECT 93.910 85.380 94.230 85.640 ;
        RECT 96.685 85.580 96.975 85.625 ;
        RECT 97.590 85.580 97.910 85.640 ;
        RECT 96.685 85.440 97.910 85.580 ;
        RECT 96.685 85.395 96.975 85.440 ;
        RECT 97.590 85.380 97.910 85.440 ;
        RECT 101.730 85.380 102.050 85.640 ;
        RECT 110.025 85.580 110.315 85.625 ;
        RECT 111.390 85.580 111.710 85.640 ;
        RECT 110.025 85.440 111.710 85.580 ;
        RECT 110.025 85.395 110.315 85.440 ;
        RECT 111.390 85.380 111.710 85.440 ;
        RECT 98.970 85.240 99.290 85.300 ;
        RECT 71.845 85.100 93.220 85.240 ;
        RECT 97.220 85.100 99.290 85.240 ;
        RECT 71.845 85.055 72.135 85.100 ;
        RECT 72.290 84.900 72.610 84.960 ;
        RECT 70.540 84.760 72.610 84.900 ;
        RECT 72.290 84.700 72.610 84.760 ;
        RECT 79.650 84.900 79.970 84.960 ;
        RECT 81.950 84.900 82.270 84.960 ;
        RECT 84.710 84.900 85.030 84.960 ;
        RECT 79.650 84.760 85.030 84.900 ;
        RECT 79.650 84.700 79.970 84.760 ;
        RECT 81.950 84.700 82.270 84.760 ;
        RECT 84.710 84.700 85.030 84.760 ;
        RECT 88.390 84.700 88.710 84.960 ;
        RECT 94.385 84.900 94.675 84.945 ;
        RECT 94.830 84.900 95.150 84.960 ;
        RECT 97.220 84.945 97.360 85.100 ;
        RECT 98.970 85.040 99.290 85.100 ;
        RECT 94.385 84.760 95.150 84.900 ;
        RECT 94.385 84.715 94.675 84.760 ;
        RECT 94.830 84.700 95.150 84.760 ;
        RECT 97.145 84.715 97.435 84.945 ;
        RECT 98.510 84.700 98.830 84.960 ;
        RECT 5.520 84.080 118.680 84.560 ;
        RECT 8.350 83.880 8.670 83.940 ;
        RECT 11.570 83.880 11.890 83.940 ;
        RECT 34.570 83.880 34.890 83.940 ;
        RECT 7.060 83.740 34.890 83.880 ;
        RECT 7.060 83.260 7.200 83.740 ;
        RECT 8.350 83.680 8.670 83.740 ;
        RECT 11.570 83.680 11.890 83.740 ;
        RECT 7.450 83.540 7.740 83.585 ;
        RECT 9.310 83.540 9.600 83.585 ;
        RECT 12.090 83.540 12.380 83.585 ;
        RECT 7.450 83.400 12.380 83.540 ;
        RECT 7.450 83.355 7.740 83.400 ;
        RECT 9.310 83.355 9.600 83.400 ;
        RECT 12.090 83.355 12.380 83.400 ;
        RECT 12.950 83.540 13.270 83.600 ;
        RECT 20.310 83.540 20.630 83.600 ;
        RECT 12.950 83.400 17.780 83.540 ;
        RECT 12.950 83.340 13.270 83.400 ;
        RECT 6.970 83.000 7.290 83.260 ;
        RECT 8.810 82.660 9.130 82.920 ;
        RECT 12.090 82.860 12.380 82.905 ;
        RECT 9.845 82.720 12.380 82.860 ;
        RECT 9.845 82.565 10.060 82.720 ;
        RECT 12.090 82.675 12.380 82.720 ;
        RECT 17.090 82.660 17.410 82.920 ;
        RECT 17.640 82.905 17.780 83.400 ;
        RECT 19.020 83.400 22.840 83.540 ;
        RECT 17.565 82.675 17.855 82.905 ;
        RECT 7.910 82.520 8.200 82.565 ;
        RECT 9.770 82.520 10.060 82.565 ;
        RECT 7.910 82.380 10.060 82.520 ;
        RECT 7.910 82.335 8.200 82.380 ;
        RECT 9.770 82.335 10.060 82.380 ;
        RECT 10.690 82.520 10.980 82.565 ;
        RECT 12.490 82.520 12.810 82.580 ;
        RECT 15.710 82.565 16.030 82.580 ;
        RECT 13.950 82.520 14.240 82.565 ;
        RECT 10.690 82.380 14.240 82.520 ;
        RECT 10.690 82.335 10.980 82.380 ;
        RECT 12.490 82.320 12.810 82.380 ;
        RECT 13.950 82.335 14.240 82.380 ;
        RECT 15.710 82.520 16.245 82.565 ;
        RECT 19.020 82.520 19.160 83.400 ;
        RECT 20.310 83.340 20.630 83.400 ;
        RECT 20.400 83.060 21.920 83.200 ;
        RECT 20.400 82.920 20.540 83.060 ;
        RECT 20.310 82.660 20.630 82.920 ;
        RECT 21.780 82.905 21.920 83.060 ;
        RECT 21.245 82.675 21.535 82.905 ;
        RECT 21.705 82.675 21.995 82.905 ;
        RECT 22.165 82.870 22.455 82.890 ;
        RECT 22.700 82.870 22.840 83.400 ;
        RECT 25.920 83.245 26.060 83.740 ;
        RECT 34.570 83.680 34.890 83.740 ;
        RECT 41.930 83.880 42.250 83.940 ;
        RECT 42.865 83.880 43.155 83.925 ;
        RECT 41.930 83.740 43.155 83.880 ;
        RECT 41.930 83.680 42.250 83.740 ;
        RECT 42.865 83.695 43.155 83.740 ;
        RECT 53.430 83.680 53.750 83.940 ;
        RECT 66.310 83.880 66.630 83.940 ;
        RECT 79.190 83.880 79.510 83.940 ;
        RECT 82.870 83.880 83.190 83.940 ;
        RECT 85.170 83.880 85.490 83.940 ;
        RECT 65.020 83.740 72.060 83.880 ;
        RECT 26.310 83.540 26.600 83.585 ;
        RECT 28.170 83.540 28.460 83.585 ;
        RECT 30.950 83.540 31.240 83.585 ;
        RECT 26.310 83.400 31.240 83.540 ;
        RECT 26.310 83.355 26.600 83.400 ;
        RECT 28.170 83.355 28.460 83.400 ;
        RECT 30.950 83.355 31.240 83.400 ;
        RECT 38.710 83.540 39.030 83.600 ;
        RECT 56.670 83.540 56.960 83.585 ;
        RECT 58.530 83.540 58.820 83.585 ;
        RECT 61.310 83.540 61.600 83.585 ;
        RECT 38.710 83.400 56.420 83.540 ;
        RECT 38.710 83.340 39.030 83.400 ;
        RECT 25.845 83.015 26.135 83.245 ;
        RECT 27.670 83.000 27.990 83.260 ;
        RECT 34.110 83.200 34.430 83.260 ;
        RECT 34.815 83.200 35.105 83.245 ;
        RECT 34.110 83.060 35.105 83.200 ;
        RECT 34.110 83.000 34.430 83.060 ;
        RECT 34.815 83.015 35.105 83.060 ;
        RECT 47.910 83.000 48.230 83.260 ;
        RECT 49.750 83.200 50.070 83.260 ;
        RECT 50.670 83.200 50.990 83.260 ;
        RECT 56.280 83.245 56.420 83.400 ;
        RECT 56.670 83.400 61.600 83.540 ;
        RECT 56.670 83.355 56.960 83.400 ;
        RECT 58.530 83.355 58.820 83.400 ;
        RECT 61.310 83.355 61.600 83.400 ;
        RECT 49.750 83.060 50.440 83.200 ;
        RECT 49.750 83.000 50.070 83.060 ;
        RECT 22.165 82.730 22.840 82.870 ;
        RECT 23.085 82.860 23.375 82.905 ;
        RECT 23.530 82.860 23.850 82.920 ;
        RECT 30.950 82.860 31.240 82.905 ;
        RECT 15.710 82.380 19.160 82.520 ;
        RECT 19.865 82.520 20.155 82.565 ;
        RECT 20.770 82.520 21.090 82.580 ;
        RECT 19.865 82.380 21.090 82.520 ;
        RECT 21.320 82.520 21.460 82.675 ;
        RECT 22.165 82.660 22.455 82.730 ;
        RECT 23.085 82.720 23.850 82.860 ;
        RECT 23.085 82.675 23.375 82.720 ;
        RECT 23.530 82.660 23.850 82.720 ;
        RECT 28.705 82.720 31.240 82.860 ;
        RECT 22.610 82.520 22.930 82.580 ;
        RECT 28.705 82.565 28.920 82.720 ;
        RECT 30.950 82.675 31.240 82.720 ;
        RECT 43.785 82.860 44.075 82.905 ;
        RECT 43.785 82.720 44.920 82.860 ;
        RECT 43.785 82.675 44.075 82.720 ;
        RECT 21.320 82.380 22.930 82.520 ;
        RECT 15.710 82.335 16.245 82.380 ;
        RECT 19.865 82.335 20.155 82.380 ;
        RECT 15.710 82.320 16.030 82.335 ;
        RECT 20.770 82.320 21.090 82.380 ;
        RECT 22.610 82.320 22.930 82.380 ;
        RECT 26.770 82.520 27.060 82.565 ;
        RECT 28.630 82.520 28.920 82.565 ;
        RECT 26.770 82.380 28.920 82.520 ;
        RECT 26.770 82.335 27.060 82.380 ;
        RECT 28.630 82.335 28.920 82.380 ;
        RECT 29.550 82.520 29.840 82.565 ;
        RECT 30.430 82.520 30.750 82.580 ;
        RECT 32.810 82.520 33.100 82.565 ;
        RECT 29.550 82.380 33.100 82.520 ;
        RECT 29.550 82.335 29.840 82.380 ;
        RECT 30.430 82.320 30.750 82.380 ;
        RECT 32.810 82.335 33.100 82.380 ;
        RECT 44.780 82.225 44.920 82.720 ;
        RECT 46.530 82.660 46.850 82.920 ;
        RECT 50.300 82.905 50.440 83.060 ;
        RECT 50.670 83.060 51.820 83.200 ;
        RECT 50.670 83.000 50.990 83.060 ;
        RECT 51.680 82.905 51.820 83.060 ;
        RECT 56.205 83.015 56.495 83.245 ;
        RECT 58.030 83.000 58.350 83.260 ;
        RECT 62.630 83.200 62.950 83.260 ;
        RECT 65.020 83.200 65.160 83.740 ;
        RECT 66.310 83.680 66.630 83.740 ;
        RECT 65.390 83.540 65.710 83.600 ;
        RECT 68.610 83.540 68.930 83.600 ;
        RECT 65.390 83.400 70.680 83.540 ;
        RECT 65.390 83.340 65.710 83.400 ;
        RECT 68.610 83.340 68.930 83.400 ;
        RECT 62.630 83.060 67.460 83.200 ;
        RECT 62.630 83.000 62.950 83.060 ;
        RECT 50.225 82.675 50.515 82.905 ;
        RECT 51.145 82.675 51.435 82.905 ;
        RECT 51.605 82.675 51.895 82.905 ;
        RECT 52.065 82.675 52.355 82.905 ;
        RECT 61.310 82.860 61.600 82.905 ;
        RECT 59.065 82.720 61.600 82.860 ;
        RECT 51.220 82.520 51.360 82.675 ;
        RECT 52.140 82.520 52.280 82.675 ;
        RECT 52.970 82.520 53.290 82.580 ;
        RECT 59.065 82.565 59.280 82.720 ;
        RECT 61.310 82.675 61.600 82.720 ;
        RECT 64.930 82.860 65.250 82.920 ;
        RECT 65.865 82.860 66.155 82.905 ;
        RECT 64.930 82.720 66.155 82.860 ;
        RECT 64.930 82.660 65.250 82.720 ;
        RECT 65.865 82.675 66.155 82.720 ;
        RECT 66.770 82.660 67.090 82.920 ;
        RECT 67.320 82.905 67.460 83.060 ;
        RECT 67.245 82.675 67.535 82.905 ;
        RECT 67.690 82.660 68.010 82.920 ;
        RECT 70.540 82.905 70.680 83.400 ;
        RECT 71.920 82.905 72.060 83.740 ;
        RECT 79.190 83.740 85.490 83.880 ;
        RECT 79.190 83.680 79.510 83.740 ;
        RECT 82.870 83.680 83.190 83.740 ;
        RECT 85.170 83.680 85.490 83.740 ;
        RECT 93.465 83.880 93.755 83.925 ;
        RECT 98.510 83.880 98.830 83.940 ;
        RECT 93.465 83.740 98.830 83.880 ;
        RECT 93.465 83.695 93.755 83.740 ;
        RECT 98.510 83.680 98.830 83.740 ;
        RECT 110.470 83.880 110.790 83.940 ;
        RECT 116.695 83.880 116.985 83.925 ;
        RECT 110.470 83.740 116.985 83.880 ;
        RECT 110.470 83.680 110.790 83.740 ;
        RECT 116.695 83.695 116.985 83.740 ;
        RECT 108.190 83.540 108.480 83.585 ;
        RECT 110.050 83.540 110.340 83.585 ;
        RECT 112.830 83.540 113.120 83.585 ;
        RECT 108.190 83.400 113.120 83.540 ;
        RECT 108.190 83.355 108.480 83.400 ;
        RECT 110.050 83.355 110.340 83.400 ;
        RECT 112.830 83.355 113.120 83.400 ;
        RECT 77.810 83.200 78.130 83.260 ;
        RECT 77.440 83.060 78.130 83.200 ;
        RECT 70.465 82.675 70.755 82.905 ;
        RECT 71.385 82.675 71.675 82.905 ;
        RECT 71.845 82.675 72.135 82.905 ;
        RECT 48.460 82.380 51.360 82.520 ;
        RECT 51.680 82.380 53.290 82.520 ;
        RECT 48.460 82.240 48.600 82.380 ;
        RECT 51.680 82.240 51.820 82.380 ;
        RECT 52.970 82.320 53.290 82.380 ;
        RECT 57.130 82.520 57.420 82.565 ;
        RECT 58.990 82.520 59.280 82.565 ;
        RECT 57.130 82.380 59.280 82.520 ;
        RECT 57.130 82.335 57.420 82.380 ;
        RECT 58.990 82.335 59.280 82.380 ;
        RECT 59.910 82.520 60.200 82.565 ;
        RECT 60.790 82.520 61.110 82.580 ;
        RECT 63.170 82.520 63.460 82.565 ;
        RECT 71.460 82.520 71.600 82.675 ;
        RECT 72.290 82.660 72.610 82.920 ;
        RECT 76.890 82.660 77.210 82.920 ;
        RECT 77.440 82.905 77.580 83.060 ;
        RECT 77.810 83.000 78.130 83.060 ;
        RECT 92.990 83.000 93.310 83.260 ;
        RECT 98.985 83.200 99.275 83.245 ;
        RECT 102.650 83.200 102.970 83.260 ;
        RECT 98.985 83.060 102.970 83.200 ;
        RECT 98.985 83.015 99.275 83.060 ;
        RECT 102.650 83.000 102.970 83.060 ;
        RECT 103.110 83.200 103.430 83.260 ;
        RECT 107.725 83.200 108.015 83.245 ;
        RECT 103.110 83.060 108.015 83.200 ;
        RECT 103.110 83.000 103.430 83.060 ;
        RECT 107.725 83.015 108.015 83.060 ;
        RECT 109.550 83.000 109.870 83.260 ;
        RECT 77.365 82.675 77.655 82.905 ;
        RECT 93.465 82.860 93.755 82.905 ;
        RECT 97.130 82.860 97.450 82.920 ;
        RECT 98.050 82.860 98.370 82.920 ;
        RECT 112.830 82.860 113.120 82.905 ;
        RECT 77.900 82.720 93.755 82.860 ;
        RECT 77.900 82.520 78.040 82.720 ;
        RECT 93.465 82.675 93.755 82.720 ;
        RECT 96.530 82.720 97.450 82.860 ;
        RECT 97.855 82.720 98.370 82.860 ;
        RECT 59.910 82.380 63.460 82.520 ;
        RECT 59.910 82.335 60.200 82.380 ;
        RECT 60.790 82.320 61.110 82.380 ;
        RECT 63.170 82.335 63.460 82.380 ;
        RECT 67.320 82.380 71.600 82.520 ;
        RECT 73.300 82.380 78.040 82.520 ;
        RECT 91.610 82.520 91.930 82.580 ;
        RECT 92.085 82.520 92.375 82.565 ;
        RECT 96.530 82.520 96.670 82.720 ;
        RECT 97.130 82.660 97.450 82.720 ;
        RECT 98.050 82.660 98.370 82.720 ;
        RECT 110.585 82.720 113.120 82.860 ;
        RECT 110.585 82.565 110.800 82.720 ;
        RECT 112.830 82.675 113.120 82.720 ;
        RECT 91.610 82.380 92.375 82.520 ;
        RECT 67.320 82.240 67.460 82.380 ;
        RECT 44.705 81.995 44.995 82.225 ;
        RECT 47.005 82.180 47.295 82.225 ;
        RECT 48.370 82.180 48.690 82.240 ;
        RECT 47.005 82.040 48.690 82.180 ;
        RECT 47.005 81.995 47.295 82.040 ;
        RECT 48.370 81.980 48.690 82.040 ;
        RECT 51.590 81.980 51.910 82.240 ;
        RECT 65.175 82.180 65.465 82.225 ;
        RECT 67.230 82.180 67.550 82.240 ;
        RECT 65.175 82.040 67.550 82.180 ;
        RECT 65.175 81.995 65.465 82.040 ;
        RECT 67.230 81.980 67.550 82.040 ;
        RECT 69.085 82.180 69.375 82.225 ;
        RECT 71.830 82.180 72.150 82.240 ;
        RECT 73.300 82.180 73.440 82.380 ;
        RECT 91.610 82.320 91.930 82.380 ;
        RECT 92.085 82.335 92.375 82.380 ;
        RECT 94.460 82.380 96.670 82.520 ;
        RECT 108.650 82.520 108.940 82.565 ;
        RECT 110.510 82.520 110.800 82.565 ;
        RECT 108.650 82.380 110.800 82.520 ;
        RECT 69.085 82.040 73.440 82.180 ;
        RECT 73.685 82.180 73.975 82.225 ;
        RECT 93.450 82.180 93.770 82.240 ;
        RECT 94.460 82.225 94.600 82.380 ;
        RECT 108.650 82.335 108.940 82.380 ;
        RECT 110.510 82.335 110.800 82.380 ;
        RECT 111.430 82.520 111.720 82.565 ;
        RECT 113.690 82.520 114.010 82.580 ;
        RECT 114.690 82.520 114.980 82.565 ;
        RECT 111.430 82.380 114.980 82.520 ;
        RECT 111.430 82.335 111.720 82.380 ;
        RECT 113.690 82.320 114.010 82.380 ;
        RECT 114.690 82.335 114.980 82.380 ;
        RECT 73.685 82.040 93.770 82.180 ;
        RECT 69.085 81.995 69.375 82.040 ;
        RECT 71.830 81.980 72.150 82.040 ;
        RECT 73.685 81.995 73.975 82.040 ;
        RECT 93.450 81.980 93.770 82.040 ;
        RECT 94.385 81.995 94.675 82.225 ;
        RECT 97.130 81.980 97.450 82.240 ;
        RECT 5.520 81.360 118.680 81.840 ;
        RECT 12.490 80.960 12.810 81.220 ;
        RECT 13.410 80.960 13.730 81.220 ;
        RECT 15.710 80.960 16.030 81.220 ;
        RECT 60.790 80.960 61.110 81.220 ;
        RECT 64.025 80.975 64.315 81.205 ;
        RECT 64.470 81.160 64.790 81.220 ;
        RECT 69.070 81.160 69.390 81.220 ;
        RECT 85.645 81.160 85.935 81.205 ;
        RECT 64.470 81.020 69.390 81.160 ;
        RECT 64.100 80.820 64.240 80.975 ;
        RECT 64.470 80.960 64.790 81.020 ;
        RECT 69.070 80.960 69.390 81.020 ;
        RECT 75.140 81.020 85.935 81.160 ;
        RECT 65.865 80.820 66.155 80.865 ;
        RECT 64.100 80.680 66.155 80.820 ;
        RECT 65.865 80.635 66.155 80.680 ;
        RECT 68.145 80.820 68.795 80.865 ;
        RECT 71.745 80.820 72.035 80.865 ;
        RECT 74.130 80.820 74.450 80.880 ;
        RECT 68.145 80.680 74.450 80.820 ;
        RECT 68.145 80.635 68.795 80.680 ;
        RECT 71.445 80.635 72.035 80.680 ;
        RECT 12.965 80.480 13.255 80.525 ;
        RECT 13.410 80.480 13.730 80.540 ;
        RECT 12.965 80.340 13.730 80.480 ;
        RECT 12.965 80.295 13.255 80.340 ;
        RECT 13.410 80.280 13.730 80.340 ;
        RECT 15.250 80.280 15.570 80.540 ;
        RECT 60.345 80.480 60.635 80.525 ;
        RECT 62.170 80.480 62.490 80.540 ;
        RECT 60.345 80.340 62.490 80.480 ;
        RECT 60.345 80.295 60.635 80.340 ;
        RECT 62.170 80.280 62.490 80.340 ;
        RECT 63.090 80.280 63.410 80.540 ;
        RECT 64.950 80.480 65.240 80.525 ;
        RECT 66.785 80.480 67.075 80.525 ;
        RECT 70.365 80.480 70.655 80.525 ;
        RECT 64.950 80.340 70.655 80.480 ;
        RECT 64.950 80.295 65.240 80.340 ;
        RECT 66.785 80.295 67.075 80.340 ;
        RECT 70.365 80.295 70.655 80.340 ;
        RECT 71.445 80.320 71.735 80.635 ;
        RECT 74.130 80.620 74.450 80.680 ;
        RECT 75.140 80.480 75.280 81.020 ;
        RECT 85.645 80.975 85.935 81.020 ;
        RECT 98.525 81.160 98.815 81.205 ;
        RECT 103.570 81.160 103.890 81.220 ;
        RECT 98.525 81.020 103.890 81.160 ;
        RECT 98.525 80.975 98.815 81.020 ;
        RECT 103.570 80.960 103.890 81.020 ;
        RECT 80.585 80.820 80.875 80.865 ;
        RECT 83.345 80.820 83.635 80.865 ;
        RECT 80.585 80.680 83.635 80.820 ;
        RECT 80.585 80.635 80.875 80.680 ;
        RECT 83.345 80.635 83.635 80.680 ;
        RECT 93.450 80.820 93.770 80.880 ;
        RECT 96.225 80.820 96.515 80.865 ;
        RECT 93.450 80.680 96.515 80.820 ;
        RECT 93.450 80.620 93.770 80.680 ;
        RECT 96.225 80.635 96.515 80.680 ;
        RECT 72.840 80.340 75.280 80.480 ;
        RECT 76.890 80.480 77.210 80.540 ;
        RECT 77.365 80.480 77.655 80.525 ;
        RECT 76.890 80.340 77.655 80.480 ;
        RECT 16.645 80.140 16.935 80.185 ;
        RECT 19.850 80.140 20.170 80.200 ;
        RECT 16.645 80.000 20.170 80.140 ;
        RECT 16.645 79.955 16.935 80.000 ;
        RECT 19.850 79.940 20.170 80.000 ;
        RECT 64.470 79.940 64.790 80.200 ;
        RECT 72.840 80.140 72.980 80.340 ;
        RECT 76.890 80.280 77.210 80.340 ;
        RECT 77.365 80.295 77.655 80.340 ;
        RECT 78.285 80.295 78.575 80.525 ;
        RECT 78.745 80.295 79.035 80.525 ;
        RECT 65.020 80.000 72.980 80.140 ;
        RECT 73.225 80.140 73.515 80.185 ;
        RECT 76.445 80.140 76.735 80.185 ;
        RECT 78.360 80.140 78.500 80.295 ;
        RECT 73.225 80.000 78.500 80.140 ;
        RECT 78.820 80.140 78.960 80.295 ;
        RECT 79.190 80.280 79.510 80.540 ;
        RECT 84.725 80.480 85.015 80.525 ;
        RECT 87.010 80.480 87.330 80.540 ;
        RECT 84.725 80.340 87.330 80.480 ;
        RECT 84.725 80.295 85.015 80.340 ;
        RECT 87.010 80.280 87.330 80.340 ;
        RECT 97.605 80.480 97.895 80.525 ;
        RECT 98.050 80.480 98.370 80.540 ;
        RECT 97.605 80.340 98.370 80.480 ;
        RECT 97.605 80.295 97.895 80.340 ;
        RECT 98.050 80.280 98.370 80.340 ;
        RECT 79.650 80.140 79.970 80.200 ;
        RECT 78.820 80.000 79.970 80.140 ;
        RECT 64.010 79.800 64.330 79.860 ;
        RECT 65.020 79.800 65.160 80.000 ;
        RECT 73.225 79.955 73.515 80.000 ;
        RECT 76.445 79.955 76.735 80.000 ;
        RECT 79.650 79.940 79.970 80.000 ;
        RECT 84.265 80.140 84.555 80.185 ;
        RECT 86.550 80.140 86.870 80.200 ;
        RECT 84.265 80.000 86.870 80.140 ;
        RECT 84.265 79.955 84.555 80.000 ;
        RECT 86.550 79.940 86.870 80.000 ;
        RECT 97.145 80.140 97.435 80.185 ;
        RECT 98.510 80.140 98.830 80.200 ;
        RECT 97.145 80.000 98.830 80.140 ;
        RECT 97.145 79.955 97.435 80.000 ;
        RECT 98.510 79.940 98.830 80.000 ;
        RECT 64.010 79.660 65.160 79.800 ;
        RECT 65.355 79.800 65.645 79.845 ;
        RECT 67.245 79.800 67.535 79.845 ;
        RECT 70.365 79.800 70.655 79.845 ;
        RECT 87.930 79.800 88.250 79.860 ;
        RECT 65.355 79.660 70.655 79.800 ;
        RECT 64.010 79.600 64.330 79.660 ;
        RECT 65.355 79.615 65.645 79.660 ;
        RECT 67.245 79.615 67.535 79.660 ;
        RECT 70.365 79.615 70.655 79.660 ;
        RECT 84.800 79.660 88.250 79.800 ;
        RECT 21.230 79.460 21.550 79.520 ;
        RECT 23.990 79.460 24.310 79.520 ;
        RECT 21.230 79.320 24.310 79.460 ;
        RECT 21.230 79.260 21.550 79.320 ;
        RECT 23.990 79.260 24.310 79.320 ;
        RECT 73.670 79.260 73.990 79.520 ;
        RECT 84.800 79.505 84.940 79.660 ;
        RECT 87.930 79.600 88.250 79.660 ;
        RECT 84.725 79.275 85.015 79.505 ;
        RECT 97.130 79.260 97.450 79.520 ;
        RECT 5.520 78.640 118.680 79.120 ;
        RECT 22.610 78.240 22.930 78.500 ;
        RECT 23.070 78.440 23.390 78.500 ;
        RECT 24.465 78.440 24.755 78.485 ;
        RECT 23.070 78.300 24.755 78.440 ;
        RECT 23.070 78.240 23.390 78.300 ;
        RECT 24.465 78.255 24.755 78.300 ;
        RECT 52.050 78.240 52.370 78.500 ;
        RECT 63.090 78.440 63.410 78.500 ;
        RECT 65.405 78.440 65.695 78.485 ;
        RECT 63.090 78.300 65.695 78.440 ;
        RECT 63.090 78.240 63.410 78.300 ;
        RECT 65.405 78.255 65.695 78.300 ;
        RECT 74.130 78.240 74.450 78.500 ;
        RECT 103.110 78.440 103.430 78.500 ;
        RECT 103.110 78.300 112.080 78.440 ;
        RECT 103.110 78.240 103.430 78.300 ;
        RECT 13.885 77.915 14.175 78.145 ;
        RECT 22.700 78.100 22.840 78.240 ;
        RECT 21.780 77.960 22.840 78.100 ;
        RECT 23.545 78.100 23.835 78.145 ;
        RECT 23.990 78.100 24.310 78.160 ;
        RECT 23.545 77.960 24.310 78.100 ;
        RECT 13.960 77.760 14.100 77.915 ;
        RECT 11.660 77.620 14.100 77.760 ;
        RECT 15.250 77.760 15.570 77.820 ;
        RECT 16.185 77.760 16.475 77.805 ;
        RECT 15.250 77.620 16.475 77.760 ;
        RECT 11.660 77.465 11.800 77.620 ;
        RECT 15.250 77.560 15.570 77.620 ;
        RECT 16.185 77.575 16.475 77.620 ;
        RECT 17.105 77.760 17.395 77.805 ;
        RECT 19.390 77.760 19.710 77.820 ;
        RECT 17.105 77.620 19.710 77.760 ;
        RECT 17.105 77.575 17.395 77.620 ;
        RECT 11.585 77.235 11.875 77.465 ;
        RECT 13.410 77.220 13.730 77.480 ;
        RECT 16.260 77.080 16.400 77.575 ;
        RECT 19.390 77.560 19.710 77.620 ;
        RECT 19.865 77.420 20.155 77.465 ;
        RECT 20.310 77.420 20.630 77.480 ;
        RECT 19.865 77.280 20.630 77.420 ;
        RECT 19.865 77.235 20.155 77.280 ;
        RECT 20.310 77.220 20.630 77.280 ;
        RECT 20.785 77.235 21.075 77.465 ;
        RECT 20.860 77.080 21.000 77.235 ;
        RECT 21.230 77.220 21.550 77.480 ;
        RECT 21.780 77.465 21.920 77.960 ;
        RECT 23.545 77.915 23.835 77.960 ;
        RECT 23.990 77.900 24.310 77.960 ;
        RECT 44.705 77.915 44.995 78.145 ;
        RECT 51.145 78.100 51.435 78.145 ;
        RECT 57.570 78.100 57.890 78.160 ;
        RECT 51.145 77.960 57.890 78.100 ;
        RECT 51.145 77.915 51.435 77.960 ;
        RECT 22.610 77.760 22.930 77.820 ;
        RECT 24.925 77.760 25.215 77.805 ;
        RECT 22.610 77.620 25.215 77.760 ;
        RECT 22.610 77.560 22.930 77.620 ;
        RECT 24.925 77.575 25.215 77.620 ;
        RECT 21.705 77.420 21.995 77.465 ;
        RECT 23.530 77.420 23.850 77.480 ;
        RECT 21.705 77.280 23.850 77.420 ;
        RECT 21.705 77.235 21.995 77.280 ;
        RECT 23.530 77.220 23.850 77.280 ;
        RECT 23.990 77.420 24.310 77.480 ;
        RECT 24.465 77.420 24.755 77.465 ;
        RECT 23.990 77.280 24.755 77.420 ;
        RECT 23.990 77.220 24.310 77.280 ;
        RECT 24.465 77.235 24.755 77.280 ;
        RECT 36.410 77.420 36.730 77.480 ;
        RECT 38.725 77.420 39.015 77.465 ;
        RECT 36.410 77.280 39.015 77.420 ;
        RECT 36.410 77.220 36.730 77.280 ;
        RECT 38.725 77.235 39.015 77.280 ;
        RECT 42.865 77.420 43.155 77.465 ;
        RECT 44.780 77.420 44.920 77.915 ;
        RECT 57.570 77.900 57.890 77.960 ;
        RECT 62.170 78.100 62.490 78.160 ;
        RECT 64.010 78.100 64.330 78.160 ;
        RECT 62.170 77.960 64.330 78.100 ;
        RECT 62.170 77.900 62.490 77.960 ;
        RECT 64.010 77.900 64.330 77.960 ;
        RECT 69.070 78.100 69.390 78.160 ;
        RECT 81.970 78.100 82.260 78.145 ;
        RECT 83.830 78.100 84.120 78.145 ;
        RECT 86.610 78.100 86.900 78.145 ;
        RECT 69.070 77.960 81.720 78.100 ;
        RECT 69.070 77.900 69.390 77.960 ;
        RECT 47.910 77.560 48.230 77.820 ;
        RECT 63.550 77.760 63.870 77.820 ;
        RECT 68.150 77.760 68.470 77.820 ;
        RECT 77.825 77.760 78.115 77.805 ;
        RECT 78.270 77.760 78.590 77.820 ;
        RECT 81.580 77.805 81.720 77.960 ;
        RECT 81.970 77.960 86.900 78.100 ;
        RECT 81.970 77.915 82.260 77.960 ;
        RECT 83.830 77.915 84.120 77.960 ;
        RECT 86.610 77.915 86.900 77.960 ;
        RECT 101.750 78.100 102.040 78.145 ;
        RECT 103.610 78.100 103.900 78.145 ;
        RECT 106.390 78.100 106.680 78.145 ;
        RECT 101.750 77.960 106.680 78.100 ;
        RECT 101.750 77.915 102.040 77.960 ;
        RECT 103.610 77.915 103.900 77.960 ;
        RECT 106.390 77.915 106.680 77.960 ;
        RECT 63.550 77.620 78.590 77.760 ;
        RECT 63.550 77.560 63.870 77.620 ;
        RECT 68.150 77.560 68.470 77.620 ;
        RECT 77.825 77.575 78.115 77.620 ;
        RECT 78.270 77.560 78.590 77.620 ;
        RECT 81.505 77.575 81.795 77.805 ;
        RECT 82.410 77.760 82.730 77.820 ;
        RECT 90.475 77.760 90.765 77.805 ;
        RECT 82.410 77.620 90.765 77.760 ;
        RECT 82.410 77.560 82.730 77.620 ;
        RECT 42.865 77.280 44.920 77.420 ;
        RECT 46.545 77.420 46.835 77.465 ;
        RECT 48.370 77.420 48.690 77.480 ;
        RECT 46.545 77.280 48.690 77.420 ;
        RECT 42.865 77.235 43.155 77.280 ;
        RECT 46.545 77.235 46.835 77.280 ;
        RECT 48.370 77.220 48.690 77.280 ;
        RECT 51.590 77.420 51.910 77.480 ;
        RECT 52.065 77.420 52.355 77.465 ;
        RECT 51.590 77.280 52.355 77.420 ;
        RECT 51.590 77.220 51.910 77.280 ;
        RECT 52.065 77.235 52.355 77.280 ;
        RECT 52.525 77.235 52.815 77.465 ;
        RECT 16.260 76.940 21.000 77.080 ;
        RECT 23.085 77.080 23.375 77.125 ;
        RECT 25.845 77.080 26.135 77.125 ;
        RECT 23.085 76.940 26.135 77.080 ;
        RECT 23.085 76.895 23.375 76.940 ;
        RECT 25.845 76.895 26.135 76.940 ;
        RECT 9.270 76.740 9.590 76.800 ;
        RECT 10.665 76.740 10.955 76.785 ;
        RECT 9.270 76.600 10.955 76.740 ;
        RECT 9.270 76.540 9.590 76.600 ;
        RECT 10.665 76.555 10.955 76.600 ;
        RECT 12.950 76.540 13.270 76.800 ;
        RECT 15.710 76.540 16.030 76.800 ;
        RECT 35.950 76.540 36.270 76.800 ;
        RECT 41.930 76.540 42.250 76.800 ;
        RECT 46.990 76.540 47.310 76.800 ;
        RECT 52.050 76.740 52.370 76.800 ;
        RECT 52.600 76.740 52.740 77.235 ;
        RECT 67.230 77.220 67.550 77.480 ;
        RECT 74.605 77.235 74.895 77.465 ;
        RECT 78.745 77.420 79.035 77.465 ;
        RECT 82.960 77.420 83.100 77.620 ;
        RECT 90.475 77.575 90.765 77.620 ;
        RECT 96.670 77.760 96.990 77.820 ;
        RECT 101.285 77.760 101.575 77.805 ;
        RECT 96.670 77.620 101.575 77.760 ;
        RECT 96.670 77.560 96.990 77.620 ;
        RECT 101.285 77.575 101.575 77.620 ;
        RECT 103.125 77.760 103.415 77.805 ;
        RECT 104.030 77.760 104.350 77.820 ;
        RECT 103.125 77.620 104.350 77.760 ;
        RECT 103.125 77.575 103.415 77.620 ;
        RECT 104.030 77.560 104.350 77.620 ;
        RECT 78.745 77.280 83.100 77.420 ;
        RECT 78.745 77.235 79.035 77.280 ;
        RECT 53.430 76.880 53.750 77.140 ;
        RECT 67.705 77.080 67.995 77.125 ;
        RECT 73.670 77.080 73.990 77.140 ;
        RECT 67.705 76.940 73.990 77.080 ;
        RECT 74.680 77.080 74.820 77.235 ;
        RECT 83.330 77.220 83.650 77.480 ;
        RECT 86.610 77.420 86.900 77.465 ;
        RECT 84.365 77.280 86.900 77.420 ;
        RECT 77.810 77.080 78.130 77.140 ;
        RECT 84.365 77.125 84.580 77.280 ;
        RECT 86.610 77.235 86.900 77.280 ;
        RECT 92.085 77.420 92.375 77.465 ;
        RECT 102.650 77.420 102.970 77.480 ;
        RECT 111.940 77.465 112.080 78.300 ;
        RECT 106.390 77.420 106.680 77.465 ;
        RECT 92.085 77.280 102.970 77.420 ;
        RECT 92.085 77.235 92.375 77.280 ;
        RECT 82.430 77.080 82.720 77.125 ;
        RECT 84.290 77.080 84.580 77.125 ;
        RECT 74.680 76.940 82.180 77.080 ;
        RECT 67.705 76.895 67.995 76.940 ;
        RECT 73.670 76.880 73.990 76.940 ;
        RECT 77.810 76.880 78.130 76.940 ;
        RECT 82.040 76.800 82.180 76.940 ;
        RECT 82.430 76.940 84.580 77.080 ;
        RECT 82.430 76.895 82.720 76.940 ;
        RECT 84.290 76.895 84.580 76.940 ;
        RECT 85.210 77.080 85.500 77.125 ;
        RECT 88.470 77.080 88.760 77.125 ;
        RECT 91.625 77.080 91.915 77.125 ;
        RECT 85.210 76.940 91.915 77.080 ;
        RECT 85.210 76.895 85.500 76.940 ;
        RECT 88.470 76.895 88.760 76.940 ;
        RECT 91.625 76.895 91.915 76.940 ;
        RECT 52.050 76.600 52.740 76.740 ;
        RECT 52.050 76.540 52.370 76.600 ;
        RECT 79.190 76.540 79.510 76.800 ;
        RECT 81.030 76.540 81.350 76.800 ;
        RECT 81.950 76.740 82.270 76.800 ;
        RECT 92.160 76.740 92.300 77.235 ;
        RECT 102.650 77.220 102.970 77.280 ;
        RECT 104.145 77.280 106.680 77.420 ;
        RECT 104.145 77.125 104.360 77.280 ;
        RECT 106.390 77.235 106.680 77.280 ;
        RECT 111.865 77.420 112.155 77.465 ;
        RECT 113.245 77.420 113.535 77.465 ;
        RECT 111.865 77.280 113.535 77.420 ;
        RECT 111.865 77.235 112.155 77.280 ;
        RECT 113.245 77.235 113.535 77.280 ;
        RECT 102.210 77.080 102.500 77.125 ;
        RECT 104.070 77.080 104.360 77.125 ;
        RECT 102.210 76.940 104.360 77.080 ;
        RECT 102.210 76.895 102.500 76.940 ;
        RECT 104.070 76.895 104.360 76.940 ;
        RECT 104.990 77.080 105.280 77.125 ;
        RECT 108.250 77.080 108.540 77.125 ;
        RECT 111.405 77.080 111.695 77.125 ;
        RECT 104.990 76.940 111.695 77.080 ;
        RECT 104.990 76.895 105.280 76.940 ;
        RECT 108.250 76.895 108.540 76.940 ;
        RECT 111.405 76.895 111.695 76.940 ;
        RECT 81.950 76.600 92.300 76.740 ;
        RECT 110.010 76.785 110.330 76.800 ;
        RECT 81.950 76.540 82.270 76.600 ;
        RECT 110.010 76.555 110.545 76.785 ;
        RECT 110.010 76.540 110.330 76.555 ;
        RECT 112.770 76.540 113.090 76.800 ;
        RECT 5.520 75.920 118.680 76.400 ;
        RECT 15.710 75.720 16.030 75.780 ;
        RECT 18.930 75.720 19.250 75.780 ;
        RECT 19.405 75.720 19.695 75.765 ;
        RECT 15.710 75.580 19.695 75.720 ;
        RECT 15.710 75.520 16.030 75.580 ;
        RECT 18.930 75.520 19.250 75.580 ;
        RECT 19.405 75.535 19.695 75.580 ;
        RECT 23.530 75.720 23.850 75.780 ;
        RECT 24.910 75.720 25.230 75.780 ;
        RECT 35.045 75.720 35.335 75.765 ;
        RECT 35.950 75.720 36.270 75.780 ;
        RECT 23.530 75.580 25.230 75.720 ;
        RECT 23.530 75.520 23.850 75.580 ;
        RECT 24.910 75.520 25.230 75.580 ;
        RECT 25.920 75.580 36.270 75.720 ;
        RECT 8.370 75.380 8.660 75.425 ;
        RECT 10.230 75.380 10.520 75.425 ;
        RECT 8.370 75.240 10.520 75.380 ;
        RECT 8.370 75.195 8.660 75.240 ;
        RECT 10.230 75.195 10.520 75.240 ;
        RECT 11.150 75.380 11.440 75.425 ;
        RECT 12.950 75.380 13.270 75.440 ;
        RECT 14.410 75.380 14.700 75.425 ;
        RECT 11.150 75.240 14.700 75.380 ;
        RECT 11.150 75.195 11.440 75.240 ;
        RECT 6.970 75.040 7.290 75.100 ;
        RECT 7.445 75.040 7.735 75.085 ;
        RECT 6.970 74.900 7.735 75.040 ;
        RECT 6.970 74.840 7.290 74.900 ;
        RECT 7.445 74.855 7.735 74.900 ;
        RECT 9.270 74.840 9.590 75.100 ;
        RECT 10.305 75.040 10.520 75.195 ;
        RECT 12.950 75.180 13.270 75.240 ;
        RECT 14.410 75.195 14.700 75.240 ;
        RECT 15.250 75.380 15.570 75.440 ;
        RECT 16.415 75.380 16.705 75.425 ;
        RECT 25.920 75.380 26.060 75.580 ;
        RECT 35.045 75.535 35.335 75.580 ;
        RECT 35.950 75.520 36.270 75.580 ;
        RECT 46.990 75.720 47.310 75.780 ;
        RECT 47.695 75.720 47.985 75.765 ;
        RECT 50.670 75.720 50.990 75.780 ;
        RECT 46.990 75.580 50.990 75.720 ;
        RECT 46.990 75.520 47.310 75.580 ;
        RECT 47.695 75.535 47.985 75.580 ;
        RECT 50.670 75.520 50.990 75.580 ;
        RECT 53.430 75.520 53.750 75.780 ;
        RECT 54.810 75.720 55.130 75.780 ;
        RECT 59.410 75.720 59.730 75.780 ;
        RECT 54.810 75.580 59.730 75.720 ;
        RECT 54.810 75.520 55.130 75.580 ;
        RECT 59.410 75.520 59.730 75.580 ;
        RECT 61.725 75.535 62.015 75.765 ;
        RECT 69.070 75.720 69.390 75.780 ;
        RECT 69.545 75.720 69.835 75.765 ;
        RECT 69.070 75.580 69.835 75.720 ;
        RECT 15.250 75.240 16.705 75.380 ;
        RECT 15.250 75.180 15.570 75.240 ;
        RECT 16.415 75.195 16.705 75.240 ;
        RECT 19.020 75.240 26.060 75.380 ;
        RECT 26.305 75.380 26.595 75.425 ;
        RECT 26.765 75.380 27.055 75.425 ;
        RECT 39.170 75.380 39.490 75.440 ;
        RECT 42.390 75.425 42.710 75.440 ;
        RECT 26.305 75.240 27.055 75.380 ;
        RECT 19.020 75.085 19.160 75.240 ;
        RECT 26.305 75.195 26.595 75.240 ;
        RECT 26.765 75.195 27.055 75.240 ;
        RECT 34.660 75.240 39.490 75.380 ;
        RECT 12.550 75.040 12.840 75.085 ;
        RECT 10.305 74.900 12.840 75.040 ;
        RECT 12.550 74.855 12.840 74.900 ;
        RECT 18.945 74.855 19.235 75.085 ;
        RECT 20.770 75.040 21.090 75.100 ;
        RECT 23.070 75.040 23.390 75.100 ;
        RECT 20.770 74.900 23.390 75.040 ;
        RECT 20.770 74.840 21.090 74.900 ;
        RECT 23.070 74.840 23.390 74.900 ;
        RECT 24.005 74.855 24.295 75.085 ;
        RECT 24.465 74.855 24.755 75.085 ;
        RECT 19.850 74.500 20.170 74.760 ;
        RECT 7.910 74.360 8.200 74.405 ;
        RECT 9.770 74.360 10.060 74.405 ;
        RECT 12.550 74.360 12.840 74.405 ;
        RECT 7.910 74.220 12.840 74.360 ;
        RECT 24.080 74.360 24.220 74.855 ;
        RECT 24.540 74.700 24.680 74.855 ;
        RECT 24.910 74.840 25.230 75.100 ;
        RECT 27.670 75.040 27.990 75.100 ;
        RECT 34.660 75.085 34.800 75.240 ;
        RECT 39.170 75.180 39.490 75.240 ;
        RECT 39.650 75.380 39.940 75.425 ;
        RECT 41.510 75.380 41.800 75.425 ;
        RECT 39.650 75.240 41.800 75.380 ;
        RECT 39.650 75.195 39.940 75.240 ;
        RECT 41.510 75.195 41.800 75.240 ;
        RECT 28.145 75.040 28.435 75.085 ;
        RECT 27.670 74.900 28.435 75.040 ;
        RECT 27.670 74.840 27.990 74.900 ;
        RECT 28.145 74.855 28.435 74.900 ;
        RECT 30.905 75.040 31.195 75.085 ;
        RECT 30.905 74.900 32.960 75.040 ;
        RECT 30.905 74.855 31.195 74.900 ;
        RECT 25.370 74.700 25.690 74.760 ;
        RECT 24.540 74.560 25.690 74.700 ;
        RECT 25.370 74.500 25.690 74.560 ;
        RECT 27.225 74.700 27.515 74.745 ;
        RECT 29.970 74.700 30.290 74.760 ;
        RECT 27.225 74.560 30.290 74.700 ;
        RECT 27.225 74.515 27.515 74.560 ;
        RECT 29.970 74.500 30.290 74.560 ;
        RECT 32.820 74.405 32.960 74.900 ;
        RECT 34.585 74.855 34.875 75.085 ;
        RECT 37.790 74.840 38.110 75.100 ;
        RECT 38.710 74.840 39.030 75.100 ;
        RECT 41.585 75.040 41.800 75.195 ;
        RECT 42.390 75.380 42.720 75.425 ;
        RECT 45.690 75.380 45.980 75.425 ;
        RECT 42.390 75.240 45.980 75.380 ;
        RECT 42.390 75.195 42.720 75.240 ;
        RECT 45.690 75.195 45.980 75.240 ;
        RECT 50.210 75.380 50.530 75.440 ;
        RECT 61.800 75.380 61.940 75.535 ;
        RECT 69.070 75.520 69.390 75.580 ;
        RECT 69.545 75.535 69.835 75.580 ;
        RECT 71.385 75.720 71.675 75.765 ;
        RECT 73.670 75.720 73.990 75.780 ;
        RECT 71.385 75.580 73.990 75.720 ;
        RECT 71.385 75.535 71.675 75.580 ;
        RECT 73.670 75.520 73.990 75.580 ;
        RECT 81.965 75.720 82.255 75.765 ;
        RECT 83.330 75.720 83.650 75.780 ;
        RECT 81.965 75.580 83.650 75.720 ;
        RECT 81.965 75.535 82.255 75.580 ;
        RECT 83.330 75.520 83.650 75.580 ;
        RECT 91.150 75.720 91.470 75.780 ;
        RECT 93.925 75.720 94.215 75.765 ;
        RECT 94.370 75.720 94.690 75.780 ;
        RECT 96.210 75.720 96.530 75.780 ;
        RECT 103.585 75.720 103.875 75.765 ;
        RECT 91.150 75.580 92.300 75.720 ;
        RECT 91.150 75.520 91.470 75.580 ;
        RECT 71.845 75.380 72.135 75.425 ;
        RECT 74.130 75.380 74.450 75.440 ;
        RECT 81.490 75.380 81.810 75.440 ;
        RECT 85.645 75.380 85.935 75.425 ;
        RECT 50.210 75.240 62.170 75.380 ;
        RECT 42.390 75.180 42.710 75.195 ;
        RECT 50.210 75.180 50.530 75.240 ;
        RECT 43.830 75.040 44.120 75.085 ;
        RECT 41.585 74.900 44.120 75.040 ;
        RECT 43.830 74.855 44.120 74.900 ;
        RECT 49.750 74.840 50.070 75.100 ;
        RECT 50.670 74.840 50.990 75.100 ;
        RECT 51.220 75.085 51.360 75.240 ;
        RECT 51.145 74.855 51.435 75.085 ;
        RECT 51.605 75.040 51.895 75.085 ;
        RECT 52.970 75.040 53.290 75.100 ;
        RECT 54.810 75.040 55.130 75.100 ;
        RECT 55.360 75.085 55.500 75.240 ;
        RECT 51.605 74.900 55.130 75.040 ;
        RECT 51.605 74.855 51.895 74.900 ;
        RECT 52.970 74.840 53.290 74.900 ;
        RECT 54.810 74.840 55.130 74.900 ;
        RECT 55.285 74.855 55.575 75.085 ;
        RECT 55.745 74.855 56.035 75.085 ;
        RECT 56.665 74.855 56.955 75.085 ;
        RECT 60.345 74.855 60.635 75.085 ;
        RECT 35.965 74.515 36.255 74.745 ;
        RECT 40.565 74.700 40.855 74.745 ;
        RECT 41.930 74.700 42.250 74.760 ;
        RECT 40.565 74.560 42.250 74.700 ;
        RECT 40.565 74.515 40.855 74.560 ;
        RECT 24.080 74.220 32.500 74.360 ;
        RECT 7.910 74.175 8.200 74.220 ;
        RECT 9.770 74.175 10.060 74.220 ;
        RECT 12.550 74.175 12.840 74.220 ;
        RECT 17.090 73.820 17.410 74.080 ;
        RECT 26.750 73.820 27.070 74.080 ;
        RECT 28.590 74.020 28.910 74.080 ;
        RECT 29.065 74.020 29.355 74.065 ;
        RECT 28.590 73.880 29.355 74.020 ;
        RECT 28.590 73.820 28.910 73.880 ;
        RECT 29.065 73.835 29.355 73.880 ;
        RECT 29.510 74.020 29.830 74.080 ;
        RECT 29.985 74.020 30.275 74.065 ;
        RECT 29.510 73.880 30.275 74.020 ;
        RECT 32.360 74.020 32.500 74.220 ;
        RECT 32.745 74.175 33.035 74.405 ;
        RECT 36.040 74.360 36.180 74.515 ;
        RECT 41.930 74.500 42.250 74.560 ;
        RECT 46.530 74.700 46.850 74.760 ;
        RECT 55.820 74.700 55.960 74.855 ;
        RECT 46.530 74.560 55.960 74.700 ;
        RECT 46.530 74.500 46.850 74.560 ;
        RECT 39.190 74.360 39.480 74.405 ;
        RECT 41.050 74.360 41.340 74.405 ;
        RECT 43.830 74.360 44.120 74.405 ;
        RECT 36.040 74.220 38.020 74.360 ;
        RECT 36.410 74.020 36.730 74.080 ;
        RECT 32.360 73.880 36.730 74.020 ;
        RECT 29.510 73.820 29.830 73.880 ;
        RECT 29.985 73.835 30.275 73.880 ;
        RECT 36.410 73.820 36.730 73.880 ;
        RECT 37.330 73.820 37.650 74.080 ;
        RECT 37.880 74.020 38.020 74.220 ;
        RECT 39.190 74.220 44.120 74.360 ;
        RECT 39.190 74.175 39.480 74.220 ;
        RECT 41.050 74.175 41.340 74.220 ;
        RECT 43.830 74.175 44.120 74.220 ;
        RECT 49.750 74.360 50.070 74.420 ;
        RECT 54.810 74.360 55.130 74.420 ;
        RECT 56.740 74.360 56.880 74.855 ;
        RECT 60.420 74.700 60.560 74.855 ;
        RECT 60.790 74.840 61.110 75.100 ;
        RECT 62.030 75.040 62.170 75.240 ;
        RECT 71.845 75.240 77.580 75.380 ;
        RECT 71.845 75.195 72.135 75.240 ;
        RECT 74.130 75.180 74.450 75.240 ;
        RECT 67.230 75.040 67.550 75.100 ;
        RECT 76.430 75.040 76.750 75.100 ;
        RECT 77.440 75.085 77.580 75.240 ;
        RECT 81.490 75.240 85.935 75.380 ;
        RECT 81.490 75.180 81.810 75.240 ;
        RECT 85.645 75.195 85.935 75.240 ;
        RECT 89.770 75.380 90.090 75.440 ;
        RECT 89.770 75.240 91.840 75.380 ;
        RECT 89.770 75.180 90.090 75.240 ;
        RECT 62.030 74.900 67.000 75.040 ;
        RECT 62.170 74.700 62.490 74.760 ;
        RECT 60.420 74.560 62.490 74.700 ;
        RECT 62.170 74.500 62.490 74.560 ;
        RECT 49.750 74.220 56.880 74.360 ;
        RECT 66.860 74.360 67.000 74.900 ;
        RECT 67.230 74.900 76.750 75.040 ;
        RECT 67.230 74.840 67.550 74.900 ;
        RECT 76.430 74.840 76.750 74.900 ;
        RECT 77.365 74.855 77.655 75.085 ;
        RECT 77.825 74.855 78.115 75.085 ;
        RECT 68.150 74.700 68.470 74.760 ;
        RECT 72.305 74.700 72.595 74.745 ;
        RECT 77.900 74.700 78.040 74.855 ;
        RECT 78.270 74.840 78.590 75.100 ;
        RECT 81.030 74.840 81.350 75.100 ;
        RECT 84.250 74.840 84.570 75.100 ;
        RECT 88.390 75.040 88.710 75.100 ;
        RECT 91.700 75.085 91.840 75.240 ;
        RECT 92.160 75.085 92.300 75.580 ;
        RECT 93.925 75.580 94.690 75.720 ;
        RECT 93.925 75.535 94.215 75.580 ;
        RECT 94.370 75.520 94.690 75.580 ;
        RECT 95.380 75.580 96.530 75.720 ;
        RECT 93.465 75.380 93.755 75.425 ;
        RECT 95.380 75.380 95.520 75.580 ;
        RECT 96.210 75.520 96.530 75.580 ;
        RECT 103.200 75.580 103.875 75.720 ;
        RECT 101.285 75.380 101.575 75.425 ;
        RECT 93.465 75.240 95.520 75.380 ;
        RECT 96.300 75.240 101.575 75.380 ;
        RECT 93.465 75.195 93.755 75.240 ;
        RECT 96.300 75.085 96.440 75.240 ;
        RECT 101.285 75.195 101.575 75.240 ;
        RECT 90.245 75.040 90.535 75.085 ;
        RECT 88.390 74.900 90.535 75.040 ;
        RECT 88.390 74.840 88.710 74.900 ;
        RECT 90.245 74.855 90.535 74.900 ;
        RECT 91.165 74.855 91.455 75.085 ;
        RECT 91.625 74.855 91.915 75.085 ;
        RECT 92.085 75.040 92.375 75.085 ;
        RECT 95.305 75.040 95.595 75.085 ;
        RECT 92.085 74.900 95.595 75.040 ;
        RECT 92.085 74.855 92.375 74.900 ;
        RECT 95.305 74.855 95.595 74.900 ;
        RECT 95.765 74.855 96.055 75.085 ;
        RECT 96.225 74.855 96.515 75.085 ;
        RECT 79.650 74.700 79.970 74.760 ;
        RECT 68.150 74.560 72.595 74.700 ;
        RECT 68.150 74.500 68.470 74.560 ;
        RECT 72.305 74.515 72.595 74.560 ;
        RECT 75.600 74.560 79.970 74.700 ;
        RECT 75.600 74.360 75.740 74.560 ;
        RECT 79.650 74.500 79.970 74.560 ;
        RECT 80.570 74.700 80.890 74.760 ;
        RECT 84.725 74.700 85.015 74.745 ;
        RECT 80.570 74.560 85.015 74.700 ;
        RECT 80.570 74.500 80.890 74.560 ;
        RECT 84.725 74.515 85.015 74.560 ;
        RECT 66.860 74.220 75.740 74.360 ;
        RECT 75.970 74.360 76.290 74.420 ;
        RECT 83.345 74.360 83.635 74.405 ;
        RECT 75.970 74.220 83.635 74.360 ;
        RECT 49.750 74.160 50.070 74.220 ;
        RECT 54.810 74.160 55.130 74.220 ;
        RECT 75.970 74.160 76.290 74.220 ;
        RECT 83.345 74.175 83.635 74.220 ;
        RECT 47.910 74.020 48.230 74.080 ;
        RECT 37.880 73.880 48.230 74.020 ;
        RECT 47.910 73.820 48.230 73.880 ;
        RECT 52.970 73.820 53.290 74.080 ;
        RECT 59.410 74.020 59.730 74.080 ;
        RECT 78.270 74.020 78.590 74.080 ;
        RECT 59.410 73.880 78.590 74.020 ;
        RECT 59.410 73.820 59.730 73.880 ;
        RECT 78.270 73.820 78.590 73.880 ;
        RECT 79.665 74.020 79.955 74.065 ;
        RECT 82.410 74.020 82.730 74.080 ;
        RECT 79.665 73.880 82.730 74.020 ;
        RECT 79.665 73.835 79.955 73.880 ;
        RECT 82.410 73.820 82.730 73.880 ;
        RECT 83.790 74.020 84.110 74.080 ;
        RECT 84.265 74.020 84.555 74.065 ;
        RECT 83.790 73.880 84.555 74.020 ;
        RECT 90.320 74.020 90.460 74.855 ;
        RECT 91.240 74.360 91.380 74.855 ;
        RECT 91.700 74.700 91.840 74.855 ;
        RECT 95.840 74.700 95.980 74.855 ;
        RECT 97.130 74.840 97.450 75.100 ;
        RECT 98.970 74.700 99.290 74.760 ;
        RECT 100.365 74.700 100.655 74.745 ;
        RECT 91.700 74.560 95.980 74.700 ;
        RECT 96.300 74.560 98.740 74.700 ;
        RECT 96.300 74.360 96.440 74.560 ;
        RECT 91.240 74.220 96.440 74.360 ;
        RECT 98.600 74.360 98.740 74.560 ;
        RECT 98.970 74.560 100.655 74.700 ;
        RECT 101.360 74.700 101.500 75.195 ;
        RECT 101.730 74.840 102.050 75.100 ;
        RECT 103.200 75.040 103.340 75.580 ;
        RECT 103.585 75.535 103.875 75.580 ;
        RECT 104.030 75.520 104.350 75.780 ;
        RECT 104.490 75.720 104.810 75.780 ;
        RECT 110.470 75.720 110.790 75.780 ;
        RECT 111.405 75.720 111.695 75.765 ;
        RECT 104.490 75.580 111.695 75.720 ;
        RECT 104.490 75.520 104.810 75.580 ;
        RECT 110.470 75.520 110.790 75.580 ;
        RECT 111.405 75.535 111.695 75.580 ;
        RECT 110.010 75.380 110.330 75.440 ;
        RECT 110.945 75.380 111.235 75.425 ;
        RECT 106.880 75.240 111.235 75.380 ;
        RECT 104.965 75.040 105.255 75.085 ;
        RECT 103.200 74.900 105.255 75.040 ;
        RECT 104.965 74.855 105.255 74.900 ;
        RECT 106.880 74.700 107.020 75.240 ;
        RECT 110.010 75.180 110.330 75.240 ;
        RECT 110.945 75.195 111.235 75.240 ;
        RECT 107.265 75.040 107.555 75.085 ;
        RECT 107.265 74.900 109.320 75.040 ;
        RECT 107.265 74.855 107.555 74.900 ;
        RECT 101.360 74.560 107.020 74.700 ;
        RECT 98.970 74.500 99.290 74.560 ;
        RECT 100.365 74.515 100.655 74.560 ;
        RECT 104.490 74.360 104.810 74.420 ;
        RECT 109.180 74.405 109.320 74.900 ;
        RECT 111.850 74.500 112.170 74.760 ;
        RECT 98.600 74.220 104.810 74.360 ;
        RECT 104.490 74.160 104.810 74.220 ;
        RECT 109.105 74.175 109.395 74.405 ;
        RECT 97.130 74.020 97.450 74.080 ;
        RECT 90.320 73.880 97.450 74.020 ;
        RECT 83.790 73.820 84.110 73.880 ;
        RECT 84.265 73.835 84.555 73.880 ;
        RECT 97.130 73.820 97.450 73.880 ;
        RECT 108.170 73.820 108.490 74.080 ;
        RECT 5.520 73.200 118.680 73.680 ;
        RECT 18.930 72.800 19.250 73.060 ;
        RECT 36.410 72.800 36.730 73.060 ;
        RECT 42.390 73.000 42.710 73.060 ;
        RECT 42.865 73.000 43.155 73.045 ;
        RECT 42.390 72.860 43.155 73.000 ;
        RECT 42.390 72.800 42.710 72.860 ;
        RECT 42.865 72.815 43.155 72.860 ;
        RECT 51.130 73.000 51.450 73.060 ;
        RECT 52.985 73.000 53.275 73.045 ;
        RECT 51.130 72.860 53.275 73.000 ;
        RECT 51.130 72.800 51.450 72.860 ;
        RECT 52.985 72.815 53.275 72.860 ;
        RECT 55.285 73.000 55.575 73.045 ;
        RECT 57.110 73.000 57.430 73.060 ;
        RECT 55.285 72.860 57.430 73.000 ;
        RECT 55.285 72.815 55.575 72.860 ;
        RECT 57.110 72.800 57.430 72.860 ;
        RECT 61.265 73.000 61.555 73.045 ;
        RECT 63.105 73.000 63.395 73.045 ;
        RECT 67.690 73.000 68.010 73.060 ;
        RECT 61.265 72.860 62.860 73.000 ;
        RECT 61.265 72.815 61.555 72.860 ;
        RECT 9.235 72.660 9.525 72.705 ;
        RECT 11.125 72.660 11.415 72.705 ;
        RECT 14.245 72.660 14.535 72.705 ;
        RECT 9.235 72.520 14.535 72.660 ;
        RECT 9.235 72.475 9.525 72.520 ;
        RECT 11.125 72.475 11.415 72.520 ;
        RECT 14.245 72.475 14.535 72.520 ;
        RECT 21.230 72.660 21.550 72.720 ;
        RECT 28.555 72.660 28.845 72.705 ;
        RECT 30.445 72.660 30.735 72.705 ;
        RECT 33.565 72.660 33.855 72.705 ;
        RECT 21.230 72.520 24.220 72.660 ;
        RECT 21.230 72.460 21.550 72.520 ;
        RECT 6.970 72.320 7.290 72.380 ;
        RECT 8.365 72.320 8.655 72.365 ;
        RECT 6.970 72.180 8.655 72.320 ;
        RECT 6.970 72.120 7.290 72.180 ;
        RECT 8.365 72.135 8.655 72.180 ;
        RECT 17.105 72.320 17.395 72.365 ;
        RECT 21.705 72.320 21.995 72.365 ;
        RECT 24.080 72.320 24.220 72.520 ;
        RECT 28.555 72.520 33.855 72.660 ;
        RECT 28.555 72.475 28.845 72.520 ;
        RECT 30.445 72.475 30.735 72.520 ;
        RECT 33.565 72.475 33.855 72.520 ;
        RECT 38.710 72.460 39.030 72.720 ;
        RECT 39.170 72.660 39.490 72.720 ;
        RECT 54.810 72.660 55.130 72.720 ;
        RECT 62.720 72.660 62.860 72.860 ;
        RECT 63.105 72.860 68.010 73.000 ;
        RECT 63.105 72.815 63.395 72.860 ;
        RECT 67.690 72.800 68.010 72.860 ;
        RECT 81.490 72.800 81.810 73.060 ;
        RECT 84.265 73.000 84.555 73.045 ;
        RECT 88.850 73.000 89.170 73.060 ;
        RECT 84.265 72.860 89.170 73.000 ;
        RECT 84.265 72.815 84.555 72.860 ;
        RECT 88.850 72.800 89.170 72.860 ;
        RECT 91.625 73.000 91.915 73.045 ;
        RECT 92.070 73.000 92.390 73.060 ;
        RECT 91.625 72.860 92.390 73.000 ;
        RECT 91.625 72.815 91.915 72.860 ;
        RECT 92.070 72.800 92.390 72.860 ;
        RECT 68.150 72.660 68.470 72.720 ;
        RECT 39.170 72.520 46.300 72.660 ;
        RECT 39.170 72.460 39.490 72.520 ;
        RECT 25.370 72.320 25.690 72.380 ;
        RECT 17.105 72.180 23.760 72.320 ;
        RECT 17.105 72.135 17.395 72.180 ;
        RECT 21.705 72.135 21.995 72.180 ;
        RECT 8.830 71.980 9.120 72.025 ;
        RECT 10.665 71.980 10.955 72.025 ;
        RECT 14.245 71.980 14.535 72.025 ;
        RECT 8.830 71.840 14.535 71.980 ;
        RECT 8.830 71.795 9.120 71.840 ;
        RECT 10.665 71.795 10.955 71.840 ;
        RECT 14.245 71.795 14.535 71.840 ;
        RECT 9.730 71.440 10.050 71.700 ;
        RECT 12.025 71.640 12.675 71.685 ;
        RECT 14.790 71.640 15.110 71.700 ;
        RECT 15.325 71.685 15.615 72.000 ;
        RECT 22.625 71.980 22.915 72.025 ;
        RECT 23.070 71.980 23.390 72.040 ;
        RECT 23.620 72.025 23.760 72.180 ;
        RECT 24.080 72.180 25.690 72.320 ;
        RECT 24.080 72.025 24.220 72.180 ;
        RECT 25.370 72.120 25.690 72.180 ;
        RECT 27.685 72.320 27.975 72.365 ;
        RECT 38.800 72.320 38.940 72.460 ;
        RECT 27.685 72.180 38.940 72.320 ;
        RECT 40.640 72.180 42.620 72.320 ;
        RECT 27.685 72.135 27.975 72.180 ;
        RECT 22.625 71.840 23.390 71.980 ;
        RECT 22.625 71.795 22.915 71.840 ;
        RECT 23.070 71.780 23.390 71.840 ;
        RECT 23.545 71.795 23.835 72.025 ;
        RECT 24.005 71.795 24.295 72.025 ;
        RECT 24.465 71.980 24.755 72.025 ;
        RECT 24.910 71.980 25.230 72.040 ;
        RECT 24.465 71.840 25.230 71.980 ;
        RECT 24.465 71.795 24.755 71.840 ;
        RECT 24.910 71.780 25.230 71.840 ;
        RECT 28.150 71.980 28.440 72.025 ;
        RECT 29.985 71.980 30.275 72.025 ;
        RECT 33.565 71.980 33.855 72.025 ;
        RECT 28.150 71.840 33.855 71.980 ;
        RECT 28.150 71.795 28.440 71.840 ;
        RECT 29.985 71.795 30.275 71.840 ;
        RECT 33.565 71.795 33.855 71.840 ;
        RECT 15.325 71.640 15.915 71.685 ;
        RECT 12.025 71.500 15.915 71.640 ;
        RECT 12.025 71.455 12.675 71.500 ;
        RECT 14.790 71.440 15.110 71.500 ;
        RECT 15.625 71.455 15.915 71.500 ;
        RECT 16.170 71.640 16.490 71.700 ;
        RECT 29.065 71.640 29.355 71.685 ;
        RECT 29.510 71.640 29.830 71.700 ;
        RECT 34.645 71.685 34.935 72.000 ;
        RECT 38.725 71.980 39.015 72.025 ;
        RECT 40.640 71.980 40.780 72.180 ;
        RECT 42.480 72.025 42.620 72.180 ;
        RECT 38.725 71.840 40.780 71.980 ;
        RECT 38.725 71.795 39.015 71.840 ;
        RECT 16.170 71.500 28.820 71.640 ;
        RECT 16.170 71.440 16.490 71.500 ;
        RECT 25.845 71.300 26.135 71.345 ;
        RECT 28.130 71.300 28.450 71.360 ;
        RECT 25.845 71.160 28.450 71.300 ;
        RECT 28.680 71.300 28.820 71.500 ;
        RECT 29.065 71.500 29.830 71.640 ;
        RECT 29.065 71.455 29.355 71.500 ;
        RECT 29.510 71.440 29.830 71.500 ;
        RECT 31.345 71.640 31.995 71.685 ;
        RECT 34.645 71.640 35.235 71.685 ;
        RECT 37.330 71.640 37.650 71.700 ;
        RECT 31.345 71.500 37.650 71.640 ;
        RECT 31.345 71.455 31.995 71.500 ;
        RECT 34.945 71.455 35.235 71.500 ;
        RECT 37.330 71.440 37.650 71.500 ;
        RECT 38.800 71.300 38.940 71.795 ;
        RECT 41.025 71.675 41.315 71.905 ;
        RECT 42.405 71.795 42.695 72.025 ;
        RECT 28.680 71.160 38.940 71.300 ;
        RECT 25.845 71.115 26.135 71.160 ;
        RECT 28.130 71.100 28.450 71.160 ;
        RECT 39.170 71.100 39.490 71.360 ;
        RECT 39.630 71.300 39.950 71.360 ;
        RECT 40.105 71.300 40.395 71.345 ;
        RECT 39.630 71.160 40.395 71.300 ;
        RECT 41.100 71.300 41.240 71.675 ;
        RECT 44.705 71.300 44.995 71.345 ;
        RECT 41.100 71.160 44.995 71.300 ;
        RECT 46.160 71.300 46.300 72.520 ;
        RECT 54.810 72.520 62.400 72.660 ;
        RECT 62.720 72.520 68.470 72.660 ;
        RECT 54.810 72.460 55.130 72.520 ;
        RECT 47.910 72.120 48.230 72.380 ;
        RECT 53.430 72.120 53.750 72.380 ;
        RECT 46.545 71.980 46.835 72.025 ;
        RECT 46.990 71.980 47.310 72.040 ;
        RECT 46.545 71.840 47.310 71.980 ;
        RECT 46.545 71.795 46.835 71.840 ;
        RECT 46.990 71.780 47.310 71.840 ;
        RECT 48.000 71.640 48.140 72.120 ;
        RECT 52.970 71.780 53.290 72.040 ;
        RECT 54.365 71.980 54.655 72.025 ;
        RECT 57.110 71.980 57.430 72.040 ;
        RECT 54.365 71.840 57.430 71.980 ;
        RECT 54.365 71.795 54.655 71.840 ;
        RECT 57.110 71.780 57.430 71.840 ;
        RECT 55.745 71.640 56.035 71.685 ;
        RECT 48.000 71.500 56.035 71.640 ;
        RECT 55.745 71.455 56.035 71.500 ;
        RECT 57.585 71.640 57.875 71.685 ;
        RECT 58.030 71.640 58.350 71.700 ;
        RECT 59.885 71.640 60.175 71.685 ;
        RECT 57.585 71.500 60.175 71.640 ;
        RECT 57.585 71.455 57.875 71.500 ;
        RECT 58.030 71.440 58.350 71.500 ;
        RECT 59.885 71.455 60.175 71.500 ;
        RECT 46.530 71.300 46.850 71.360 ;
        RECT 47.005 71.300 47.295 71.345 ;
        RECT 46.160 71.160 47.295 71.300 ;
        RECT 61.800 71.300 61.940 72.520 ;
        RECT 62.260 72.320 62.400 72.520 ;
        RECT 68.150 72.460 68.470 72.520 ;
        RECT 72.750 72.660 73.070 72.720 ;
        RECT 81.965 72.660 82.255 72.705 ;
        RECT 72.750 72.520 82.255 72.660 ;
        RECT 72.750 72.460 73.070 72.520 ;
        RECT 81.965 72.475 82.255 72.520 ;
        RECT 107.730 72.660 108.020 72.705 ;
        RECT 109.590 72.660 109.880 72.705 ;
        RECT 112.370 72.660 112.660 72.705 ;
        RECT 107.730 72.520 112.660 72.660 ;
        RECT 107.730 72.475 108.020 72.520 ;
        RECT 109.590 72.475 109.880 72.520 ;
        RECT 112.370 72.475 112.660 72.520 ;
        RECT 67.230 72.320 67.550 72.380 ;
        RECT 62.260 72.180 67.550 72.320 ;
        RECT 68.240 72.320 68.380 72.460 ;
        RECT 75.065 72.320 75.355 72.365 ;
        RECT 68.240 72.180 75.355 72.320 ;
        RECT 67.230 72.120 67.550 72.180 ;
        RECT 75.065 72.135 75.355 72.180 ;
        RECT 78.730 72.320 79.050 72.380 ;
        RECT 82.410 72.320 82.730 72.380 ;
        RECT 96.670 72.320 96.990 72.380 ;
        RECT 107.265 72.320 107.555 72.365 ;
        RECT 78.730 72.180 80.340 72.320 ;
        RECT 78.730 72.120 79.050 72.180 ;
        RECT 62.170 71.780 62.490 72.040 ;
        RECT 63.550 71.980 63.870 72.040 ;
        RECT 65.405 71.980 65.695 72.025 ;
        RECT 63.550 71.840 65.695 71.980 ;
        RECT 63.550 71.780 63.870 71.840 ;
        RECT 65.405 71.795 65.695 71.840 ;
        RECT 69.070 71.780 69.390 72.040 ;
        RECT 70.465 71.980 70.755 72.025 ;
        RECT 70.465 71.840 72.520 71.980 ;
        RECT 70.465 71.795 70.755 71.840 ;
        RECT 64.485 71.300 64.775 71.345 ;
        RECT 61.800 71.160 64.775 71.300 ;
        RECT 39.630 71.100 39.950 71.160 ;
        RECT 40.105 71.115 40.395 71.160 ;
        RECT 44.705 71.115 44.995 71.160 ;
        RECT 46.530 71.100 46.850 71.160 ;
        RECT 47.005 71.115 47.295 71.160 ;
        RECT 64.485 71.115 64.775 71.160 ;
        RECT 67.230 71.300 67.550 71.360 ;
        RECT 68.165 71.300 68.455 71.345 ;
        RECT 67.230 71.160 68.455 71.300 ;
        RECT 67.230 71.100 67.550 71.160 ;
        RECT 68.165 71.115 68.455 71.160 ;
        RECT 71.385 71.300 71.675 71.345 ;
        RECT 71.830 71.300 72.150 71.360 ;
        RECT 72.380 71.345 72.520 71.840 ;
        RECT 74.130 71.780 74.450 72.040 ;
        RECT 76.430 71.980 76.750 72.040 ;
        RECT 78.285 71.980 78.575 72.025 ;
        RECT 76.430 71.840 78.575 71.980 ;
        RECT 76.430 71.780 76.750 71.840 ;
        RECT 78.285 71.795 78.575 71.840 ;
        RECT 79.190 71.780 79.510 72.040 ;
        RECT 79.650 71.780 79.970 72.040 ;
        RECT 80.200 72.025 80.340 72.180 ;
        RECT 82.410 72.180 84.480 72.320 ;
        RECT 82.410 72.120 82.730 72.180 ;
        RECT 80.125 71.795 80.415 72.025 ;
        RECT 82.870 71.780 83.190 72.040 ;
        RECT 83.330 71.780 83.650 72.040 ;
        RECT 84.340 72.025 84.480 72.180 ;
        RECT 96.670 72.180 107.555 72.320 ;
        RECT 96.670 72.120 96.990 72.180 ;
        RECT 107.265 72.135 107.555 72.180 ;
        RECT 108.170 72.320 108.490 72.380 ;
        RECT 109.105 72.320 109.395 72.365 ;
        RECT 108.170 72.180 109.395 72.320 ;
        RECT 108.170 72.120 108.490 72.180 ;
        RECT 109.105 72.135 109.395 72.180 ;
        RECT 110.470 72.320 110.790 72.380 ;
        RECT 116.235 72.320 116.525 72.365 ;
        RECT 110.470 72.180 116.525 72.320 ;
        RECT 110.470 72.120 110.790 72.180 ;
        RECT 116.235 72.135 116.525 72.180 ;
        RECT 84.265 71.795 84.555 72.025 ;
        RECT 87.930 71.980 88.250 72.040 ;
        RECT 88.405 71.980 88.695 72.025 ;
        RECT 87.930 71.840 88.695 71.980 ;
        RECT 87.930 71.780 88.250 71.840 ;
        RECT 88.405 71.795 88.695 71.840 ;
        RECT 89.325 71.795 89.615 72.025 ;
        RECT 74.605 71.640 74.895 71.685 ;
        RECT 79.280 71.640 79.420 71.780 ;
        RECT 74.605 71.500 79.420 71.640 ;
        RECT 89.400 71.640 89.540 71.795 ;
        RECT 89.770 71.780 90.090 72.040 ;
        RECT 90.245 71.980 90.535 72.025 ;
        RECT 91.150 71.980 91.470 72.040 ;
        RECT 90.245 71.840 91.470 71.980 ;
        RECT 90.245 71.795 90.535 71.840 ;
        RECT 91.150 71.780 91.470 71.840 ;
        RECT 97.130 71.780 97.450 72.040 ;
        RECT 99.905 71.980 100.195 72.025 ;
        RECT 103.110 71.980 103.430 72.040 ;
        RECT 112.370 71.980 112.660 72.025 ;
        RECT 99.905 71.840 103.430 71.980 ;
        RECT 99.905 71.795 100.195 71.840 ;
        RECT 103.110 71.780 103.430 71.840 ;
        RECT 110.125 71.840 112.660 71.980 ;
        RECT 101.730 71.640 102.050 71.700 ;
        RECT 110.125 71.685 110.340 71.840 ;
        RECT 112.370 71.795 112.660 71.840 ;
        RECT 89.400 71.500 102.050 71.640 ;
        RECT 74.605 71.455 74.895 71.500 ;
        RECT 101.730 71.440 102.050 71.500 ;
        RECT 108.190 71.640 108.480 71.685 ;
        RECT 110.050 71.640 110.340 71.685 ;
        RECT 108.190 71.500 110.340 71.640 ;
        RECT 108.190 71.455 108.480 71.500 ;
        RECT 110.050 71.455 110.340 71.500 ;
        RECT 110.970 71.640 111.260 71.685 ;
        RECT 112.770 71.640 113.090 71.700 ;
        RECT 114.230 71.640 114.520 71.685 ;
        RECT 110.970 71.500 114.520 71.640 ;
        RECT 110.970 71.455 111.260 71.500 ;
        RECT 112.770 71.440 113.090 71.500 ;
        RECT 114.230 71.455 114.520 71.500 ;
        RECT 71.385 71.160 72.150 71.300 ;
        RECT 71.385 71.115 71.675 71.160 ;
        RECT 71.830 71.100 72.150 71.160 ;
        RECT 72.305 71.115 72.595 71.345 ;
        RECT 95.750 71.300 96.070 71.360 ;
        RECT 96.225 71.300 96.515 71.345 ;
        RECT 95.750 71.160 96.515 71.300 ;
        RECT 95.750 71.100 96.070 71.160 ;
        RECT 96.225 71.115 96.515 71.160 ;
        RECT 99.430 71.100 99.750 71.360 ;
        RECT 5.520 70.480 118.680 70.960 ;
        RECT 9.730 70.280 10.050 70.340 ;
        RECT 11.585 70.280 11.875 70.325 ;
        RECT 9.730 70.140 11.875 70.280 ;
        RECT 9.730 70.080 10.050 70.140 ;
        RECT 11.585 70.095 11.875 70.140 ;
        RECT 13.885 70.280 14.175 70.325 ;
        RECT 14.790 70.280 15.110 70.340 ;
        RECT 20.770 70.280 21.090 70.340 ;
        RECT 24.450 70.280 24.770 70.340 ;
        RECT 13.885 70.140 15.110 70.280 ;
        RECT 13.885 70.095 14.175 70.140 ;
        RECT 14.790 70.080 15.110 70.140 ;
        RECT 20.400 70.140 21.090 70.280 ;
        RECT 17.090 69.940 17.410 70.000 ;
        RECT 12.580 69.800 17.410 69.940 ;
        RECT 12.580 69.645 12.720 69.800 ;
        RECT 17.090 69.740 17.410 69.800 ;
        RECT 12.505 69.415 12.795 69.645 ;
        RECT 13.410 69.600 13.730 69.660 ;
        RECT 20.400 69.600 20.540 70.140 ;
        RECT 20.770 70.080 21.090 70.140 ;
        RECT 21.320 70.140 24.770 70.280 ;
        RECT 13.410 69.460 20.540 69.600 ;
        RECT 20.785 69.600 21.075 69.645 ;
        RECT 21.320 69.600 21.460 70.140 ;
        RECT 24.450 70.080 24.770 70.140 ;
        RECT 27.670 70.080 27.990 70.340 ;
        RECT 30.445 70.280 30.735 70.325 ;
        RECT 31.350 70.280 31.670 70.340 ;
        RECT 30.445 70.140 31.670 70.280 ;
        RECT 30.445 70.095 30.735 70.140 ;
        RECT 31.350 70.080 31.670 70.140 ;
        RECT 39.170 70.280 39.490 70.340 ;
        RECT 46.530 70.325 46.850 70.340 ;
        RECT 39.170 70.140 40.780 70.280 ;
        RECT 39.170 70.080 39.490 70.140 ;
        RECT 24.005 69.940 24.295 69.985 ;
        RECT 24.005 69.800 26.980 69.940 ;
        RECT 24.005 69.755 24.295 69.800 ;
        RECT 20.785 69.460 21.460 69.600 ;
        RECT 13.410 69.400 13.730 69.460 ;
        RECT 20.785 69.415 21.075 69.460 ;
        RECT 21.705 69.415 21.995 69.645 ;
        RECT 22.165 69.415 22.455 69.645 ;
        RECT 22.625 69.600 22.915 69.645 ;
        RECT 23.530 69.600 23.850 69.660 ;
        RECT 22.625 69.460 23.850 69.600 ;
        RECT 22.625 69.415 22.915 69.460 ;
        RECT 16.630 69.260 16.950 69.320 ;
        RECT 21.780 69.260 21.920 69.415 ;
        RECT 16.630 69.120 21.920 69.260 ;
        RECT 22.240 69.260 22.380 69.415 ;
        RECT 23.530 69.400 23.850 69.460 ;
        RECT 24.450 69.400 24.770 69.660 ;
        RECT 25.370 69.400 25.690 69.660 ;
        RECT 25.845 69.415 26.135 69.645 ;
        RECT 23.070 69.260 23.390 69.320 ;
        RECT 22.240 69.120 23.390 69.260 ;
        RECT 16.630 69.060 16.950 69.120 ;
        RECT 23.070 69.060 23.390 69.120 ;
        RECT 25.920 69.260 26.060 69.415 ;
        RECT 26.290 69.400 26.610 69.660 ;
        RECT 26.840 69.600 26.980 69.800 ;
        RECT 28.130 69.740 28.450 70.000 ;
        RECT 38.270 69.940 38.560 69.985 ;
        RECT 40.130 69.940 40.420 69.985 ;
        RECT 38.270 69.800 40.420 69.940 ;
        RECT 40.640 69.940 40.780 70.140 ;
        RECT 46.315 70.095 46.850 70.325 ;
        RECT 46.530 70.080 46.850 70.095 ;
        RECT 58.030 70.080 58.350 70.340 ;
        RECT 62.630 70.280 62.950 70.340 ;
        RECT 58.580 70.140 62.950 70.280 ;
        RECT 41.050 69.940 41.340 69.985 ;
        RECT 44.310 69.940 44.600 69.985 ;
        RECT 40.640 69.800 44.600 69.940 ;
        RECT 38.270 69.755 38.560 69.800 ;
        RECT 40.130 69.755 40.420 69.800 ;
        RECT 41.050 69.755 41.340 69.800 ;
        RECT 44.310 69.755 44.600 69.800 ;
        RECT 45.150 69.940 45.470 70.000 ;
        RECT 58.580 69.940 58.720 70.140 ;
        RECT 62.630 70.080 62.950 70.140 ;
        RECT 74.130 70.325 74.450 70.340 ;
        RECT 74.130 70.095 74.665 70.325 ;
        RECT 82.410 70.280 82.730 70.340 ;
        RECT 91.150 70.280 91.470 70.340 ;
        RECT 93.465 70.280 93.755 70.325 ;
        RECT 98.050 70.280 98.370 70.340 ;
        RECT 82.410 70.140 92.300 70.280 ;
        RECT 74.130 70.080 74.450 70.095 ;
        RECT 82.410 70.080 82.730 70.140 ;
        RECT 91.150 70.080 91.470 70.140 ;
        RECT 45.150 69.800 58.720 69.940 ;
        RECT 59.410 69.940 59.730 70.000 ;
        RECT 60.790 69.940 61.110 70.000 ;
        RECT 66.330 69.940 66.620 69.985 ;
        RECT 68.190 69.940 68.480 69.985 ;
        RECT 59.410 69.800 61.940 69.940 ;
        RECT 29.525 69.600 29.815 69.645 ;
        RECT 26.840 69.460 29.815 69.600 ;
        RECT 29.525 69.415 29.815 69.460 ;
        RECT 37.345 69.600 37.635 69.645 ;
        RECT 40.205 69.600 40.420 69.755 ;
        RECT 45.150 69.740 45.470 69.800 ;
        RECT 59.410 69.740 59.730 69.800 ;
        RECT 60.790 69.740 61.110 69.800 ;
        RECT 42.450 69.600 42.740 69.645 ;
        RECT 37.345 69.460 39.860 69.600 ;
        RECT 40.205 69.460 42.740 69.600 ;
        RECT 37.345 69.415 37.635 69.460 ;
        RECT 25.920 69.120 27.900 69.260 ;
        RECT 18.470 68.920 18.790 68.980 ;
        RECT 24.910 68.920 25.230 68.980 ;
        RECT 18.470 68.780 25.230 68.920 ;
        RECT 18.470 68.720 18.790 68.780 ;
        RECT 24.910 68.720 25.230 68.780 ;
        RECT 23.070 68.580 23.390 68.640 ;
        RECT 25.920 68.580 26.060 69.120 ;
        RECT 27.760 68.980 27.900 69.120 ;
        RECT 28.590 69.060 28.910 69.320 ;
        RECT 39.170 69.060 39.490 69.320 ;
        RECT 39.720 69.260 39.860 69.460 ;
        RECT 42.450 69.415 42.740 69.460 ;
        RECT 58.045 69.600 58.335 69.645 ;
        RECT 59.885 69.600 60.175 69.645 ;
        RECT 61.250 69.600 61.570 69.660 ;
        RECT 61.800 69.645 61.940 69.800 ;
        RECT 66.330 69.800 68.480 69.940 ;
        RECT 66.330 69.755 66.620 69.800 ;
        RECT 68.190 69.755 68.480 69.800 ;
        RECT 69.110 69.940 69.400 69.985 ;
        RECT 72.370 69.940 72.660 69.985 ;
        RECT 75.525 69.940 75.815 69.985 ;
        RECT 69.110 69.800 75.815 69.940 ;
        RECT 69.110 69.755 69.400 69.800 ;
        RECT 72.370 69.755 72.660 69.800 ;
        RECT 75.525 69.755 75.815 69.800 ;
        RECT 89.770 69.940 90.090 70.000 ;
        RECT 89.770 69.800 91.840 69.940 ;
        RECT 58.045 69.460 59.640 69.600 ;
        RECT 58.045 69.415 58.335 69.460 ;
        RECT 41.010 69.260 41.330 69.320 ;
        RECT 39.720 69.120 41.330 69.260 ;
        RECT 41.010 69.060 41.330 69.120 ;
        RECT 58.505 69.260 58.795 69.305 ;
        RECT 58.950 69.260 59.270 69.320 ;
        RECT 58.505 69.120 59.270 69.260 ;
        RECT 59.500 69.260 59.640 69.460 ;
        RECT 59.885 69.460 61.570 69.600 ;
        RECT 59.885 69.415 60.175 69.460 ;
        RECT 61.250 69.400 61.570 69.460 ;
        RECT 61.725 69.415 62.015 69.645 ;
        RECT 62.170 69.600 62.490 69.660 ;
        RECT 64.470 69.600 64.790 69.660 ;
        RECT 65.405 69.600 65.695 69.645 ;
        RECT 62.170 69.460 64.240 69.600 ;
        RECT 62.170 69.400 62.490 69.460 ;
        RECT 63.550 69.260 63.870 69.320 ;
        RECT 59.500 69.120 63.870 69.260 ;
        RECT 64.100 69.260 64.240 69.460 ;
        RECT 64.470 69.460 65.695 69.600 ;
        RECT 64.470 69.400 64.790 69.460 ;
        RECT 65.405 69.415 65.695 69.460 ;
        RECT 67.230 69.400 67.550 69.660 ;
        RECT 68.265 69.600 68.480 69.755 ;
        RECT 89.770 69.740 90.090 69.800 ;
        RECT 70.510 69.600 70.800 69.645 ;
        RECT 68.265 69.460 70.800 69.600 ;
        RECT 70.510 69.415 70.800 69.460 ;
        RECT 75.970 69.600 76.290 69.660 ;
        RECT 81.950 69.600 82.270 69.660 ;
        RECT 75.970 69.460 82.270 69.600 ;
        RECT 75.970 69.400 76.290 69.460 ;
        RECT 81.950 69.400 82.270 69.460 ;
        RECT 88.390 69.600 88.710 69.660 ;
        RECT 90.245 69.600 90.535 69.645 ;
        RECT 88.390 69.460 90.535 69.600 ;
        RECT 88.390 69.400 88.710 69.460 ;
        RECT 90.245 69.415 90.535 69.460 ;
        RECT 68.610 69.260 68.930 69.320 ;
        RECT 64.100 69.120 68.930 69.260 ;
        RECT 58.505 69.075 58.795 69.120 ;
        RECT 58.950 69.060 59.270 69.120 ;
        RECT 63.550 69.060 63.870 69.120 ;
        RECT 68.610 69.060 68.930 69.120 ;
        RECT 27.670 68.920 27.990 68.980 ;
        RECT 37.810 68.920 38.100 68.965 ;
        RECT 39.670 68.920 39.960 68.965 ;
        RECT 42.450 68.920 42.740 68.965 ;
        RECT 63.090 68.920 63.410 68.980 ;
        RECT 27.670 68.780 34.340 68.920 ;
        RECT 27.670 68.720 27.990 68.780 ;
        RECT 34.200 68.640 34.340 68.780 ;
        RECT 37.810 68.780 42.740 68.920 ;
        RECT 37.810 68.735 38.100 68.780 ;
        RECT 39.670 68.735 39.960 68.780 ;
        RECT 42.450 68.735 42.740 68.780 ;
        RECT 48.230 68.780 63.410 68.920 ;
        RECT 23.070 68.440 26.060 68.580 ;
        RECT 29.525 68.580 29.815 68.625 ;
        RECT 29.970 68.580 30.290 68.640 ;
        RECT 29.525 68.440 30.290 68.580 ;
        RECT 23.070 68.380 23.390 68.440 ;
        RECT 29.525 68.395 29.815 68.440 ;
        RECT 29.970 68.380 30.290 68.440 ;
        RECT 34.110 68.580 34.430 68.640 ;
        RECT 48.230 68.580 48.370 68.780 ;
        RECT 63.090 68.720 63.410 68.780 ;
        RECT 65.870 68.920 66.160 68.965 ;
        RECT 67.730 68.920 68.020 68.965 ;
        RECT 70.510 68.920 70.800 68.965 ;
        RECT 65.870 68.780 70.800 68.920 ;
        RECT 65.870 68.735 66.160 68.780 ;
        RECT 67.730 68.735 68.020 68.780 ;
        RECT 70.510 68.735 70.800 68.780 ;
        RECT 78.730 68.920 79.050 68.980 ;
        RECT 90.780 68.920 90.920 69.800 ;
        RECT 91.700 69.645 91.840 69.800 ;
        RECT 92.160 69.645 92.300 70.140 ;
        RECT 93.465 70.140 98.370 70.280 ;
        RECT 93.465 70.095 93.755 70.140 ;
        RECT 98.050 70.080 98.370 70.140 ;
        RECT 101.730 70.280 102.050 70.340 ;
        RECT 102.895 70.280 103.185 70.325 ;
        RECT 101.730 70.140 103.185 70.280 ;
        RECT 101.730 70.080 102.050 70.140 ;
        RECT 102.895 70.095 103.185 70.140 ;
        RECT 110.470 70.280 110.790 70.340 ;
        RECT 110.945 70.280 111.235 70.325 ;
        RECT 110.470 70.140 111.235 70.280 ;
        RECT 110.470 70.080 110.790 70.140 ;
        RECT 110.945 70.095 111.235 70.140 ;
        RECT 94.850 69.940 95.140 69.985 ;
        RECT 96.710 69.940 97.000 69.985 ;
        RECT 94.850 69.800 97.000 69.940 ;
        RECT 94.850 69.755 95.140 69.800 ;
        RECT 96.710 69.755 97.000 69.800 ;
        RECT 97.630 69.940 97.920 69.985 ;
        RECT 99.430 69.940 99.750 70.000 ;
        RECT 100.890 69.940 101.180 69.985 ;
        RECT 97.630 69.800 101.180 69.940 ;
        RECT 97.630 69.755 97.920 69.800 ;
        RECT 91.165 69.415 91.455 69.645 ;
        RECT 91.625 69.415 91.915 69.645 ;
        RECT 92.085 69.415 92.375 69.645 ;
        RECT 93.925 69.600 94.215 69.645 ;
        RECT 96.210 69.600 96.530 69.660 ;
        RECT 93.925 69.460 96.530 69.600 ;
        RECT 96.785 69.600 97.000 69.755 ;
        RECT 99.430 69.740 99.750 69.800 ;
        RECT 100.890 69.755 101.180 69.800 ;
        RECT 99.030 69.600 99.320 69.645 ;
        RECT 96.785 69.460 99.320 69.600 ;
        RECT 93.925 69.415 94.215 69.460 ;
        RECT 91.240 69.260 91.380 69.415 ;
        RECT 96.210 69.400 96.530 69.460 ;
        RECT 99.030 69.415 99.320 69.460 ;
        RECT 95.290 69.260 95.610 69.320 ;
        RECT 91.240 69.120 95.610 69.260 ;
        RECT 95.290 69.060 95.610 69.120 ;
        RECT 95.750 69.060 96.070 69.320 ;
        RECT 110.930 69.260 111.250 69.320 ;
        RECT 111.405 69.260 111.695 69.305 ;
        RECT 110.930 69.120 111.695 69.260 ;
        RECT 110.930 69.060 111.250 69.120 ;
        RECT 111.405 69.075 111.695 69.120 ;
        RECT 111.850 69.060 112.170 69.320 ;
        RECT 78.730 68.780 90.920 68.920 ;
        RECT 94.390 68.920 94.680 68.965 ;
        RECT 96.250 68.920 96.540 68.965 ;
        RECT 99.030 68.920 99.320 68.965 ;
        RECT 94.390 68.780 99.320 68.920 ;
        RECT 78.730 68.720 79.050 68.780 ;
        RECT 94.390 68.735 94.680 68.780 ;
        RECT 96.250 68.735 96.540 68.780 ;
        RECT 99.030 68.735 99.320 68.780 ;
        RECT 34.110 68.440 48.370 68.580 ;
        RECT 34.110 68.380 34.430 68.440 ;
        RECT 59.410 68.380 59.730 68.640 ;
        RECT 60.805 68.580 61.095 68.625 ;
        RECT 62.630 68.580 62.950 68.640 ;
        RECT 60.805 68.440 62.950 68.580 ;
        RECT 60.805 68.395 61.095 68.440 ;
        RECT 62.630 68.380 62.950 68.440 ;
        RECT 105.410 68.580 105.730 68.640 ;
        RECT 109.105 68.580 109.395 68.625 ;
        RECT 105.410 68.440 109.395 68.580 ;
        RECT 105.410 68.380 105.730 68.440 ;
        RECT 109.105 68.395 109.395 68.440 ;
        RECT 5.520 67.760 118.680 68.240 ;
        RECT 22.150 67.560 22.470 67.620 ;
        RECT 22.625 67.560 22.915 67.605 ;
        RECT 26.290 67.560 26.610 67.620 ;
        RECT 29.050 67.560 29.370 67.620 ;
        RECT 29.525 67.560 29.815 67.605 ;
        RECT 22.150 67.420 22.915 67.560 ;
        RECT 22.150 67.360 22.470 67.420 ;
        RECT 22.625 67.375 22.915 67.420 ;
        RECT 24.540 67.420 28.360 67.560 ;
        RECT 24.540 67.220 24.680 67.420 ;
        RECT 26.290 67.360 26.610 67.420 ;
        RECT 24.080 67.080 24.680 67.220 ;
        RECT 15.250 66.680 15.570 66.940 ;
        RECT 16.645 66.540 16.935 66.585 ;
        RECT 19.850 66.540 20.170 66.600 ;
        RECT 16.645 66.400 20.170 66.540 ;
        RECT 16.645 66.355 16.935 66.400 ;
        RECT 19.850 66.340 20.170 66.400 ;
        RECT 23.530 66.540 23.850 66.600 ;
        RECT 24.080 66.585 24.220 67.080 ;
        RECT 24.540 66.740 27.900 66.880 ;
        RECT 24.540 66.585 24.680 66.740 ;
        RECT 27.760 66.600 27.900 66.740 ;
        RECT 24.005 66.540 24.295 66.585 ;
        RECT 23.530 66.400 24.295 66.540 ;
        RECT 23.530 66.340 23.850 66.400 ;
        RECT 24.005 66.355 24.295 66.400 ;
        RECT 24.465 66.355 24.755 66.585 ;
        RECT 24.925 66.355 25.215 66.585 ;
        RECT 25.845 66.540 26.135 66.585 ;
        RECT 26.305 66.540 26.595 66.585 ;
        RECT 27.225 66.540 27.515 66.585 ;
        RECT 25.845 66.400 26.595 66.540 ;
        RECT 25.845 66.355 26.135 66.400 ;
        RECT 26.305 66.355 26.595 66.400 ;
        RECT 26.840 66.400 27.515 66.540 ;
        RECT 22.150 66.200 22.470 66.260 ;
        RECT 25.000 66.200 25.140 66.355 ;
        RECT 22.150 66.060 25.140 66.200 ;
        RECT 22.150 66.000 22.470 66.060 ;
        RECT 21.230 65.860 21.550 65.920 ;
        RECT 24.450 65.860 24.770 65.920 ;
        RECT 26.380 65.860 26.520 66.355 ;
        RECT 26.840 66.200 26.980 66.400 ;
        RECT 27.225 66.355 27.515 66.400 ;
        RECT 27.670 66.340 27.990 66.600 ;
        RECT 28.220 66.585 28.360 67.420 ;
        RECT 29.050 67.420 29.815 67.560 ;
        RECT 29.050 67.360 29.370 67.420 ;
        RECT 29.525 67.375 29.815 67.420 ;
        RECT 32.285 67.560 32.575 67.605 ;
        RECT 33.190 67.560 33.510 67.620 ;
        RECT 32.285 67.420 33.510 67.560 ;
        RECT 32.285 67.375 32.575 67.420 ;
        RECT 33.190 67.360 33.510 67.420 ;
        RECT 52.510 67.360 52.830 67.620 ;
        RECT 56.205 67.560 56.495 67.605 ;
        RECT 56.650 67.560 56.970 67.620 ;
        RECT 56.205 67.420 56.970 67.560 ;
        RECT 56.205 67.375 56.495 67.420 ;
        RECT 56.650 67.360 56.970 67.420 ;
        RECT 63.090 67.560 63.410 67.620 ;
        RECT 78.730 67.560 79.050 67.620 ;
        RECT 63.090 67.420 79.050 67.560 ;
        RECT 63.090 67.360 63.410 67.420 ;
        RECT 78.730 67.360 79.050 67.420 ;
        RECT 79.190 67.605 79.510 67.620 ;
        RECT 79.190 67.375 79.725 67.605 ;
        RECT 83.790 67.560 84.110 67.620 ;
        RECT 85.645 67.560 85.935 67.605 ;
        RECT 87.930 67.560 88.250 67.620 ;
        RECT 83.790 67.420 85.935 67.560 ;
        RECT 79.190 67.360 79.510 67.375 ;
        RECT 83.790 67.360 84.110 67.420 ;
        RECT 85.645 67.375 85.935 67.420 ;
        RECT 86.180 67.420 88.250 67.560 ;
        RECT 86.180 67.280 86.320 67.420 ;
        RECT 87.930 67.360 88.250 67.420 ;
        RECT 89.310 67.360 89.630 67.620 ;
        RECT 92.990 67.360 93.310 67.620 ;
        RECT 96.225 67.560 96.515 67.605 ;
        RECT 97.130 67.560 97.450 67.620 ;
        RECT 96.225 67.420 97.450 67.560 ;
        RECT 96.225 67.375 96.515 67.420 ;
        RECT 97.130 67.360 97.450 67.420 ;
        RECT 30.430 67.220 30.750 67.280 ;
        RECT 50.670 67.220 50.990 67.280 ;
        RECT 54.350 67.220 54.670 67.280 ;
        RECT 30.430 67.080 35.720 67.220 ;
        RECT 30.430 67.020 30.750 67.080 ;
        RECT 33.740 66.740 35.260 66.880 ;
        RECT 33.740 66.585 33.880 66.740 ;
        RECT 28.145 66.540 28.435 66.585 ;
        RECT 33.665 66.540 33.955 66.585 ;
        RECT 28.145 66.400 33.955 66.540 ;
        RECT 28.145 66.355 28.435 66.400 ;
        RECT 33.665 66.355 33.955 66.400 ;
        RECT 34.110 66.340 34.430 66.600 ;
        RECT 34.570 66.340 34.890 66.600 ;
        RECT 29.970 66.200 30.290 66.260 ;
        RECT 26.840 66.060 30.290 66.200 ;
        RECT 35.120 66.200 35.260 66.740 ;
        RECT 35.580 66.585 35.720 67.080 ;
        RECT 50.670 67.080 54.670 67.220 ;
        RECT 50.670 67.020 50.990 67.080 ;
        RECT 54.350 67.020 54.670 67.080 ;
        RECT 70.930 67.220 71.220 67.265 ;
        RECT 72.790 67.220 73.080 67.265 ;
        RECT 75.570 67.220 75.860 67.265 ;
        RECT 86.090 67.220 86.410 67.280 ;
        RECT 100.810 67.220 101.130 67.280 ;
        RECT 70.930 67.080 75.860 67.220 ;
        RECT 70.930 67.035 71.220 67.080 ;
        RECT 72.790 67.035 73.080 67.080 ;
        RECT 75.570 67.035 75.860 67.080 ;
        RECT 82.500 67.080 86.410 67.220 ;
        RECT 56.650 66.880 56.970 66.940 ;
        RECT 49.380 66.740 56.970 66.880 ;
        RECT 35.505 66.540 35.795 66.585 ;
        RECT 48.370 66.540 48.690 66.600 ;
        RECT 49.380 66.585 49.520 66.740 ;
        RECT 35.505 66.400 48.690 66.540 ;
        RECT 35.505 66.355 35.795 66.400 ;
        RECT 48.370 66.340 48.690 66.400 ;
        RECT 49.305 66.355 49.595 66.585 ;
        RECT 50.210 66.340 50.530 66.600 ;
        RECT 50.670 66.340 50.990 66.600 ;
        RECT 51.130 66.340 51.450 66.600 ;
        RECT 53.060 66.585 53.200 66.740 ;
        RECT 56.650 66.680 56.970 66.740 ;
        RECT 67.230 66.680 67.550 66.940 ;
        RECT 71.830 66.880 72.150 66.940 ;
        RECT 72.305 66.880 72.595 66.925 ;
        RECT 71.830 66.740 72.595 66.880 ;
        RECT 71.830 66.680 72.150 66.740 ;
        RECT 72.305 66.695 72.595 66.740 ;
        RECT 52.985 66.355 53.275 66.585 ;
        RECT 53.905 66.540 54.195 66.585 ;
        RECT 53.520 66.400 54.195 66.540 ;
        RECT 52.050 66.200 52.370 66.260 ;
        RECT 53.520 66.200 53.660 66.400 ;
        RECT 53.905 66.355 54.195 66.400 ;
        RECT 54.350 66.340 54.670 66.600 ;
        RECT 54.810 66.340 55.130 66.600 ;
        RECT 58.490 66.340 58.810 66.600 ;
        RECT 69.070 66.540 69.390 66.600 ;
        RECT 70.465 66.540 70.755 66.585 ;
        RECT 75.570 66.540 75.860 66.585 ;
        RECT 69.070 66.400 70.755 66.540 ;
        RECT 69.070 66.340 69.390 66.400 ;
        RECT 70.465 66.355 70.755 66.400 ;
        RECT 73.325 66.400 75.860 66.540 ;
        RECT 35.120 66.060 48.370 66.200 ;
        RECT 29.970 66.000 30.290 66.060 ;
        RECT 30.430 65.860 30.750 65.920 ;
        RECT 21.230 65.720 30.750 65.860 ;
        RECT 48.230 65.860 48.370 66.060 ;
        RECT 52.050 66.060 53.660 66.200 ;
        RECT 54.900 66.200 55.040 66.340 ;
        RECT 58.950 66.200 59.270 66.260 ;
        RECT 73.325 66.245 73.540 66.400 ;
        RECT 75.570 66.355 75.860 66.400 ;
        RECT 79.190 66.540 79.510 66.600 ;
        RECT 82.500 66.585 82.640 67.080 ;
        RECT 86.090 67.020 86.410 67.080 ;
        RECT 87.100 67.080 101.130 67.220 ;
        RECT 82.960 66.740 84.020 66.880 ;
        RECT 82.425 66.540 82.715 66.585 ;
        RECT 79.190 66.400 82.715 66.540 ;
        RECT 79.190 66.340 79.510 66.400 ;
        RECT 82.425 66.355 82.715 66.400 ;
        RECT 54.900 66.060 59.270 66.200 ;
        RECT 52.050 66.000 52.370 66.060 ;
        RECT 58.950 66.000 59.270 66.060 ;
        RECT 71.390 66.200 71.680 66.245 ;
        RECT 73.250 66.200 73.540 66.245 ;
        RECT 71.390 66.060 73.540 66.200 ;
        RECT 71.390 66.015 71.680 66.060 ;
        RECT 73.250 66.015 73.540 66.060 ;
        RECT 74.130 66.245 74.450 66.260 ;
        RECT 74.130 66.200 74.460 66.245 ;
        RECT 77.430 66.200 77.720 66.245 ;
        RECT 74.130 66.060 77.720 66.200 ;
        RECT 74.130 66.015 74.460 66.060 ;
        RECT 77.430 66.015 77.720 66.060 ;
        RECT 79.650 66.200 79.970 66.260 ;
        RECT 82.960 66.200 83.100 66.740 ;
        RECT 83.880 66.585 84.020 66.740 ;
        RECT 83.345 66.355 83.635 66.585 ;
        RECT 83.805 66.355 84.095 66.585 ;
        RECT 84.265 66.355 84.555 66.585 ;
        RECT 79.650 66.060 83.100 66.200 ;
        RECT 74.130 66.000 74.450 66.015 ;
        RECT 79.650 66.000 79.970 66.060 ;
        RECT 65.850 65.860 66.170 65.920 ;
        RECT 82.410 65.860 82.730 65.920 ;
        RECT 48.230 65.720 82.730 65.860 ;
        RECT 83.420 65.860 83.560 66.355 ;
        RECT 84.340 66.200 84.480 66.355 ;
        RECT 86.090 66.340 86.410 66.600 ;
        RECT 87.100 66.585 87.240 67.080 ;
        RECT 100.810 67.020 101.130 67.080 ;
        RECT 106.345 67.035 106.635 67.265 ;
        RECT 107.270 67.220 107.560 67.265 ;
        RECT 109.130 67.220 109.420 67.265 ;
        RECT 111.910 67.220 112.200 67.265 ;
        RECT 107.270 67.080 112.200 67.220 ;
        RECT 107.270 67.035 107.560 67.080 ;
        RECT 109.130 67.035 109.420 67.080 ;
        RECT 111.910 67.035 112.200 67.080 ;
        RECT 89.310 66.880 89.630 66.940 ;
        RECT 98.970 66.880 99.290 66.940 ;
        RECT 102.190 66.880 102.510 66.940 ;
        RECT 87.560 66.740 89.630 66.880 ;
        RECT 87.560 66.585 87.700 66.740 ;
        RECT 89.310 66.680 89.630 66.740 ;
        RECT 90.780 66.740 98.740 66.880 ;
        RECT 90.780 66.585 90.920 66.740 ;
        RECT 87.000 66.355 87.290 66.585 ;
        RECT 87.500 66.355 87.790 66.585 ;
        RECT 87.945 66.355 88.235 66.585 ;
        RECT 89.785 66.355 90.075 66.585 ;
        RECT 90.705 66.355 90.995 66.585 ;
        RECT 88.020 66.200 88.160 66.355 ;
        RECT 84.340 66.060 88.160 66.200 ;
        RECT 89.860 66.200 90.000 66.355 ;
        RECT 91.150 66.340 91.470 66.600 ;
        RECT 91.625 66.540 91.915 66.585 ;
        RECT 91.625 66.400 92.760 66.540 ;
        RECT 91.625 66.355 91.915 66.400 ;
        RECT 92.070 66.200 92.390 66.260 ;
        RECT 89.860 66.060 92.390 66.200 ;
        RECT 88.020 65.920 88.160 66.060 ;
        RECT 92.070 66.000 92.390 66.060 ;
        RECT 83.790 65.860 84.110 65.920 ;
        RECT 83.420 65.720 84.110 65.860 ;
        RECT 21.230 65.660 21.550 65.720 ;
        RECT 24.450 65.660 24.770 65.720 ;
        RECT 30.430 65.660 30.750 65.720 ;
        RECT 65.850 65.660 66.170 65.720 ;
        RECT 82.410 65.660 82.730 65.720 ;
        RECT 83.790 65.660 84.110 65.720 ;
        RECT 87.930 65.860 88.250 65.920 ;
        RECT 91.150 65.860 91.470 65.920 ;
        RECT 92.620 65.860 92.760 66.400 ;
        RECT 98.600 66.200 98.740 66.740 ;
        RECT 98.970 66.740 102.510 66.880 ;
        RECT 106.420 66.880 106.560 67.035 ;
        RECT 108.645 66.880 108.935 66.925 ;
        RECT 106.420 66.740 108.935 66.880 ;
        RECT 98.970 66.680 99.290 66.740 ;
        RECT 102.190 66.680 102.510 66.740 ;
        RECT 108.645 66.695 108.935 66.740 ;
        RECT 99.430 66.540 99.750 66.600 ;
        RECT 101.730 66.540 102.050 66.600 ;
        RECT 99.430 66.400 102.050 66.540 ;
        RECT 99.430 66.340 99.750 66.400 ;
        RECT 101.730 66.340 102.050 66.400 ;
        RECT 105.410 66.340 105.730 66.600 ;
        RECT 105.870 66.540 106.190 66.600 ;
        RECT 106.805 66.540 107.095 66.585 ;
        RECT 111.910 66.540 112.200 66.585 ;
        RECT 105.870 66.400 107.095 66.540 ;
        RECT 105.870 66.340 106.190 66.400 ;
        RECT 106.805 66.355 107.095 66.400 ;
        RECT 109.665 66.400 112.200 66.540 ;
        RECT 109.665 66.245 109.880 66.400 ;
        RECT 111.910 66.355 112.200 66.400 ;
        RECT 113.690 66.245 114.010 66.260 ;
        RECT 107.730 66.200 108.020 66.245 ;
        RECT 109.590 66.200 109.880 66.245 ;
        RECT 98.600 66.060 100.580 66.200 ;
        RECT 87.930 65.720 92.760 65.860 ;
        RECT 87.930 65.660 88.250 65.720 ;
        RECT 91.150 65.660 91.470 65.720 ;
        RECT 98.050 65.660 98.370 65.920 ;
        RECT 98.525 65.860 98.815 65.905 ;
        RECT 99.430 65.860 99.750 65.920 ;
        RECT 98.525 65.720 99.750 65.860 ;
        RECT 100.440 65.860 100.580 66.060 ;
        RECT 107.730 66.060 109.880 66.200 ;
        RECT 107.730 66.015 108.020 66.060 ;
        RECT 109.590 66.015 109.880 66.060 ;
        RECT 110.510 66.200 110.800 66.245 ;
        RECT 113.690 66.200 114.060 66.245 ;
        RECT 110.510 66.060 114.060 66.200 ;
        RECT 110.510 66.015 110.800 66.060 ;
        RECT 113.690 66.015 114.060 66.060 ;
        RECT 113.690 66.000 114.010 66.015 ;
        RECT 110.930 65.860 111.250 65.920 ;
        RECT 115.775 65.860 116.065 65.905 ;
        RECT 100.440 65.720 116.065 65.860 ;
        RECT 98.525 65.675 98.815 65.720 ;
        RECT 99.430 65.660 99.750 65.720 ;
        RECT 110.930 65.660 111.250 65.720 ;
        RECT 115.775 65.675 116.065 65.720 ;
        RECT 5.520 65.040 118.680 65.520 ;
        RECT 23.990 64.840 24.310 64.900 ;
        RECT 24.925 64.840 25.215 64.885 ;
        RECT 23.990 64.700 25.215 64.840 ;
        RECT 23.990 64.640 24.310 64.700 ;
        RECT 24.925 64.655 25.215 64.700 ;
        RECT 57.110 64.840 57.430 64.900 ;
        RECT 57.585 64.840 57.875 64.885 ;
        RECT 57.110 64.700 57.875 64.840 ;
        RECT 57.110 64.640 57.430 64.700 ;
        RECT 57.585 64.655 57.875 64.700 ;
        RECT 58.950 64.840 59.270 64.900 ;
        RECT 72.305 64.840 72.595 64.885 ;
        RECT 74.130 64.840 74.450 64.900 ;
        RECT 58.950 64.700 72.060 64.840 ;
        RECT 58.950 64.640 59.270 64.700 ;
        RECT 20.770 64.500 21.090 64.560 ;
        RECT 37.790 64.500 38.110 64.560 ;
        RECT 49.750 64.545 50.070 64.560 ;
        RECT 43.790 64.500 44.080 64.545 ;
        RECT 45.650 64.500 45.940 64.545 ;
        RECT 20.770 64.360 40.320 64.500 ;
        RECT 20.770 64.300 21.090 64.360 ;
        RECT 21.230 64.160 21.550 64.220 ;
        RECT 21.705 64.160 21.995 64.205 ;
        RECT 21.230 64.020 21.995 64.160 ;
        RECT 21.230 63.960 21.550 64.020 ;
        RECT 21.705 63.975 21.995 64.020 ;
        RECT 22.625 63.975 22.915 64.205 ;
        RECT 16.170 63.620 16.490 63.880 ;
        RECT 12.030 63.140 12.350 63.200 ;
        RECT 13.425 63.140 13.715 63.185 ;
        RECT 12.030 63.000 13.715 63.140 ;
        RECT 12.030 62.940 12.350 63.000 ;
        RECT 13.425 62.955 13.715 63.000 ;
        RECT 20.770 63.140 21.090 63.200 ;
        RECT 22.700 63.140 22.840 63.975 ;
        RECT 23.070 63.960 23.390 64.220 ;
        RECT 23.530 63.960 23.850 64.220 ;
        RECT 23.990 64.160 24.310 64.220 ;
        RECT 27.225 64.160 27.515 64.205 ;
        RECT 23.990 64.020 27.515 64.160 ;
        RECT 23.990 63.960 24.310 64.020 ;
        RECT 27.225 63.975 27.515 64.020 ;
        RECT 27.670 63.960 27.990 64.220 ;
        RECT 33.280 64.205 33.420 64.360 ;
        RECT 37.790 64.300 38.110 64.360 ;
        RECT 33.205 63.975 33.495 64.205 ;
        RECT 36.410 63.960 36.730 64.220 ;
        RECT 40.180 64.205 40.320 64.360 ;
        RECT 43.790 64.360 45.940 64.500 ;
        RECT 43.790 64.315 44.080 64.360 ;
        RECT 45.650 64.315 45.940 64.360 ;
        RECT 46.570 64.500 46.860 64.545 ;
        RECT 49.750 64.500 50.120 64.545 ;
        RECT 46.570 64.360 50.120 64.500 ;
        RECT 46.570 64.315 46.860 64.360 ;
        RECT 49.750 64.315 50.120 64.360 ;
        RECT 50.670 64.500 50.990 64.560 ;
        RECT 56.650 64.500 56.970 64.560 ;
        RECT 71.920 64.500 72.060 64.700 ;
        RECT 72.305 64.700 74.450 64.840 ;
        RECT 72.305 64.655 72.595 64.700 ;
        RECT 74.130 64.640 74.450 64.700 ;
        RECT 79.650 64.840 79.970 64.900 ;
        RECT 82.425 64.840 82.715 64.885 ;
        RECT 82.870 64.840 83.190 64.900 ;
        RECT 79.650 64.700 80.800 64.840 ;
        RECT 79.650 64.640 79.970 64.700 ;
        RECT 80.660 64.500 80.800 64.700 ;
        RECT 82.425 64.700 83.190 64.840 ;
        RECT 82.425 64.655 82.715 64.700 ;
        RECT 82.870 64.640 83.190 64.700 ;
        RECT 87.010 64.640 87.330 64.900 ;
        RECT 89.770 64.640 90.090 64.900 ;
        RECT 90.690 64.640 91.010 64.900 ;
        RECT 98.050 64.640 98.370 64.900 ;
        RECT 109.105 64.655 109.395 64.885 ;
        RECT 89.860 64.500 90.000 64.640 ;
        RECT 96.670 64.500 96.990 64.560 ;
        RECT 50.670 64.360 55.040 64.500 ;
        RECT 40.105 63.975 40.395 64.205 ;
        RECT 41.930 64.160 42.250 64.220 ;
        RECT 42.865 64.160 43.155 64.205 ;
        RECT 41.930 64.020 43.155 64.160 ;
        RECT 45.725 64.160 45.940 64.315 ;
        RECT 49.750 64.300 50.070 64.315 ;
        RECT 50.670 64.300 50.990 64.360 ;
        RECT 47.970 64.160 48.260 64.205 ;
        RECT 45.725 64.020 48.260 64.160 ;
        RECT 40.180 63.820 40.320 63.975 ;
        RECT 41.930 63.960 42.250 64.020 ;
        RECT 42.865 63.975 43.155 64.020 ;
        RECT 47.970 63.975 48.260 64.020 ;
        RECT 51.130 64.160 51.450 64.220 ;
        RECT 53.890 64.160 54.210 64.220 ;
        RECT 54.900 64.205 55.040 64.360 ;
        RECT 56.650 64.360 61.020 64.500 ;
        RECT 71.920 64.360 79.880 64.500 ;
        RECT 56.650 64.300 56.970 64.360 ;
        RECT 54.365 64.160 54.655 64.205 ;
        RECT 51.130 64.020 54.655 64.160 ;
        RECT 51.130 63.960 51.450 64.020 ;
        RECT 53.890 63.960 54.210 64.020 ;
        RECT 54.365 63.975 54.655 64.020 ;
        RECT 54.825 63.975 55.115 64.205 ;
        RECT 55.285 63.975 55.575 64.205 ;
        RECT 56.205 64.160 56.495 64.205 ;
        RECT 56.740 64.160 56.880 64.300 ;
        RECT 56.205 64.020 56.880 64.160 ;
        RECT 56.205 63.975 56.495 64.020 ;
        RECT 44.230 63.820 44.550 63.880 ;
        RECT 40.180 63.680 44.550 63.820 ;
        RECT 44.230 63.620 44.550 63.680 ;
        RECT 44.690 63.620 45.010 63.880 ;
        RECT 23.530 63.480 23.850 63.540 ;
        RECT 26.305 63.480 26.595 63.525 ;
        RECT 23.530 63.340 26.595 63.480 ;
        RECT 23.530 63.280 23.850 63.340 ;
        RECT 26.305 63.295 26.595 63.340 ;
        RECT 43.330 63.480 43.620 63.525 ;
        RECT 45.190 63.480 45.480 63.525 ;
        RECT 47.970 63.480 48.260 63.525 ;
        RECT 43.330 63.340 48.260 63.480 ;
        RECT 54.900 63.480 55.040 63.975 ;
        RECT 55.360 63.820 55.500 63.975 ;
        RECT 58.950 63.960 59.270 64.220 ;
        RECT 59.425 63.975 59.715 64.205 ;
        RECT 56.650 63.820 56.970 63.880 ;
        RECT 55.360 63.680 56.970 63.820 ;
        RECT 56.650 63.620 56.970 63.680 ;
        RECT 59.500 63.480 59.640 63.975 ;
        RECT 59.870 63.960 60.190 64.220 ;
        RECT 60.880 64.205 61.020 64.360 ;
        RECT 60.805 63.975 61.095 64.205 ;
        RECT 62.630 64.160 62.950 64.220 ;
        RECT 63.550 64.160 63.870 64.220 ;
        RECT 64.485 64.160 64.775 64.205 ;
        RECT 62.630 64.020 64.775 64.160 ;
        RECT 60.880 63.820 61.020 63.975 ;
        RECT 62.630 63.960 62.950 64.020 ;
        RECT 63.550 63.960 63.870 64.020 ;
        RECT 64.485 63.975 64.775 64.020 ;
        RECT 69.085 64.160 69.375 64.205 ;
        RECT 69.990 64.160 70.310 64.220 ;
        RECT 69.085 64.020 70.310 64.160 ;
        RECT 69.085 63.975 69.375 64.020 ;
        RECT 69.990 63.960 70.310 64.020 ;
        RECT 70.465 64.160 70.755 64.205 ;
        RECT 71.845 64.160 72.135 64.205 ;
        RECT 75.970 64.160 76.290 64.220 ;
        RECT 70.465 64.020 76.290 64.160 ;
        RECT 70.465 63.975 70.755 64.020 ;
        RECT 71.845 63.975 72.135 64.020 ;
        RECT 75.970 63.960 76.290 64.020 ;
        RECT 79.190 63.960 79.510 64.220 ;
        RECT 79.280 63.820 79.420 63.960 ;
        RECT 60.880 63.680 79.420 63.820 ;
        RECT 79.740 63.820 79.880 64.360 ;
        RECT 80.660 64.360 92.760 64.500 ;
        RECT 80.110 63.960 80.430 64.220 ;
        RECT 80.660 64.205 80.800 64.360 ;
        RECT 80.585 63.975 80.875 64.205 ;
        RECT 81.045 64.160 81.335 64.205 ;
        RECT 87.930 64.160 88.250 64.220 ;
        RECT 88.940 64.205 89.080 64.360 ;
        RECT 88.405 64.160 88.695 64.205 ;
        RECT 81.045 64.020 88.695 64.160 ;
        RECT 81.045 63.975 81.335 64.020 ;
        RECT 81.120 63.820 81.260 63.975 ;
        RECT 87.930 63.960 88.250 64.020 ;
        RECT 88.405 63.975 88.695 64.020 ;
        RECT 88.865 63.975 89.155 64.205 ;
        RECT 89.325 64.160 89.615 64.205 ;
        RECT 89.770 64.160 90.090 64.220 ;
        RECT 89.325 64.020 90.090 64.160 ;
        RECT 89.325 63.975 89.615 64.020 ;
        RECT 89.770 63.960 90.090 64.020 ;
        RECT 90.305 64.160 90.595 64.205 ;
        RECT 91.150 64.160 91.470 64.220 ;
        RECT 92.620 64.205 92.760 64.360 ;
        RECT 93.080 64.360 104.720 64.500 ;
        RECT 93.080 64.205 93.220 64.360 ;
        RECT 96.670 64.300 96.990 64.360 ;
        RECT 92.085 64.160 92.375 64.205 ;
        RECT 90.305 63.975 90.690 64.160 ;
        RECT 79.740 63.680 81.260 63.820 ;
        RECT 82.410 63.820 82.730 63.880 ;
        RECT 86.105 63.820 86.395 63.865 ;
        RECT 82.410 63.680 86.395 63.820 ;
        RECT 62.170 63.480 62.490 63.540 ;
        RECT 63.640 63.525 63.780 63.680 ;
        RECT 54.900 63.340 62.490 63.480 ;
        RECT 43.330 63.295 43.620 63.340 ;
        RECT 45.190 63.295 45.480 63.340 ;
        RECT 47.970 63.295 48.260 63.340 ;
        RECT 62.170 63.280 62.490 63.340 ;
        RECT 63.565 63.295 63.855 63.525 ;
        RECT 79.280 63.480 79.420 63.680 ;
        RECT 82.410 63.620 82.730 63.680 ;
        RECT 86.105 63.635 86.395 63.680 ;
        RECT 90.550 63.820 90.690 63.975 ;
        RECT 91.150 64.020 92.375 64.160 ;
        RECT 91.150 63.960 91.470 64.020 ;
        RECT 92.085 63.975 92.375 64.020 ;
        RECT 92.545 63.975 92.835 64.205 ;
        RECT 93.005 63.975 93.295 64.205 ;
        RECT 93.925 63.975 94.215 64.205 ;
        RECT 97.130 64.160 97.450 64.220 ;
        RECT 100.810 64.160 101.130 64.220 ;
        RECT 104.580 64.205 104.720 64.360 ;
        RECT 97.130 64.020 101.130 64.160 ;
        RECT 94.000 63.820 94.140 63.975 ;
        RECT 97.130 63.960 97.450 64.020 ;
        RECT 100.810 63.960 101.130 64.020 ;
        RECT 104.505 63.975 104.795 64.205 ;
        RECT 108.185 64.160 108.475 64.205 ;
        RECT 109.180 64.160 109.320 64.655 ;
        RECT 110.930 64.640 111.250 64.900 ;
        RECT 113.690 64.640 114.010 64.900 ;
        RECT 114.165 64.160 114.455 64.205 ;
        RECT 114.625 64.160 114.915 64.205 ;
        RECT 108.185 64.020 109.320 64.160 ;
        RECT 110.330 64.020 114.915 64.160 ;
        RECT 108.185 63.975 108.475 64.020 ;
        RECT 90.550 63.680 94.140 63.820 ;
        RECT 103.110 63.820 103.430 63.880 ;
        RECT 110.330 63.820 110.470 64.020 ;
        RECT 114.165 63.975 114.455 64.020 ;
        RECT 114.625 63.975 114.915 64.020 ;
        RECT 103.110 63.680 110.470 63.820 ;
        RECT 90.550 63.480 90.690 63.680 ;
        RECT 103.110 63.620 103.430 63.680 ;
        RECT 111.390 63.620 111.710 63.880 ;
        RECT 111.850 63.620 112.170 63.880 ;
        RECT 79.280 63.340 90.690 63.480 ;
        RECT 102.190 63.480 102.510 63.540 ;
        RECT 111.940 63.480 112.080 63.620 ;
        RECT 102.190 63.340 112.080 63.480 ;
        RECT 102.190 63.280 102.510 63.340 ;
        RECT 20.770 63.000 22.840 63.140 ;
        RECT 28.130 63.140 28.450 63.200 ;
        RECT 28.605 63.140 28.895 63.185 ;
        RECT 28.130 63.000 28.895 63.140 ;
        RECT 20.770 62.940 21.090 63.000 ;
        RECT 28.130 62.940 28.450 63.000 ;
        RECT 28.605 62.955 28.895 63.000 ;
        RECT 32.730 62.940 33.050 63.200 ;
        RECT 35.505 63.140 35.795 63.185 ;
        RECT 35.950 63.140 36.270 63.200 ;
        RECT 35.505 63.000 36.270 63.140 ;
        RECT 35.505 62.955 35.795 63.000 ;
        RECT 35.950 62.940 36.270 63.000 ;
        RECT 38.710 63.140 39.030 63.200 ;
        RECT 52.050 63.185 52.370 63.200 ;
        RECT 39.645 63.140 39.935 63.185 ;
        RECT 38.710 63.000 39.935 63.140 ;
        RECT 38.710 62.940 39.030 63.000 ;
        RECT 39.645 62.955 39.935 63.000 ;
        RECT 51.835 62.955 52.370 63.185 ;
        RECT 52.050 62.940 52.370 62.955 ;
        RECT 52.970 62.940 53.290 63.200 ;
        RECT 61.250 63.140 61.570 63.200 ;
        RECT 61.725 63.140 62.015 63.185 ;
        RECT 61.250 63.000 62.015 63.140 ;
        RECT 61.250 62.940 61.570 63.000 ;
        RECT 61.725 62.955 62.015 63.000 ;
        RECT 80.110 63.140 80.430 63.200 ;
        RECT 82.410 63.140 82.730 63.200 ;
        RECT 80.110 63.000 82.730 63.140 ;
        RECT 80.110 62.940 80.430 63.000 ;
        RECT 82.410 62.940 82.730 63.000 ;
        RECT 83.330 62.940 83.650 63.200 ;
        RECT 101.730 62.940 102.050 63.200 ;
        RECT 107.250 62.940 107.570 63.200 ;
        RECT 114.150 63.140 114.470 63.200 ;
        RECT 115.085 63.140 115.375 63.185 ;
        RECT 114.150 63.000 115.375 63.140 ;
        RECT 114.150 62.940 114.470 63.000 ;
        RECT 115.085 62.955 115.375 63.000 ;
        RECT 5.520 62.320 118.680 62.800 ;
        RECT 14.345 62.120 14.635 62.165 ;
        RECT 16.170 62.120 16.490 62.180 ;
        RECT 14.345 61.980 16.490 62.120 ;
        RECT 14.345 61.935 14.635 61.980 ;
        RECT 16.170 61.920 16.490 61.980 ;
        RECT 22.150 62.120 22.470 62.180 ;
        RECT 44.690 62.120 45.010 62.180 ;
        RECT 45.625 62.120 45.915 62.165 ;
        RECT 49.750 62.120 50.070 62.180 ;
        RECT 51.605 62.120 51.895 62.165 ;
        RECT 22.150 61.980 22.840 62.120 ;
        RECT 22.150 61.920 22.470 61.980 ;
        RECT 17.565 61.440 17.855 61.485 ;
        RECT 20.310 61.440 20.630 61.500 ;
        RECT 21.705 61.440 21.995 61.485 ;
        RECT 17.565 61.300 21.995 61.440 ;
        RECT 17.565 61.255 17.855 61.300 ;
        RECT 20.310 61.240 20.630 61.300 ;
        RECT 21.705 61.255 21.995 61.300 ;
        RECT 22.700 61.160 22.840 61.980 ;
        RECT 44.690 61.980 45.915 62.120 ;
        RECT 44.690 61.920 45.010 61.980 ;
        RECT 45.625 61.935 45.915 61.980 ;
        RECT 46.620 61.980 47.680 62.120 ;
        RECT 34.590 61.780 34.880 61.825 ;
        RECT 36.450 61.780 36.740 61.825 ;
        RECT 39.230 61.780 39.520 61.825 ;
        RECT 34.590 61.640 39.520 61.780 ;
        RECT 34.590 61.595 34.880 61.640 ;
        RECT 36.450 61.595 36.740 61.640 ;
        RECT 39.230 61.595 39.520 61.640 ;
        RECT 44.230 61.780 44.550 61.840 ;
        RECT 46.620 61.780 46.760 61.980 ;
        RECT 44.230 61.640 46.760 61.780 ;
        RECT 44.230 61.580 44.550 61.640 ;
        RECT 47.005 61.595 47.295 61.825 ;
        RECT 27.210 61.440 27.530 61.500 ;
        RECT 27.210 61.300 31.120 61.440 ;
        RECT 27.210 61.240 27.530 61.300 ;
        RECT 12.030 60.900 12.350 61.160 ;
        RECT 13.870 60.900 14.190 61.160 ;
        RECT 16.645 61.100 16.935 61.145 ;
        RECT 18.930 61.100 19.250 61.160 ;
        RECT 20.785 61.100 21.075 61.145 ;
        RECT 16.645 60.960 21.075 61.100 ;
        RECT 16.645 60.915 16.935 60.960 ;
        RECT 18.930 60.900 19.250 60.960 ;
        RECT 20.785 60.915 21.075 60.960 ;
        RECT 22.610 61.100 22.930 61.160 ;
        RECT 25.845 61.100 26.135 61.145 ;
        RECT 22.610 60.960 26.135 61.100 ;
        RECT 22.610 60.900 22.930 60.960 ;
        RECT 25.845 60.915 26.135 60.960 ;
        RECT 30.430 60.900 30.750 61.160 ;
        RECT 30.980 61.145 31.120 61.300 ;
        RECT 35.950 61.240 36.270 61.500 ;
        RECT 30.905 61.100 31.195 61.145 ;
        RECT 34.125 61.100 34.415 61.145 ;
        RECT 35.490 61.100 35.810 61.160 ;
        RECT 39.230 61.100 39.520 61.145 ;
        RECT 30.905 60.960 35.810 61.100 ;
        RECT 30.905 60.915 31.195 60.960 ;
        RECT 34.125 60.915 34.415 60.960 ;
        RECT 35.490 60.900 35.810 60.960 ;
        RECT 36.985 60.960 39.520 61.100 ;
        RECT 9.270 60.760 9.590 60.820 ;
        RECT 36.985 60.805 37.200 60.960 ;
        RECT 39.230 60.915 39.520 60.960 ;
        RECT 46.545 61.100 46.835 61.145 ;
        RECT 47.080 61.100 47.220 61.595 ;
        RECT 46.545 60.960 47.220 61.100 ;
        RECT 47.540 61.100 47.680 61.980 ;
        RECT 49.750 61.980 51.895 62.120 ;
        RECT 49.750 61.920 50.070 61.980 ;
        RECT 51.605 61.935 51.895 61.980 ;
        RECT 58.950 62.120 59.270 62.180 ;
        RECT 61.725 62.120 62.015 62.165 ;
        RECT 58.950 61.980 62.015 62.120 ;
        RECT 58.950 61.920 59.270 61.980 ;
        RECT 61.725 61.935 62.015 61.980 ;
        RECT 63.090 62.120 63.410 62.180 ;
        RECT 63.565 62.120 63.855 62.165 ;
        RECT 63.090 61.980 63.855 62.120 ;
        RECT 63.090 61.920 63.410 61.980 ;
        RECT 63.565 61.935 63.855 61.980 ;
        RECT 65.850 61.920 66.170 62.180 ;
        RECT 98.050 62.120 98.370 62.180 ;
        RECT 98.970 62.120 99.290 62.180 ;
        RECT 111.390 62.120 111.710 62.180 ;
        RECT 114.855 62.120 115.145 62.165 ;
        RECT 98.050 61.980 99.290 62.120 ;
        RECT 98.050 61.920 98.370 61.980 ;
        RECT 98.970 61.920 99.290 61.980 ;
        RECT 103.660 61.980 115.145 62.120 ;
        RECT 52.050 61.780 52.370 61.840 ;
        RECT 49.380 61.640 52.370 61.780 ;
        RECT 49.380 61.485 49.520 61.640 ;
        RECT 52.050 61.580 52.370 61.640 ;
        RECT 62.170 61.780 62.490 61.840 ;
        RECT 67.705 61.780 67.995 61.825 ;
        RECT 79.650 61.780 79.970 61.840 ;
        RECT 89.325 61.780 89.615 61.825 ;
        RECT 95.290 61.780 95.610 61.840 ;
        RECT 103.660 61.780 103.800 61.980 ;
        RECT 111.390 61.920 111.710 61.980 ;
        RECT 114.855 61.935 115.145 61.980 ;
        RECT 62.170 61.640 79.970 61.780 ;
        RECT 62.170 61.580 62.490 61.640 ;
        RECT 67.705 61.595 67.995 61.640 ;
        RECT 79.650 61.580 79.970 61.640 ;
        RECT 80.660 61.640 86.320 61.780 ;
        RECT 49.305 61.255 49.595 61.485 ;
        RECT 50.225 61.440 50.515 61.485 ;
        RECT 52.970 61.440 53.290 61.500 ;
        RECT 65.850 61.440 66.170 61.500 ;
        RECT 80.660 61.485 80.800 61.640 ;
        RECT 78.745 61.440 79.035 61.485 ;
        RECT 80.585 61.440 80.875 61.485 ;
        RECT 50.225 61.300 53.290 61.440 ;
        RECT 50.225 61.255 50.515 61.300 ;
        RECT 52.970 61.240 53.290 61.300 ;
        RECT 64.560 61.300 65.620 61.440 ;
        RECT 51.145 61.100 51.435 61.145 ;
        RECT 47.540 60.960 51.435 61.100 ;
        RECT 46.545 60.915 46.835 60.960 ;
        RECT 51.145 60.915 51.435 60.960 ;
        RECT 61.710 61.100 62.030 61.160 ;
        RECT 64.560 61.145 64.700 61.300 ;
        RECT 62.645 61.100 62.935 61.145 ;
        RECT 61.710 60.960 62.935 61.100 ;
        RECT 61.710 60.900 62.030 60.960 ;
        RECT 62.645 60.915 62.935 60.960 ;
        RECT 64.485 60.915 64.775 61.145 ;
        RECT 64.945 60.915 65.235 61.145 ;
        RECT 65.480 61.100 65.620 61.300 ;
        RECT 65.850 61.300 80.875 61.440 ;
        RECT 65.850 61.240 66.170 61.300 ;
        RECT 78.745 61.255 79.035 61.300 ;
        RECT 80.585 61.255 80.875 61.300 ;
        RECT 81.505 61.440 81.795 61.485 ;
        RECT 83.790 61.440 84.110 61.500 ;
        RECT 86.180 61.485 86.320 61.640 ;
        RECT 89.325 61.640 92.760 61.780 ;
        RECT 89.325 61.595 89.615 61.640 ;
        RECT 92.620 61.485 92.760 61.640 ;
        RECT 95.290 61.640 103.800 61.780 ;
        RECT 95.290 61.580 95.610 61.640 ;
        RECT 81.505 61.300 84.110 61.440 ;
        RECT 81.505 61.255 81.795 61.300 ;
        RECT 83.790 61.240 84.110 61.300 ;
        RECT 86.105 61.440 86.395 61.485 ;
        RECT 86.105 61.300 92.300 61.440 ;
        RECT 86.105 61.255 86.395 61.300 ;
        RECT 66.310 61.100 66.630 61.160 ;
        RECT 66.785 61.100 67.075 61.145 ;
        RECT 65.480 60.960 67.075 61.100 ;
        RECT 35.050 60.760 35.340 60.805 ;
        RECT 36.910 60.760 37.200 60.805 ;
        RECT 9.270 60.620 19.160 60.760 ;
        RECT 9.270 60.560 9.590 60.620 ;
        RECT 11.125 60.420 11.415 60.465 ;
        RECT 11.570 60.420 11.890 60.480 ;
        RECT 11.125 60.280 11.890 60.420 ;
        RECT 11.125 60.235 11.415 60.280 ;
        RECT 11.570 60.220 11.890 60.280 ;
        RECT 13.410 60.220 13.730 60.480 ;
        RECT 15.710 60.420 16.030 60.480 ;
        RECT 16.185 60.420 16.475 60.465 ;
        RECT 16.630 60.420 16.950 60.480 ;
        RECT 19.020 60.465 19.160 60.620 ;
        RECT 35.050 60.620 37.200 60.760 ;
        RECT 35.050 60.575 35.340 60.620 ;
        RECT 36.910 60.575 37.200 60.620 ;
        RECT 37.830 60.760 38.120 60.805 ;
        RECT 38.710 60.760 39.030 60.820 ;
        RECT 41.090 60.760 41.380 60.805 ;
        RECT 48.845 60.760 49.135 60.805 ;
        RECT 37.830 60.620 41.380 60.760 ;
        RECT 37.830 60.575 38.120 60.620 ;
        RECT 38.710 60.560 39.030 60.620 ;
        RECT 41.090 60.575 41.380 60.620 ;
        RECT 45.240 60.620 49.135 60.760 ;
        RECT 62.720 60.760 62.860 60.915 ;
        RECT 65.020 60.760 65.160 60.915 ;
        RECT 66.310 60.900 66.630 60.960 ;
        RECT 66.785 60.915 67.075 60.960 ;
        RECT 73.225 61.100 73.515 61.145 ;
        RECT 78.285 61.100 78.575 61.145 ;
        RECT 81.965 61.100 82.255 61.145 ;
        RECT 83.330 61.100 83.650 61.160 ;
        RECT 73.225 60.960 76.200 61.100 ;
        RECT 73.225 60.915 73.515 60.960 ;
        RECT 62.720 60.620 65.160 60.760 ;
        RECT 15.710 60.280 16.950 60.420 ;
        RECT 15.710 60.220 16.030 60.280 ;
        RECT 16.185 60.235 16.475 60.280 ;
        RECT 16.630 60.220 16.950 60.280 ;
        RECT 18.945 60.235 19.235 60.465 ;
        RECT 21.245 60.420 21.535 60.465 ;
        RECT 23.070 60.420 23.390 60.480 ;
        RECT 21.245 60.280 23.390 60.420 ;
        RECT 21.245 60.235 21.535 60.280 ;
        RECT 23.070 60.220 23.390 60.280 ;
        RECT 26.750 60.420 27.070 60.480 ;
        RECT 27.225 60.420 27.515 60.465 ;
        RECT 26.750 60.280 27.515 60.420 ;
        RECT 26.750 60.220 27.070 60.280 ;
        RECT 27.225 60.235 27.515 60.280 ;
        RECT 38.250 60.420 38.570 60.480 ;
        RECT 43.095 60.420 43.385 60.465 ;
        RECT 45.240 60.420 45.380 60.620 ;
        RECT 48.845 60.575 49.135 60.620 ;
        RECT 38.250 60.280 45.380 60.420 ;
        RECT 48.920 60.420 49.060 60.575 ;
        RECT 50.210 60.420 50.530 60.480 ;
        RECT 48.920 60.280 50.530 60.420 ;
        RECT 38.250 60.220 38.570 60.280 ;
        RECT 43.095 60.235 43.385 60.280 ;
        RECT 50.210 60.220 50.530 60.280 ;
        RECT 70.450 60.420 70.770 60.480 ;
        RECT 76.060 60.465 76.200 60.960 ;
        RECT 78.285 60.960 83.650 61.100 ;
        RECT 78.285 60.915 78.575 60.960 ;
        RECT 81.965 60.915 82.255 60.960 ;
        RECT 83.330 60.900 83.650 60.960 ;
        RECT 83.880 60.760 84.020 61.240 ;
        RECT 84.265 61.100 84.555 61.145 ;
        RECT 89.785 61.100 90.075 61.145 ;
        RECT 84.265 60.960 90.075 61.100 ;
        RECT 92.160 61.100 92.300 61.300 ;
        RECT 92.545 61.255 92.835 61.485 ;
        RECT 96.685 61.440 96.975 61.485 ;
        RECT 102.190 61.440 102.510 61.500 ;
        RECT 93.080 61.300 102.510 61.440 ;
        RECT 93.080 61.100 93.220 61.300 ;
        RECT 96.685 61.255 96.975 61.300 ;
        RECT 102.190 61.240 102.510 61.300 ;
        RECT 98.970 61.100 99.290 61.160 ;
        RECT 92.160 60.960 93.220 61.100 ;
        RECT 97.680 60.960 99.290 61.100 ;
        RECT 84.265 60.915 84.555 60.960 ;
        RECT 89.785 60.915 90.075 60.960 ;
        RECT 83.420 60.620 84.020 60.760 ;
        RECT 87.025 60.760 87.315 60.805 ;
        RECT 96.670 60.760 96.990 60.820 ;
        RECT 97.680 60.805 97.820 60.960 ;
        RECT 98.970 60.900 99.290 60.960 ;
        RECT 87.025 60.620 96.990 60.760 ;
        RECT 83.420 60.480 83.560 60.620 ;
        RECT 87.025 60.575 87.315 60.620 ;
        RECT 96.670 60.560 96.990 60.620 ;
        RECT 97.605 60.575 97.895 60.805 ;
        RECT 98.065 60.760 98.355 60.805 ;
        RECT 101.730 60.760 102.050 60.820 ;
        RECT 103.660 60.805 103.800 61.640 ;
        RECT 106.350 61.780 106.640 61.825 ;
        RECT 108.210 61.780 108.500 61.825 ;
        RECT 110.990 61.780 111.280 61.825 ;
        RECT 106.350 61.640 111.280 61.780 ;
        RECT 106.350 61.595 106.640 61.640 ;
        RECT 108.210 61.595 108.500 61.640 ;
        RECT 110.990 61.595 111.280 61.640 ;
        RECT 107.250 61.440 107.570 61.500 ;
        RECT 107.725 61.440 108.015 61.485 ;
        RECT 107.250 61.300 108.015 61.440 ;
        RECT 107.250 61.240 107.570 61.300 ;
        RECT 107.725 61.255 108.015 61.300 ;
        RECT 104.030 61.100 104.350 61.160 ;
        RECT 105.870 61.100 106.190 61.160 ;
        RECT 110.990 61.100 111.280 61.145 ;
        RECT 104.030 60.960 106.190 61.100 ;
        RECT 104.030 60.900 104.350 60.960 ;
        RECT 105.870 60.900 106.190 60.960 ;
        RECT 108.745 60.960 111.280 61.100 ;
        RECT 108.745 60.805 108.960 60.960 ;
        RECT 110.990 60.915 111.280 60.960 ;
        RECT 98.065 60.620 102.050 60.760 ;
        RECT 98.065 60.575 98.355 60.620 ;
        RECT 101.730 60.560 102.050 60.620 ;
        RECT 103.585 60.575 103.875 60.805 ;
        RECT 106.810 60.760 107.100 60.805 ;
        RECT 108.670 60.760 108.960 60.805 ;
        RECT 106.810 60.620 108.960 60.760 ;
        RECT 106.810 60.575 107.100 60.620 ;
        RECT 108.670 60.575 108.960 60.620 ;
        RECT 109.590 60.760 109.880 60.805 ;
        RECT 112.850 60.760 113.140 60.805 ;
        RECT 114.150 60.760 114.470 60.820 ;
        RECT 109.590 60.620 114.470 60.760 ;
        RECT 109.590 60.575 109.880 60.620 ;
        RECT 112.850 60.575 113.140 60.620 ;
        RECT 114.150 60.560 114.470 60.620 ;
        RECT 72.305 60.420 72.595 60.465 ;
        RECT 70.450 60.280 72.595 60.420 ;
        RECT 70.450 60.220 70.770 60.280 ;
        RECT 72.305 60.235 72.595 60.280 ;
        RECT 75.985 60.235 76.275 60.465 ;
        RECT 77.825 60.420 78.115 60.465 ;
        RECT 78.730 60.420 79.050 60.480 ;
        RECT 77.825 60.280 79.050 60.420 ;
        RECT 77.825 60.235 78.115 60.280 ;
        RECT 78.730 60.220 79.050 60.280 ;
        RECT 83.330 60.220 83.650 60.480 ;
        RECT 83.790 60.220 84.110 60.480 ;
        RECT 85.185 60.420 85.475 60.465 ;
        RECT 86.550 60.420 86.870 60.480 ;
        RECT 85.185 60.280 86.870 60.420 ;
        RECT 85.185 60.235 85.475 60.280 ;
        RECT 86.550 60.220 86.870 60.280 ;
        RECT 87.485 60.420 87.775 60.465 ;
        RECT 90.230 60.420 90.550 60.480 ;
        RECT 87.485 60.280 90.550 60.420 ;
        RECT 87.485 60.235 87.775 60.280 ;
        RECT 90.230 60.220 90.550 60.280 ;
        RECT 98.510 60.420 98.830 60.480 ;
        RECT 99.905 60.420 100.195 60.465 ;
        RECT 98.510 60.280 100.195 60.420 ;
        RECT 98.510 60.220 98.830 60.280 ;
        RECT 99.905 60.235 100.195 60.280 ;
        RECT 103.110 60.220 103.430 60.480 ;
        RECT 105.425 60.420 105.715 60.465 ;
        RECT 106.330 60.420 106.650 60.480 ;
        RECT 105.425 60.280 106.650 60.420 ;
        RECT 105.425 60.235 105.715 60.280 ;
        RECT 106.330 60.220 106.650 60.280 ;
        RECT 5.520 59.600 118.680 60.080 ;
        RECT 10.205 59.400 10.495 59.445 ;
        RECT 23.070 59.400 23.390 59.460 ;
        RECT 24.465 59.400 24.755 59.445 ;
        RECT 10.205 59.260 12.260 59.400 ;
        RECT 10.205 59.215 10.495 59.260 ;
        RECT 12.120 59.105 12.260 59.260 ;
        RECT 23.070 59.260 24.755 59.400 ;
        RECT 23.070 59.200 23.390 59.260 ;
        RECT 24.465 59.215 24.755 59.260 ;
        RECT 27.225 59.400 27.515 59.445 ;
        RECT 27.670 59.400 27.990 59.460 ;
        RECT 27.225 59.260 27.990 59.400 ;
        RECT 27.225 59.215 27.515 59.260 ;
        RECT 27.670 59.200 27.990 59.260 ;
        RECT 35.490 59.400 35.810 59.460 ;
        RECT 38.265 59.400 38.555 59.445 ;
        RECT 41.930 59.400 42.250 59.460 ;
        RECT 35.490 59.260 42.250 59.400 ;
        RECT 35.490 59.200 35.810 59.260 ;
        RECT 38.265 59.215 38.555 59.260 ;
        RECT 41.930 59.200 42.250 59.260 ;
        RECT 51.145 59.215 51.435 59.445 ;
        RECT 52.050 59.400 52.370 59.460 ;
        RECT 52.985 59.400 53.275 59.445 ;
        RECT 52.050 59.260 53.275 59.400 ;
        RECT 12.045 58.875 12.335 59.105 ;
        RECT 14.325 59.060 14.975 59.105 ;
        RECT 17.925 59.060 18.215 59.105 ;
        RECT 19.390 59.060 19.710 59.120 ;
        RECT 14.325 58.920 19.710 59.060 ;
        RECT 14.325 58.875 14.975 58.920 ;
        RECT 17.625 58.875 18.215 58.920 ;
        RECT 9.270 58.520 9.590 58.780 ;
        RECT 11.130 58.720 11.420 58.765 ;
        RECT 12.965 58.720 13.255 58.765 ;
        RECT 16.545 58.720 16.835 58.765 ;
        RECT 11.130 58.580 16.835 58.720 ;
        RECT 11.130 58.535 11.420 58.580 ;
        RECT 12.965 58.535 13.255 58.580 ;
        RECT 16.545 58.535 16.835 58.580 ;
        RECT 17.625 58.560 17.915 58.875 ;
        RECT 19.390 58.860 19.710 58.920 ;
        RECT 21.230 58.860 21.550 59.120 ;
        RECT 24.005 59.060 24.295 59.105 ;
        RECT 26.750 59.060 27.070 59.120 ;
        RECT 29.065 59.060 29.355 59.105 ;
        RECT 24.005 58.920 29.355 59.060 ;
        RECT 24.005 58.875 24.295 58.920 ;
        RECT 26.750 58.860 27.070 58.920 ;
        RECT 29.065 58.875 29.355 58.920 ;
        RECT 29.525 59.060 29.815 59.105 ;
        RECT 34.570 59.060 34.890 59.120 ;
        RECT 29.525 58.920 34.890 59.060 ;
        RECT 29.525 58.875 29.815 58.920 ;
        RECT 34.570 58.860 34.890 58.920 ;
        RECT 19.850 58.520 20.170 58.780 ;
        RECT 20.310 58.720 20.630 58.780 ;
        RECT 20.310 58.580 23.760 58.720 ;
        RECT 20.310 58.520 20.630 58.580 ;
        RECT 8.350 58.380 8.670 58.440 ;
        RECT 10.665 58.380 10.955 58.425 ;
        RECT 8.350 58.240 10.955 58.380 ;
        RECT 8.350 58.180 8.670 58.240 ;
        RECT 10.665 58.195 10.955 58.240 ;
        RECT 19.405 58.380 19.695 58.425 ;
        RECT 22.610 58.380 22.930 58.440 ;
        RECT 23.620 58.425 23.760 58.580 ;
        RECT 31.810 58.520 32.130 58.780 ;
        RECT 47.465 58.720 47.755 58.765 ;
        RECT 49.750 58.720 50.070 58.780 ;
        RECT 47.465 58.580 50.070 58.720 ;
        RECT 47.465 58.535 47.755 58.580 ;
        RECT 49.750 58.520 50.070 58.580 ;
        RECT 50.685 58.720 50.975 58.765 ;
        RECT 51.220 58.720 51.360 59.215 ;
        RECT 52.050 59.200 52.370 59.260 ;
        RECT 52.985 59.215 53.275 59.260 ;
        RECT 65.405 59.400 65.695 59.445 ;
        RECT 65.850 59.400 66.170 59.460 ;
        RECT 65.405 59.260 66.170 59.400 ;
        RECT 65.405 59.215 65.695 59.260 ;
        RECT 65.850 59.200 66.170 59.260 ;
        RECT 77.825 59.400 78.115 59.445 ;
        RECT 80.110 59.400 80.430 59.460 ;
        RECT 77.825 59.260 80.430 59.400 ;
        RECT 77.825 59.215 78.115 59.260 ;
        RECT 80.110 59.200 80.430 59.260 ;
        RECT 96.670 59.200 96.990 59.460 ;
        RECT 97.130 59.200 97.450 59.460 ;
        RECT 53.890 58.860 54.210 59.120 ;
        RECT 57.570 59.060 57.890 59.120 ;
        RECT 67.705 59.060 67.995 59.105 ;
        RECT 57.570 58.920 67.995 59.060 ;
        RECT 57.570 58.860 57.890 58.920 ;
        RECT 67.705 58.875 67.995 58.920 ;
        RECT 50.685 58.580 51.360 58.720 ;
        RECT 53.445 58.720 53.735 58.765 ;
        RECT 53.980 58.720 54.120 58.860 ;
        RECT 59.870 58.720 60.190 58.780 ;
        RECT 53.445 58.580 60.190 58.720 ;
        RECT 50.685 58.535 50.975 58.580 ;
        RECT 53.445 58.535 53.735 58.580 ;
        RECT 59.870 58.520 60.190 58.580 ;
        RECT 64.025 58.720 64.315 58.765 ;
        RECT 64.470 58.720 64.790 58.780 ;
        RECT 64.025 58.580 64.790 58.720 ;
        RECT 64.025 58.535 64.315 58.580 ;
        RECT 64.470 58.520 64.790 58.580 ;
        RECT 66.325 58.720 66.615 58.765 ;
        RECT 66.325 58.580 67.460 58.720 ;
        RECT 66.325 58.535 66.615 58.580 ;
        RECT 19.405 58.240 22.930 58.380 ;
        RECT 19.405 58.195 19.695 58.240 ;
        RECT 22.610 58.180 22.930 58.240 ;
        RECT 23.545 58.380 23.835 58.425 ;
        RECT 30.445 58.380 30.735 58.425 ;
        RECT 39.170 58.380 39.490 58.440 ;
        RECT 23.545 58.240 39.490 58.380 ;
        RECT 23.545 58.195 23.835 58.240 ;
        RECT 30.445 58.195 30.735 58.240 ;
        RECT 39.170 58.180 39.490 58.240 ;
        RECT 54.350 58.180 54.670 58.440 ;
        RECT 11.535 58.040 11.825 58.085 ;
        RECT 13.425 58.040 13.715 58.085 ;
        RECT 16.545 58.040 16.835 58.085 ;
        RECT 11.535 57.900 16.835 58.040 ;
        RECT 11.535 57.855 11.825 57.900 ;
        RECT 13.425 57.855 13.715 57.900 ;
        RECT 16.545 57.855 16.835 57.900 ;
        RECT 23.990 58.040 24.310 58.100 ;
        RECT 26.305 58.040 26.595 58.085 ;
        RECT 23.990 57.900 26.595 58.040 ;
        RECT 23.990 57.840 24.310 57.900 ;
        RECT 26.305 57.855 26.595 57.900 ;
        RECT 27.300 57.900 62.170 58.040 ;
        RECT 19.850 57.700 20.170 57.760 ;
        RECT 27.300 57.700 27.440 57.900 ;
        RECT 19.850 57.560 27.440 57.700 ;
        RECT 45.150 57.700 45.470 57.760 ;
        RECT 46.545 57.700 46.835 57.745 ;
        RECT 45.150 57.560 46.835 57.700 ;
        RECT 19.850 57.500 20.170 57.560 ;
        RECT 45.150 57.500 45.470 57.560 ;
        RECT 46.545 57.515 46.835 57.560 ;
        RECT 49.765 57.700 50.055 57.745 ;
        RECT 50.210 57.700 50.530 57.760 ;
        RECT 49.765 57.560 50.530 57.700 ;
        RECT 62.030 57.700 62.170 57.900 ;
        RECT 67.320 57.700 67.460 58.580 ;
        RECT 67.780 58.380 67.920 58.875 ;
        RECT 70.450 58.860 70.770 59.120 ;
        RECT 72.745 59.060 73.395 59.105 ;
        RECT 74.130 59.060 74.450 59.120 ;
        RECT 76.345 59.060 76.635 59.105 ;
        RECT 72.745 58.920 76.635 59.060 ;
        RECT 72.745 58.875 73.395 58.920 ;
        RECT 74.130 58.860 74.450 58.920 ;
        RECT 76.045 58.875 76.635 58.920 ;
        RECT 86.550 59.060 86.870 59.120 ;
        RECT 89.325 59.060 89.615 59.105 ;
        RECT 86.550 58.920 89.615 59.060 ;
        RECT 69.070 58.520 69.390 58.780 ;
        RECT 69.550 58.720 69.840 58.765 ;
        RECT 71.385 58.720 71.675 58.765 ;
        RECT 74.965 58.720 75.255 58.765 ;
        RECT 69.550 58.580 75.255 58.720 ;
        RECT 69.550 58.535 69.840 58.580 ;
        RECT 71.385 58.535 71.675 58.580 ;
        RECT 74.965 58.535 75.255 58.580 ;
        RECT 76.045 58.560 76.335 58.875 ;
        RECT 86.550 58.860 86.870 58.920 ;
        RECT 89.325 58.875 89.615 58.920 ;
        RECT 91.605 59.060 92.255 59.105 ;
        RECT 95.205 59.060 95.495 59.105 ;
        RECT 91.605 58.920 95.495 59.060 ;
        RECT 91.605 58.875 92.255 58.920 ;
        RECT 94.905 58.875 95.495 58.920 ;
        RECT 98.625 59.060 98.915 59.105 ;
        RECT 101.865 59.060 102.515 59.105 ;
        RECT 98.625 58.920 102.515 59.060 ;
        RECT 98.625 58.875 99.215 58.920 ;
        RECT 101.865 58.875 102.515 58.920 ;
        RECT 104.030 59.060 104.350 59.120 ;
        RECT 104.030 58.920 106.100 59.060 ;
        RECT 94.905 58.780 95.195 58.875 ;
        RECT 79.205 58.535 79.495 58.765 ;
        RECT 79.650 58.720 79.970 58.780 ;
        RECT 81.505 58.720 81.795 58.765 ;
        RECT 79.650 58.580 81.795 58.720 ;
        RECT 72.290 58.380 72.610 58.440 ;
        RECT 67.780 58.240 72.610 58.380 ;
        RECT 79.280 58.380 79.420 58.535 ;
        RECT 79.650 58.520 79.970 58.580 ;
        RECT 81.505 58.535 81.795 58.580 ;
        RECT 83.790 58.720 84.110 58.780 ;
        RECT 86.105 58.720 86.395 58.765 ;
        RECT 83.790 58.580 86.395 58.720 ;
        RECT 83.790 58.520 84.110 58.580 ;
        RECT 86.105 58.535 86.395 58.580 ;
        RECT 88.410 58.720 88.700 58.765 ;
        RECT 90.245 58.720 90.535 58.765 ;
        RECT 93.825 58.720 94.115 58.765 ;
        RECT 88.410 58.580 94.115 58.720 ;
        RECT 88.410 58.535 88.700 58.580 ;
        RECT 90.245 58.535 90.535 58.580 ;
        RECT 93.825 58.535 94.115 58.580 ;
        RECT 94.830 58.560 95.195 58.780 ;
        RECT 98.925 58.780 99.215 58.875 ;
        RECT 104.030 58.860 104.350 58.920 ;
        RECT 105.960 58.780 106.100 58.920 ;
        RECT 98.925 58.560 99.290 58.780 ;
        RECT 94.830 58.520 95.150 58.560 ;
        RECT 98.970 58.520 99.290 58.560 ;
        RECT 100.005 58.720 100.295 58.765 ;
        RECT 103.585 58.720 103.875 58.765 ;
        RECT 105.420 58.720 105.710 58.765 ;
        RECT 100.005 58.580 105.710 58.720 ;
        RECT 100.005 58.535 100.295 58.580 ;
        RECT 103.585 58.535 103.875 58.580 ;
        RECT 105.420 58.535 105.710 58.580 ;
        RECT 105.870 58.520 106.190 58.780 ;
        RECT 106.330 58.520 106.650 58.780 ;
        RECT 83.345 58.380 83.635 58.425 ;
        RECT 79.280 58.240 83.635 58.380 ;
        RECT 72.290 58.180 72.610 58.240 ;
        RECT 83.345 58.195 83.635 58.240 ;
        RECT 87.945 58.380 88.235 58.425 ;
        RECT 96.210 58.380 96.530 58.440 ;
        RECT 104.030 58.380 104.350 58.440 ;
        RECT 87.945 58.240 104.350 58.380 ;
        RECT 87.945 58.195 88.235 58.240 ;
        RECT 69.955 58.040 70.245 58.085 ;
        RECT 71.845 58.040 72.135 58.085 ;
        RECT 74.965 58.040 75.255 58.085 ;
        RECT 69.955 57.900 75.255 58.040 ;
        RECT 69.955 57.855 70.245 57.900 ;
        RECT 71.845 57.855 72.135 57.900 ;
        RECT 74.965 57.855 75.255 57.900 ;
        RECT 75.510 58.040 75.830 58.100 ;
        RECT 88.020 58.040 88.160 58.195 ;
        RECT 96.210 58.180 96.530 58.240 ;
        RECT 104.030 58.180 104.350 58.240 ;
        RECT 104.490 58.180 104.810 58.440 ;
        RECT 75.510 57.900 88.160 58.040 ;
        RECT 88.815 58.040 89.105 58.085 ;
        RECT 90.705 58.040 90.995 58.085 ;
        RECT 93.825 58.040 94.115 58.085 ;
        RECT 88.815 57.900 94.115 58.040 ;
        RECT 75.510 57.840 75.830 57.900 ;
        RECT 88.815 57.855 89.105 57.900 ;
        RECT 90.705 57.855 90.995 57.900 ;
        RECT 93.825 57.855 94.115 57.900 ;
        RECT 100.005 58.040 100.295 58.085 ;
        RECT 103.125 58.040 103.415 58.085 ;
        RECT 105.015 58.040 105.305 58.085 ;
        RECT 100.005 57.900 105.305 58.040 ;
        RECT 100.005 57.855 100.295 57.900 ;
        RECT 103.125 57.855 103.415 57.900 ;
        RECT 105.015 57.855 105.305 57.900 ;
        RECT 71.370 57.700 71.690 57.760 ;
        RECT 62.030 57.560 71.690 57.700 ;
        RECT 49.765 57.515 50.055 57.560 ;
        RECT 50.210 57.500 50.530 57.560 ;
        RECT 71.370 57.500 71.690 57.560 ;
        RECT 78.270 57.500 78.590 57.760 ;
        RECT 81.950 57.500 82.270 57.760 ;
        RECT 107.265 57.700 107.555 57.745 ;
        RECT 108.170 57.700 108.490 57.760 ;
        RECT 107.265 57.560 108.490 57.700 ;
        RECT 107.265 57.515 107.555 57.560 ;
        RECT 108.170 57.500 108.490 57.560 ;
        RECT 5.520 56.880 118.680 57.360 ;
        RECT 9.680 56.680 9.970 56.725 ;
        RECT 11.570 56.680 11.890 56.740 ;
        RECT 9.680 56.540 11.890 56.680 ;
        RECT 9.680 56.495 9.970 56.540 ;
        RECT 11.570 56.480 11.890 56.540 ;
        RECT 18.930 56.480 19.250 56.740 ;
        RECT 35.965 56.680 36.255 56.725 ;
        RECT 36.410 56.680 36.730 56.740 ;
        RECT 35.965 56.540 36.730 56.680 ;
        RECT 35.965 56.495 36.255 56.540 ;
        RECT 36.410 56.480 36.730 56.540 ;
        RECT 41.010 56.680 41.330 56.740 ;
        RECT 52.970 56.680 53.290 56.740 ;
        RECT 57.355 56.680 57.645 56.725 ;
        RECT 59.870 56.680 60.190 56.740 ;
        RECT 41.010 56.540 54.580 56.680 ;
        RECT 41.010 56.480 41.330 56.540 ;
        RECT 52.970 56.480 53.290 56.540 ;
        RECT 54.440 56.400 54.580 56.540 ;
        RECT 57.355 56.540 60.190 56.680 ;
        RECT 57.355 56.495 57.645 56.540 ;
        RECT 59.870 56.480 60.190 56.540 ;
        RECT 64.010 56.680 64.330 56.740 ;
        RECT 66.325 56.680 66.615 56.725 ;
        RECT 64.010 56.540 66.615 56.680 ;
        RECT 64.010 56.480 64.330 56.540 ;
        RECT 66.325 56.495 66.615 56.540 ;
        RECT 74.130 56.480 74.450 56.740 ;
        RECT 83.330 56.680 83.650 56.740 ;
        RECT 85.645 56.680 85.935 56.725 ;
        RECT 83.330 56.540 85.935 56.680 ;
        RECT 83.330 56.480 83.650 56.540 ;
        RECT 85.645 56.495 85.935 56.540 ;
        RECT 9.235 56.340 9.525 56.385 ;
        RECT 11.125 56.340 11.415 56.385 ;
        RECT 14.245 56.340 14.535 56.385 ;
        RECT 9.235 56.200 14.535 56.340 ;
        RECT 9.235 56.155 9.525 56.200 ;
        RECT 11.125 56.155 11.415 56.200 ;
        RECT 14.245 56.155 14.535 56.200 ;
        RECT 17.105 56.340 17.395 56.385 ;
        RECT 20.770 56.340 21.090 56.400 ;
        RECT 17.105 56.200 21.090 56.340 ;
        RECT 17.105 56.155 17.395 56.200 ;
        RECT 20.770 56.140 21.090 56.200 ;
        RECT 22.150 56.340 22.470 56.400 ;
        RECT 23.990 56.340 24.310 56.400 ;
        RECT 22.150 56.200 24.310 56.340 ;
        RECT 22.150 56.140 22.470 56.200 ;
        RECT 23.990 56.140 24.310 56.200 ;
        RECT 26.770 56.340 27.060 56.385 ;
        RECT 28.630 56.340 28.920 56.385 ;
        RECT 31.410 56.340 31.700 56.385 ;
        RECT 26.770 56.200 31.700 56.340 ;
        RECT 26.770 56.155 27.060 56.200 ;
        RECT 28.630 56.155 28.920 56.200 ;
        RECT 31.410 56.155 31.700 56.200 ;
        RECT 48.850 56.340 49.140 56.385 ;
        RECT 50.710 56.340 51.000 56.385 ;
        RECT 53.490 56.340 53.780 56.385 ;
        RECT 48.850 56.200 53.780 56.340 ;
        RECT 48.850 56.155 49.140 56.200 ;
        RECT 50.710 56.155 51.000 56.200 ;
        RECT 53.490 56.155 53.780 56.200 ;
        RECT 54.350 56.340 54.670 56.400 ;
        RECT 63.105 56.340 63.395 56.385 ;
        RECT 54.350 56.200 63.395 56.340 ;
        RECT 54.350 56.140 54.670 56.200 ;
        RECT 63.105 56.155 63.395 56.200 ;
        RECT 77.775 56.340 78.065 56.385 ;
        RECT 79.665 56.340 79.955 56.385 ;
        RECT 82.785 56.340 83.075 56.385 ;
        RECT 77.775 56.200 83.075 56.340 ;
        RECT 77.775 56.155 78.065 56.200 ;
        RECT 79.665 56.155 79.955 56.200 ;
        RECT 82.785 56.155 83.075 56.200 ;
        RECT 21.230 56.000 21.550 56.060 ;
        RECT 26.305 56.000 26.595 56.045 ;
        RECT 27.210 56.000 27.530 56.060 ;
        RECT 8.440 55.860 27.530 56.000 ;
        RECT 8.440 55.720 8.580 55.860 ;
        RECT 21.230 55.800 21.550 55.860 ;
        RECT 26.305 55.815 26.595 55.860 ;
        RECT 27.210 55.800 27.530 55.860 ;
        RECT 28.130 55.800 28.450 56.060 ;
        RECT 34.570 56.000 34.890 56.060 ;
        RECT 35.275 56.000 35.565 56.045 ;
        RECT 34.570 55.860 38.020 56.000 ;
        RECT 34.570 55.800 34.890 55.860 ;
        RECT 35.275 55.815 35.565 55.860 ;
        RECT 8.350 55.460 8.670 55.720 ;
        RECT 8.830 55.660 9.120 55.705 ;
        RECT 10.665 55.660 10.955 55.705 ;
        RECT 14.245 55.660 14.535 55.705 ;
        RECT 8.830 55.520 14.535 55.660 ;
        RECT 8.830 55.475 9.120 55.520 ;
        RECT 10.665 55.475 10.955 55.520 ;
        RECT 14.245 55.475 14.535 55.520 ;
        RECT 12.025 55.320 12.675 55.365 ;
        RECT 13.410 55.320 13.730 55.380 ;
        RECT 15.325 55.365 15.615 55.680 ;
        RECT 20.770 55.660 21.090 55.720 ;
        RECT 21.705 55.660 21.995 55.705 ;
        RECT 20.770 55.520 21.995 55.660 ;
        RECT 20.770 55.460 21.090 55.520 ;
        RECT 21.705 55.475 21.995 55.520 ;
        RECT 22.150 55.660 22.470 55.720 ;
        RECT 37.880 55.705 38.020 55.860 ;
        RECT 38.250 55.800 38.570 56.060 ;
        RECT 39.170 56.000 39.490 56.060 ;
        RECT 41.010 56.000 41.330 56.060 ;
        RECT 39.170 55.860 41.330 56.000 ;
        RECT 39.170 55.800 39.490 55.860 ;
        RECT 41.010 55.800 41.330 55.860 ;
        RECT 41.930 56.000 42.250 56.060 ;
        RECT 48.385 56.000 48.675 56.045 ;
        RECT 41.930 55.860 48.675 56.000 ;
        RECT 41.930 55.800 42.250 55.860 ;
        RECT 48.385 55.815 48.675 55.860 ;
        RECT 50.210 55.800 50.530 56.060 ;
        RECT 58.030 56.000 58.350 56.060 ;
        RECT 58.950 56.000 59.270 56.060 ;
        RECT 60.805 56.000 61.095 56.045 ;
        RECT 50.760 55.860 54.120 56.000 ;
        RECT 25.385 55.660 25.675 55.705 ;
        RECT 31.410 55.660 31.700 55.705 ;
        RECT 22.150 55.520 25.675 55.660 ;
        RECT 22.150 55.460 22.470 55.520 ;
        RECT 25.385 55.475 25.675 55.520 ;
        RECT 29.165 55.520 31.700 55.660 ;
        RECT 29.165 55.365 29.380 55.520 ;
        RECT 31.410 55.475 31.700 55.520 ;
        RECT 37.805 55.475 38.095 55.705 ;
        RECT 44.230 55.660 44.550 55.720 ;
        RECT 45.625 55.660 45.915 55.705 ;
        RECT 47.005 55.660 47.295 55.705 ;
        RECT 44.230 55.520 47.295 55.660 ;
        RECT 44.230 55.460 44.550 55.520 ;
        RECT 45.625 55.475 45.915 55.520 ;
        RECT 47.005 55.475 47.295 55.520 ;
        RECT 47.465 55.660 47.755 55.705 ;
        RECT 50.760 55.660 50.900 55.860 ;
        RECT 53.490 55.660 53.780 55.705 ;
        RECT 47.465 55.520 50.900 55.660 ;
        RECT 51.245 55.520 53.780 55.660 ;
        RECT 47.465 55.475 47.755 55.520 ;
        RECT 15.325 55.320 15.915 55.365 ;
        RECT 12.025 55.180 15.915 55.320 ;
        RECT 12.025 55.135 12.675 55.180 ;
        RECT 13.410 55.120 13.730 55.180 ;
        RECT 15.625 55.135 15.915 55.180 ;
        RECT 27.230 55.320 27.520 55.365 ;
        RECT 29.090 55.320 29.380 55.365 ;
        RECT 27.230 55.180 29.380 55.320 ;
        RECT 27.230 55.135 27.520 55.180 ;
        RECT 29.090 55.135 29.380 55.180 ;
        RECT 30.010 55.320 30.300 55.365 ;
        RECT 32.730 55.320 33.050 55.380 ;
        RECT 33.270 55.320 33.560 55.365 ;
        RECT 30.010 55.180 33.560 55.320 ;
        RECT 30.010 55.135 30.300 55.180 ;
        RECT 32.730 55.120 33.050 55.180 ;
        RECT 33.270 55.135 33.560 55.180 ;
        RECT 46.085 55.320 46.375 55.365 ;
        RECT 48.830 55.320 49.150 55.380 ;
        RECT 51.245 55.365 51.460 55.520 ;
        RECT 53.490 55.475 53.780 55.520 ;
        RECT 46.085 55.180 49.150 55.320 ;
        RECT 46.085 55.135 46.375 55.180 ;
        RECT 48.830 55.120 49.150 55.180 ;
        RECT 49.310 55.320 49.600 55.365 ;
        RECT 51.170 55.320 51.460 55.365 ;
        RECT 49.310 55.180 51.460 55.320 ;
        RECT 49.310 55.135 49.600 55.180 ;
        RECT 51.170 55.135 51.460 55.180 ;
        RECT 52.090 55.320 52.380 55.365 ;
        RECT 53.980 55.320 54.120 55.860 ;
        RECT 58.030 55.860 61.095 56.000 ;
        RECT 58.030 55.800 58.350 55.860 ;
        RECT 58.950 55.800 59.270 55.860 ;
        RECT 60.805 55.815 61.095 55.860 ;
        RECT 61.725 56.000 62.015 56.045 ;
        RECT 66.310 56.000 66.630 56.060 ;
        RECT 61.725 55.860 66.630 56.000 ;
        RECT 61.725 55.815 62.015 55.860 ;
        RECT 66.310 55.800 66.630 55.860 ;
        RECT 69.070 56.000 69.390 56.060 ;
        RECT 75.510 56.000 75.830 56.060 ;
        RECT 76.905 56.000 77.195 56.045 ;
        RECT 69.070 55.860 77.195 56.000 ;
        RECT 69.070 55.800 69.390 55.860 ;
        RECT 75.510 55.800 75.830 55.860 ;
        RECT 76.905 55.815 77.195 55.860 ;
        RECT 78.270 55.800 78.590 56.060 ;
        RECT 78.730 56.000 79.050 56.060 ;
        RECT 85.720 56.000 85.860 56.495 ;
        RECT 90.230 56.480 90.550 56.740 ;
        RECT 94.830 56.480 95.150 56.740 ;
        RECT 100.365 56.680 100.655 56.725 ;
        RECT 104.490 56.680 104.810 56.740 ;
        RECT 100.365 56.540 104.810 56.680 ;
        RECT 100.365 56.495 100.655 56.540 ;
        RECT 104.490 56.480 104.810 56.540 ;
        RECT 90.705 56.340 90.995 56.385 ;
        RECT 103.110 56.340 103.430 56.400 ;
        RECT 87.560 56.200 103.430 56.340 ;
        RECT 87.025 56.000 87.315 56.045 ;
        RECT 78.730 55.860 84.480 56.000 ;
        RECT 85.720 55.860 87.315 56.000 ;
        RECT 78.730 55.800 79.050 55.860 ;
        RECT 60.345 55.660 60.635 55.705 ;
        RECT 59.500 55.520 60.635 55.660 ;
        RECT 55.350 55.320 55.640 55.365 ;
        RECT 52.090 55.180 55.640 55.320 ;
        RECT 52.090 55.135 52.380 55.180 ;
        RECT 55.350 55.135 55.640 55.180 ;
        RECT 22.610 54.780 22.930 55.040 ;
        RECT 59.500 54.980 59.640 55.520 ;
        RECT 60.345 55.475 60.635 55.520 ;
        RECT 62.170 55.460 62.490 55.720 ;
        RECT 64.470 55.460 64.790 55.720 ;
        RECT 65.865 55.660 66.155 55.705 ;
        RECT 70.465 55.660 70.755 55.705 ;
        RECT 71.370 55.660 71.690 55.720 ;
        RECT 65.865 55.520 71.690 55.660 ;
        RECT 65.865 55.475 66.155 55.520 ;
        RECT 70.465 55.475 70.755 55.520 ;
        RECT 71.370 55.460 71.690 55.520 ;
        RECT 71.845 55.660 72.135 55.705 ;
        RECT 73.685 55.660 73.975 55.705 ;
        RECT 71.845 55.520 73.975 55.660 ;
        RECT 71.845 55.475 72.135 55.520 ;
        RECT 73.685 55.475 73.975 55.520 ;
        RECT 77.370 55.660 77.660 55.705 ;
        RECT 79.205 55.660 79.495 55.705 ;
        RECT 82.785 55.660 83.075 55.705 ;
        RECT 77.370 55.520 83.075 55.660 ;
        RECT 77.370 55.475 77.660 55.520 ;
        RECT 79.205 55.475 79.495 55.520 ;
        RECT 82.785 55.475 83.075 55.520 ;
        RECT 59.885 55.320 60.175 55.365 ;
        RECT 64.560 55.320 64.700 55.460 ;
        RECT 59.885 55.180 64.700 55.320 ;
        RECT 73.760 55.320 73.900 55.475 ;
        RECT 79.650 55.320 79.970 55.380 ;
        RECT 80.565 55.320 81.215 55.365 ;
        RECT 81.950 55.320 82.270 55.380 ;
        RECT 83.865 55.365 84.155 55.680 ;
        RECT 84.340 55.660 84.480 55.860 ;
        RECT 87.025 55.815 87.315 55.860 ;
        RECT 87.560 55.660 87.700 56.200 ;
        RECT 90.705 56.155 90.995 56.200 ;
        RECT 103.110 56.140 103.430 56.200 ;
        RECT 103.685 56.340 103.975 56.385 ;
        RECT 106.805 56.340 107.095 56.385 ;
        RECT 108.695 56.340 108.985 56.385 ;
        RECT 103.685 56.200 108.985 56.340 ;
        RECT 103.685 56.155 103.975 56.200 ;
        RECT 106.805 56.155 107.095 56.200 ;
        RECT 108.695 56.155 108.985 56.200 ;
        RECT 89.770 56.000 90.090 56.060 ;
        RECT 93.465 56.000 93.755 56.045 ;
        RECT 100.825 56.000 101.115 56.045 ;
        RECT 89.770 55.860 101.115 56.000 ;
        RECT 89.770 55.800 90.090 55.860 ;
        RECT 93.465 55.815 93.755 55.860 ;
        RECT 100.825 55.815 101.115 55.860 ;
        RECT 105.870 56.000 106.190 56.060 ;
        RECT 109.565 56.000 109.855 56.045 ;
        RECT 105.870 55.860 109.855 56.000 ;
        RECT 105.870 55.800 106.190 55.860 ;
        RECT 109.565 55.815 109.855 55.860 ;
        RECT 84.340 55.520 87.700 55.660 ;
        RECT 95.305 55.475 95.595 55.705 ;
        RECT 96.210 55.660 96.530 55.720 ;
        RECT 96.685 55.660 96.975 55.705 ;
        RECT 96.210 55.520 96.975 55.660 ;
        RECT 83.865 55.320 84.455 55.365 ;
        RECT 95.380 55.320 95.520 55.475 ;
        RECT 96.210 55.460 96.530 55.520 ;
        RECT 96.685 55.475 96.975 55.520 ;
        RECT 98.510 55.660 98.830 55.720 ;
        RECT 99.445 55.660 99.735 55.705 ;
        RECT 98.510 55.520 99.735 55.660 ;
        RECT 98.510 55.460 98.830 55.520 ;
        RECT 99.445 55.475 99.735 55.520 ;
        RECT 97.130 55.320 97.450 55.380 ;
        RECT 102.605 55.365 102.895 55.680 ;
        RECT 103.685 55.660 103.975 55.705 ;
        RECT 107.265 55.660 107.555 55.705 ;
        RECT 109.100 55.660 109.390 55.705 ;
        RECT 103.685 55.520 109.390 55.660 ;
        RECT 103.685 55.475 103.975 55.520 ;
        RECT 107.265 55.475 107.555 55.520 ;
        RECT 109.100 55.475 109.390 55.520 ;
        RECT 73.760 55.180 80.340 55.320 ;
        RECT 59.885 55.135 60.175 55.180 ;
        RECT 79.650 55.120 79.970 55.180 ;
        RECT 62.630 54.980 62.950 55.040 ;
        RECT 59.500 54.840 62.950 54.980 ;
        RECT 80.200 54.980 80.340 55.180 ;
        RECT 80.565 55.180 84.455 55.320 ;
        RECT 80.565 55.135 81.215 55.180 ;
        RECT 81.950 55.120 82.270 55.180 ;
        RECT 84.165 55.135 84.455 55.180 ;
        RECT 84.800 55.180 97.450 55.320 ;
        RECT 84.800 54.980 84.940 55.180 ;
        RECT 97.130 55.120 97.450 55.180 ;
        RECT 102.305 55.320 102.895 55.365 ;
        RECT 103.110 55.320 103.430 55.380 ;
        RECT 105.545 55.320 106.195 55.365 ;
        RECT 102.305 55.180 106.195 55.320 ;
        RECT 102.305 55.135 102.595 55.180 ;
        RECT 103.110 55.120 103.430 55.180 ;
        RECT 105.545 55.135 106.195 55.180 ;
        RECT 108.170 55.120 108.490 55.380 ;
        RECT 80.200 54.840 84.940 54.980 ;
        RECT 62.630 54.780 62.950 54.840 ;
        RECT 5.520 54.160 118.680 54.640 ;
        RECT 10.665 53.960 10.955 54.005 ;
        RECT 19.850 53.960 20.170 54.020 ;
        RECT 10.665 53.820 20.170 53.960 ;
        RECT 10.665 53.775 10.955 53.820 ;
        RECT 19.850 53.760 20.170 53.820 ;
        RECT 20.325 53.960 20.615 54.005 ;
        RECT 22.150 53.960 22.470 54.020 ;
        RECT 20.325 53.820 22.470 53.960 ;
        RECT 20.325 53.775 20.615 53.820 ;
        RECT 22.150 53.760 22.470 53.820 ;
        RECT 29.985 53.960 30.275 54.005 ;
        RECT 30.430 53.960 30.750 54.020 ;
        RECT 29.985 53.820 30.750 53.960 ;
        RECT 29.985 53.775 30.275 53.820 ;
        RECT 30.430 53.760 30.750 53.820 ;
        RECT 49.750 53.960 50.070 54.020 ;
        RECT 52.985 53.960 53.275 54.005 ;
        RECT 49.750 53.820 53.275 53.960 ;
        RECT 49.750 53.760 50.070 53.820 ;
        RECT 52.985 53.775 53.275 53.820 ;
        RECT 53.890 53.960 54.210 54.020 ;
        RECT 54.825 53.960 55.115 54.005 ;
        RECT 53.890 53.820 55.115 53.960 ;
        RECT 53.890 53.760 54.210 53.820 ;
        RECT 54.825 53.775 55.115 53.820 ;
        RECT 55.285 53.960 55.575 54.005 ;
        RECT 56.650 53.960 56.970 54.020 ;
        RECT 55.285 53.820 56.970 53.960 ;
        RECT 55.285 53.775 55.575 53.820 ;
        RECT 22.610 53.620 22.930 53.680 ;
        RECT 12.580 53.480 22.930 53.620 ;
        RECT 5.130 53.280 5.450 53.340 ;
        RECT 12.580 53.325 12.720 53.480 ;
        RECT 22.610 53.420 22.930 53.480 ;
        RECT 24.905 53.620 25.555 53.665 ;
        RECT 25.830 53.620 26.150 53.680 ;
        RECT 28.505 53.620 28.795 53.665 ;
        RECT 24.905 53.480 28.795 53.620 ;
        RECT 24.905 53.435 25.555 53.480 ;
        RECT 25.830 53.420 26.150 53.480 ;
        RECT 28.205 53.435 28.795 53.480 ;
        RECT 44.250 53.620 44.540 53.665 ;
        RECT 46.110 53.620 46.400 53.665 ;
        RECT 44.250 53.480 46.400 53.620 ;
        RECT 44.250 53.435 44.540 53.480 ;
        RECT 46.110 53.435 46.400 53.480 ;
        RECT 47.030 53.620 47.320 53.665 ;
        RECT 48.830 53.620 49.150 53.680 ;
        RECT 50.290 53.620 50.580 53.665 ;
        RECT 52.295 53.620 52.585 53.665 ;
        RECT 55.360 53.620 55.500 53.775 ;
        RECT 56.650 53.760 56.970 53.820 ;
        RECT 96.210 53.760 96.530 54.020 ;
        RECT 98.970 53.960 99.290 54.020 ;
        RECT 99.905 53.960 100.195 54.005 ;
        RECT 98.970 53.820 100.195 53.960 ;
        RECT 98.970 53.760 99.290 53.820 ;
        RECT 99.905 53.775 100.195 53.820 ;
        RECT 103.110 53.960 103.430 54.020 ;
        RECT 105.425 53.960 105.715 54.005 ;
        RECT 103.110 53.820 105.715 53.960 ;
        RECT 103.110 53.760 103.430 53.820 ;
        RECT 105.425 53.775 105.715 53.820 ;
        RECT 47.030 53.480 50.580 53.620 ;
        RECT 47.030 53.435 47.320 53.480 ;
        RECT 10.205 53.280 10.495 53.325 ;
        RECT 5.130 53.140 10.495 53.280 ;
        RECT 5.130 53.080 5.450 53.140 ;
        RECT 10.205 53.095 10.495 53.140 ;
        RECT 12.505 53.095 12.795 53.325 ;
        RECT 16.185 53.280 16.475 53.325 ;
        RECT 18.025 53.280 18.315 53.325 ;
        RECT 16.185 53.140 18.315 53.280 ;
        RECT 16.185 53.095 16.475 53.140 ;
        RECT 18.025 53.095 18.315 53.140 ;
        RECT 18.470 53.080 18.790 53.340 ;
        RECT 21.230 53.080 21.550 53.340 ;
        RECT 21.710 53.280 22.000 53.325 ;
        RECT 23.545 53.280 23.835 53.325 ;
        RECT 27.125 53.280 27.415 53.325 ;
        RECT 21.710 53.140 27.415 53.280 ;
        RECT 21.710 53.095 22.000 53.140 ;
        RECT 23.545 53.095 23.835 53.140 ;
        RECT 27.125 53.095 27.415 53.140 ;
        RECT 28.205 53.120 28.495 53.435 ;
        RECT 36.885 53.280 37.175 53.325 ;
        RECT 39.645 53.280 39.935 53.325 ;
        RECT 41.930 53.280 42.250 53.340 ;
        RECT 43.325 53.280 43.615 53.325 ;
        RECT 36.885 53.140 38.020 53.280 ;
        RECT 36.885 53.095 37.175 53.140 ;
        RECT 13.425 52.940 13.715 52.985 ;
        RECT 15.710 52.940 16.030 53.000 ;
        RECT 13.425 52.800 16.030 52.940 ;
        RECT 13.425 52.755 13.715 52.800 ;
        RECT 15.710 52.740 16.030 52.800 ;
        RECT 17.565 52.940 17.855 52.985 ;
        RECT 20.310 52.940 20.630 53.000 ;
        RECT 17.565 52.800 20.630 52.940 ;
        RECT 17.565 52.755 17.855 52.800 ;
        RECT 20.310 52.740 20.630 52.800 ;
        RECT 22.625 52.940 22.915 52.985 ;
        RECT 23.070 52.940 23.390 53.000 ;
        RECT 22.625 52.800 23.390 52.940 ;
        RECT 22.625 52.755 22.915 52.800 ;
        RECT 23.070 52.740 23.390 52.800 ;
        RECT 37.880 52.645 38.020 53.140 ;
        RECT 39.645 53.140 41.700 53.280 ;
        RECT 39.645 53.095 39.935 53.140 ;
        RECT 40.105 52.755 40.395 52.985 ;
        RECT 22.115 52.600 22.405 52.645 ;
        RECT 24.005 52.600 24.295 52.645 ;
        RECT 27.125 52.600 27.415 52.645 ;
        RECT 22.115 52.460 27.415 52.600 ;
        RECT 22.115 52.415 22.405 52.460 ;
        RECT 24.005 52.415 24.295 52.460 ;
        RECT 27.125 52.415 27.415 52.460 ;
        RECT 37.805 52.415 38.095 52.645 ;
        RECT 40.180 52.600 40.320 52.755 ;
        RECT 41.010 52.740 41.330 53.000 ;
        RECT 41.560 52.940 41.700 53.140 ;
        RECT 41.930 53.140 43.615 53.280 ;
        RECT 41.930 53.080 42.250 53.140 ;
        RECT 43.325 53.095 43.615 53.140 ;
        RECT 45.150 53.080 45.470 53.340 ;
        RECT 46.185 53.280 46.400 53.435 ;
        RECT 48.830 53.420 49.150 53.480 ;
        RECT 50.290 53.435 50.580 53.480 ;
        RECT 51.220 53.480 55.500 53.620 ;
        RECT 48.430 53.280 48.720 53.325 ;
        RECT 46.185 53.140 48.720 53.280 ;
        RECT 48.430 53.095 48.720 53.140 ;
        RECT 51.220 52.940 51.360 53.480 ;
        RECT 52.295 53.435 52.585 53.480 ;
        RECT 61.265 53.280 61.555 53.325 ;
        RECT 62.630 53.280 62.950 53.340 ;
        RECT 63.105 53.280 63.395 53.325 ;
        RECT 61.265 53.140 63.395 53.280 ;
        RECT 61.265 53.095 61.555 53.140 ;
        RECT 62.630 53.080 62.950 53.140 ;
        RECT 63.105 53.095 63.395 53.140 ;
        RECT 88.850 53.080 89.170 53.340 ;
        RECT 97.130 53.280 97.450 53.340 ;
        RECT 99.445 53.280 99.735 53.325 ;
        RECT 102.650 53.280 102.970 53.340 ;
        RECT 105.885 53.280 106.175 53.325 ;
        RECT 97.130 53.140 106.175 53.280 ;
        RECT 97.130 53.080 97.450 53.140 ;
        RECT 99.445 53.095 99.735 53.140 ;
        RECT 102.650 53.080 102.970 53.140 ;
        RECT 105.885 53.095 106.175 53.140 ;
        RECT 41.560 52.800 51.360 52.940 ;
        RECT 52.970 52.940 53.290 53.000 ;
        RECT 55.745 52.940 56.035 52.985 ;
        RECT 52.970 52.800 56.035 52.940 ;
        RECT 52.970 52.740 53.290 52.800 ;
        RECT 55.745 52.755 56.035 52.800 ;
        RECT 43.310 52.600 43.630 52.660 ;
        RECT 40.180 52.460 43.630 52.600 ;
        RECT 43.310 52.400 43.630 52.460 ;
        RECT 43.790 52.600 44.080 52.645 ;
        RECT 45.650 52.600 45.940 52.645 ;
        RECT 48.430 52.600 48.720 52.645 ;
        RECT 92.070 52.600 92.390 52.660 ;
        RECT 43.790 52.460 48.720 52.600 ;
        RECT 43.790 52.415 44.080 52.460 ;
        RECT 45.650 52.415 45.940 52.460 ;
        RECT 48.430 52.415 48.720 52.460 ;
        RECT 62.260 52.460 92.390 52.600 ;
        RECT 62.260 52.320 62.400 52.460 ;
        RECT 92.070 52.400 92.390 52.460 ;
        RECT 11.570 52.060 11.890 52.320 ;
        RECT 34.570 52.260 34.890 52.320 ;
        RECT 35.965 52.260 36.255 52.305 ;
        RECT 34.570 52.120 36.255 52.260 ;
        RECT 34.570 52.060 34.890 52.120 ;
        RECT 35.965 52.075 36.255 52.120 ;
        RECT 62.170 52.060 62.490 52.320 ;
        RECT 64.025 52.260 64.315 52.305 ;
        RECT 65.390 52.260 65.710 52.320 ;
        RECT 85.630 52.260 85.950 52.320 ;
        RECT 64.025 52.120 85.950 52.260 ;
        RECT 64.025 52.075 64.315 52.120 ;
        RECT 65.390 52.060 65.710 52.120 ;
        RECT 85.630 52.060 85.950 52.120 ;
        RECT 5.520 51.440 118.680 51.920 ;
        RECT 15.710 51.240 16.030 51.300 ;
        RECT 17.105 51.240 17.395 51.285 ;
        RECT 15.710 51.100 17.395 51.240 ;
        RECT 15.710 51.040 16.030 51.100 ;
        RECT 17.105 51.055 17.395 51.100 ;
        RECT 19.390 51.040 19.710 51.300 ;
        RECT 21.690 51.040 22.010 51.300 ;
        RECT 25.830 51.040 26.150 51.300 ;
        RECT 41.945 51.240 42.235 51.285 ;
        RECT 33.280 51.100 42.235 51.240 ;
        RECT 9.235 50.900 9.525 50.945 ;
        RECT 11.125 50.900 11.415 50.945 ;
        RECT 14.245 50.900 14.535 50.945 ;
        RECT 9.235 50.760 14.535 50.900 ;
        RECT 9.235 50.715 9.525 50.760 ;
        RECT 11.125 50.715 11.415 50.760 ;
        RECT 14.245 50.715 14.535 50.760 ;
        RECT 18.470 50.900 18.790 50.960 ;
        RECT 33.280 50.900 33.420 51.100 ;
        RECT 41.945 51.055 42.235 51.100 ;
        RECT 43.310 51.240 43.630 51.300 ;
        RECT 44.705 51.240 44.995 51.285 ;
        RECT 43.310 51.100 44.995 51.240 ;
        RECT 18.470 50.760 33.420 50.900 ;
        RECT 34.075 50.900 34.365 50.945 ;
        RECT 35.965 50.900 36.255 50.945 ;
        RECT 39.085 50.900 39.375 50.945 ;
        RECT 34.075 50.760 39.375 50.900 ;
        RECT 18.470 50.700 18.790 50.760 ;
        RECT 34.075 50.715 34.365 50.760 ;
        RECT 35.965 50.715 36.255 50.760 ;
        RECT 39.085 50.715 39.375 50.760 ;
        RECT 8.350 50.360 8.670 50.620 ;
        RECT 9.745 50.560 10.035 50.605 ;
        RECT 11.570 50.560 11.890 50.620 ;
        RECT 27.210 50.560 27.530 50.620 ;
        RECT 33.205 50.560 33.495 50.605 ;
        RECT 9.745 50.420 11.890 50.560 ;
        RECT 9.745 50.375 10.035 50.420 ;
        RECT 11.570 50.360 11.890 50.420 ;
        RECT 19.940 50.420 25.600 50.560 ;
        RECT 19.940 50.265 20.080 50.420 ;
        RECT 8.830 50.220 9.120 50.265 ;
        RECT 10.665 50.220 10.955 50.265 ;
        RECT 14.245 50.220 14.535 50.265 ;
        RECT 8.830 50.080 14.535 50.220 ;
        RECT 8.830 50.035 9.120 50.080 ;
        RECT 10.665 50.035 10.955 50.080 ;
        RECT 14.245 50.035 14.535 50.080 ;
        RECT 12.025 49.880 12.675 49.925 ;
        RECT 14.790 49.880 15.110 49.940 ;
        RECT 15.325 49.925 15.615 50.240 ;
        RECT 19.865 50.035 20.155 50.265 ;
        RECT 15.325 49.880 15.915 49.925 ;
        RECT 12.025 49.740 15.915 49.880 ;
        RECT 12.025 49.695 12.675 49.740 ;
        RECT 14.790 49.680 15.110 49.740 ;
        RECT 15.625 49.695 15.915 49.740 ;
        RECT 13.870 49.540 14.190 49.600 ;
        RECT 19.940 49.540 20.080 50.035 ;
        RECT 23.070 50.020 23.390 50.280 ;
        RECT 23.530 50.020 23.850 50.280 ;
        RECT 25.460 50.265 25.600 50.420 ;
        RECT 27.210 50.420 33.495 50.560 ;
        RECT 27.210 50.360 27.530 50.420 ;
        RECT 33.205 50.375 33.495 50.420 ;
        RECT 34.570 50.360 34.890 50.620 ;
        RECT 42.020 50.560 42.160 51.055 ;
        RECT 43.310 51.040 43.630 51.100 ;
        RECT 44.705 51.055 44.995 51.100 ;
        RECT 80.570 51.240 80.890 51.300 ;
        RECT 81.505 51.240 81.795 51.285 ;
        RECT 80.570 51.100 81.795 51.240 ;
        RECT 80.570 51.040 80.890 51.100 ;
        RECT 81.505 51.055 81.795 51.100 ;
        RECT 85.185 51.240 85.475 51.285 ;
        RECT 87.010 51.240 87.330 51.300 ;
        RECT 85.185 51.100 87.330 51.240 ;
        RECT 85.185 51.055 85.475 51.100 ;
        RECT 87.010 51.040 87.330 51.100 ;
        RECT 88.865 51.240 89.155 51.285 ;
        RECT 91.610 51.240 91.930 51.300 ;
        RECT 88.865 51.100 91.930 51.240 ;
        RECT 88.865 51.055 89.155 51.100 ;
        RECT 91.610 51.040 91.930 51.100 ;
        RECT 95.305 51.240 95.595 51.285 ;
        RECT 97.590 51.240 97.910 51.300 ;
        RECT 95.305 51.100 97.910 51.240 ;
        RECT 95.305 51.055 95.595 51.100 ;
        RECT 97.590 51.040 97.910 51.100 ;
        RECT 83.330 50.900 83.650 50.960 ;
        RECT 79.740 50.760 83.650 50.900 ;
        RECT 47.465 50.560 47.755 50.605 ;
        RECT 42.020 50.420 47.755 50.560 ;
        RECT 47.465 50.375 47.755 50.420 ;
        RECT 79.740 50.280 79.880 50.760 ;
        RECT 83.330 50.700 83.650 50.760 ;
        RECT 97.130 50.560 97.450 50.620 ;
        RECT 80.200 50.420 84.020 50.560 ;
        RECT 24.005 50.035 24.295 50.265 ;
        RECT 24.925 50.035 25.215 50.265 ;
        RECT 25.385 50.220 25.675 50.265 ;
        RECT 33.670 50.220 33.960 50.265 ;
        RECT 35.505 50.220 35.795 50.265 ;
        RECT 39.085 50.220 39.375 50.265 ;
        RECT 25.385 50.080 33.420 50.220 ;
        RECT 25.385 50.035 25.675 50.080 ;
        RECT 22.610 49.880 22.930 49.940 ;
        RECT 24.080 49.880 24.220 50.035 ;
        RECT 22.610 49.740 24.220 49.880 ;
        RECT 25.000 49.880 25.140 50.035 ;
        RECT 26.750 49.880 27.070 49.940 ;
        RECT 25.000 49.740 27.070 49.880 ;
        RECT 22.610 49.680 22.930 49.740 ;
        RECT 26.750 49.680 27.070 49.740 ;
        RECT 13.870 49.400 20.080 49.540 ;
        RECT 33.280 49.540 33.420 50.080 ;
        RECT 33.670 50.080 39.375 50.220 ;
        RECT 33.670 50.035 33.960 50.080 ;
        RECT 35.505 50.035 35.795 50.080 ;
        RECT 39.085 50.035 39.375 50.080 ;
        RECT 40.165 49.925 40.455 50.240 ;
        RECT 43.325 50.035 43.615 50.265 ;
        RECT 50.685 50.220 50.975 50.265 ;
        RECT 64.010 50.220 64.330 50.280 ;
        RECT 50.685 50.080 64.330 50.220 ;
        RECT 50.685 50.035 50.975 50.080 ;
        RECT 36.865 49.880 37.515 49.925 ;
        RECT 40.165 49.880 40.755 49.925 ;
        RECT 42.865 49.880 43.155 49.925 ;
        RECT 36.865 49.740 43.155 49.880 ;
        RECT 36.865 49.695 37.515 49.740 ;
        RECT 40.465 49.695 40.755 49.740 ;
        RECT 42.865 49.695 43.155 49.740 ;
        RECT 43.400 49.880 43.540 50.035 ;
        RECT 64.010 50.020 64.330 50.080 ;
        RECT 71.385 50.035 71.675 50.265 ;
        RECT 71.845 50.220 72.135 50.265 ;
        RECT 72.290 50.220 72.610 50.280 ;
        RECT 71.845 50.080 72.610 50.220 ;
        RECT 71.845 50.035 72.135 50.080 ;
        RECT 49.305 49.880 49.595 49.925 ;
        RECT 43.400 49.740 49.595 49.880 ;
        RECT 71.460 49.880 71.600 50.035 ;
        RECT 72.290 50.020 72.610 50.080 ;
        RECT 78.270 50.020 78.590 50.280 ;
        RECT 79.190 50.020 79.510 50.280 ;
        RECT 79.650 50.020 79.970 50.280 ;
        RECT 80.200 50.265 80.340 50.420 ;
        RECT 83.880 50.280 84.020 50.420 ;
        RECT 86.640 50.420 97.450 50.560 ;
        RECT 80.125 50.035 80.415 50.265 ;
        RECT 81.950 50.020 82.270 50.280 ;
        RECT 82.885 50.035 83.175 50.265 ;
        RECT 75.970 49.880 76.290 49.940 ;
        RECT 71.460 49.740 76.290 49.880 ;
        RECT 41.930 49.540 42.250 49.600 ;
        RECT 43.400 49.540 43.540 49.740 ;
        RECT 49.305 49.695 49.595 49.740 ;
        RECT 75.970 49.680 76.290 49.740 ;
        RECT 33.280 49.400 43.540 49.540 ;
        RECT 68.150 49.540 68.470 49.600 ;
        RECT 70.465 49.540 70.755 49.585 ;
        RECT 68.150 49.400 70.755 49.540 ;
        RECT 13.870 49.340 14.190 49.400 ;
        RECT 41.930 49.340 42.250 49.400 ;
        RECT 68.150 49.340 68.470 49.400 ;
        RECT 70.465 49.355 70.755 49.400 ;
        RECT 71.830 49.540 72.150 49.600 ;
        RECT 72.305 49.540 72.595 49.585 ;
        RECT 71.830 49.400 72.595 49.540 ;
        RECT 71.830 49.340 72.150 49.400 ;
        RECT 72.305 49.355 72.595 49.400 ;
        RECT 78.270 49.540 78.590 49.600 ;
        RECT 81.950 49.540 82.270 49.600 ;
        RECT 78.270 49.400 82.270 49.540 ;
        RECT 82.960 49.540 83.100 50.035 ;
        RECT 83.330 50.020 83.650 50.280 ;
        RECT 83.790 50.020 84.110 50.280 ;
        RECT 85.630 50.020 85.950 50.280 ;
        RECT 86.640 50.265 86.780 50.420 ;
        RECT 97.130 50.360 97.450 50.420 ;
        RECT 86.565 50.035 86.855 50.265 ;
        RECT 87.025 50.035 87.315 50.265 ;
        RECT 87.485 50.035 87.775 50.265 ;
        RECT 83.420 49.880 83.560 50.020 ;
        RECT 87.100 49.880 87.240 50.035 ;
        RECT 83.420 49.740 87.240 49.880 ;
        RECT 83.330 49.540 83.650 49.600 ;
        RECT 82.960 49.400 83.650 49.540 ;
        RECT 78.270 49.340 78.590 49.400 ;
        RECT 81.950 49.340 82.270 49.400 ;
        RECT 83.330 49.340 83.650 49.400 ;
        RECT 83.790 49.540 84.110 49.600 ;
        RECT 87.560 49.540 87.700 50.035 ;
        RECT 90.230 50.020 90.550 50.280 ;
        RECT 92.070 50.020 92.390 50.280 ;
        RECT 93.005 50.035 93.295 50.265 ;
        RECT 93.080 49.880 93.220 50.035 ;
        RECT 93.450 50.020 93.770 50.280 ;
        RECT 93.925 50.220 94.215 50.265 ;
        RECT 94.830 50.220 95.150 50.280 ;
        RECT 93.925 50.080 95.150 50.220 ;
        RECT 93.925 50.035 94.215 50.080 ;
        RECT 94.830 50.020 95.150 50.080 ;
        RECT 95.750 49.880 96.070 49.940 ;
        RECT 93.080 49.740 96.070 49.880 ;
        RECT 95.750 49.680 96.070 49.740 ;
        RECT 88.390 49.540 88.710 49.600 ;
        RECT 83.790 49.400 88.710 49.540 ;
        RECT 83.790 49.340 84.110 49.400 ;
        RECT 88.390 49.340 88.710 49.400 ;
        RECT 91.165 49.540 91.455 49.585 ;
        RECT 97.590 49.540 97.910 49.600 ;
        RECT 91.165 49.400 97.910 49.540 ;
        RECT 91.165 49.355 91.455 49.400 ;
        RECT 97.590 49.340 97.910 49.400 ;
        RECT 5.520 48.720 118.680 49.200 ;
        RECT 14.790 48.520 15.110 48.580 ;
        RECT 14.420 48.380 15.110 48.520 ;
        RECT 14.420 48.225 14.560 48.380 ;
        RECT 14.790 48.320 15.110 48.380 ;
        RECT 23.070 48.520 23.390 48.580 ;
        RECT 34.570 48.520 34.890 48.580 ;
        RECT 62.170 48.520 62.490 48.580 ;
        RECT 69.990 48.520 70.310 48.580 ;
        RECT 23.070 48.380 24.220 48.520 ;
        RECT 23.070 48.320 23.390 48.380 ;
        RECT 14.345 47.995 14.635 48.225 ;
        RECT 13.870 47.840 14.190 47.900 ;
        RECT 14.805 47.840 15.095 47.885 ;
        RECT 13.870 47.700 15.095 47.840 ;
        RECT 13.870 47.640 14.190 47.700 ;
        RECT 14.805 47.655 15.095 47.700 ;
        RECT 22.165 47.840 22.455 47.885 ;
        RECT 22.165 47.700 22.840 47.840 ;
        RECT 22.165 47.655 22.455 47.700 ;
        RECT 22.700 46.820 22.840 47.700 ;
        RECT 23.070 47.640 23.390 47.900 ;
        RECT 23.530 47.640 23.850 47.900 ;
        RECT 24.080 47.885 24.220 48.380 ;
        RECT 34.570 48.380 62.490 48.520 ;
        RECT 34.570 48.320 34.890 48.380 ;
        RECT 62.170 48.320 62.490 48.380 ;
        RECT 67.780 48.380 70.310 48.520 ;
        RECT 25.385 48.180 25.675 48.225 ;
        RECT 28.590 48.180 28.910 48.240 ;
        RECT 25.385 48.040 28.910 48.180 ;
        RECT 25.385 47.995 25.675 48.040 ;
        RECT 28.590 47.980 28.910 48.040 ;
        RECT 51.130 48.180 51.450 48.240 ;
        RECT 52.065 48.180 52.355 48.225 ;
        RECT 67.780 48.180 67.920 48.380 ;
        RECT 69.990 48.320 70.310 48.380 ;
        RECT 75.970 48.320 76.290 48.580 ;
        RECT 85.260 48.380 89.080 48.520 ;
        RECT 85.260 48.240 85.400 48.380 ;
        RECT 51.130 48.040 52.355 48.180 ;
        RECT 51.130 47.980 51.450 48.040 ;
        RECT 52.065 47.995 52.355 48.040 ;
        RECT 63.640 48.040 67.920 48.180 ;
        RECT 24.005 47.840 24.295 47.885 ;
        RECT 27.210 47.840 27.530 47.900 ;
        RECT 24.005 47.700 27.530 47.840 ;
        RECT 24.005 47.655 24.295 47.700 ;
        RECT 27.210 47.640 27.530 47.700 ;
        RECT 27.685 47.655 27.975 47.885 ;
        RECT 23.620 47.500 23.760 47.640 ;
        RECT 26.290 47.500 26.610 47.560 ;
        RECT 27.760 47.500 27.900 47.655 ;
        RECT 28.130 47.640 28.450 47.900 ;
        RECT 29.065 47.840 29.355 47.885 ;
        RECT 34.570 47.840 34.890 47.900 ;
        RECT 29.065 47.700 34.890 47.840 ;
        RECT 29.065 47.655 29.355 47.700 ;
        RECT 23.620 47.360 27.900 47.500 ;
        RECT 26.290 47.300 26.610 47.360 ;
        RECT 23.990 47.160 24.310 47.220 ;
        RECT 25.845 47.160 26.135 47.205 ;
        RECT 23.990 47.020 26.135 47.160 ;
        RECT 23.990 46.960 24.310 47.020 ;
        RECT 25.845 46.975 26.135 47.020 ;
        RECT 24.910 46.820 25.230 46.880 ;
        RECT 26.750 46.820 27.070 46.880 ;
        RECT 29.140 46.820 29.280 47.655 ;
        RECT 34.570 47.640 34.890 47.700 ;
        RECT 48.830 47.640 49.150 47.900 ;
        RECT 49.765 47.655 50.055 47.885 ;
        RECT 50.225 47.655 50.515 47.885 ;
        RECT 50.685 47.840 50.975 47.885 ;
        RECT 54.810 47.840 55.130 47.900 ;
        RECT 50.685 47.700 55.130 47.840 ;
        RECT 50.685 47.655 50.975 47.700 ;
        RECT 45.610 47.500 45.930 47.560 ;
        RECT 49.840 47.500 49.980 47.655 ;
        RECT 45.610 47.360 49.980 47.500 ;
        RECT 50.300 47.500 50.440 47.655 ;
        RECT 54.810 47.640 55.130 47.700 ;
        RECT 60.330 47.640 60.650 47.900 ;
        RECT 50.300 47.360 51.360 47.500 ;
        RECT 45.610 47.300 45.930 47.360 ;
        RECT 51.220 46.880 51.360 47.360 ;
        RECT 63.090 47.300 63.410 47.560 ;
        RECT 56.650 47.160 56.970 47.220 ;
        RECT 61.265 47.160 61.555 47.205 ;
        RECT 63.640 47.160 63.780 48.040 ;
        RECT 68.150 47.980 68.470 48.240 ;
        RECT 70.445 48.180 71.095 48.225 ;
        RECT 71.830 48.180 72.150 48.240 ;
        RECT 74.045 48.180 74.335 48.225 ;
        RECT 79.650 48.180 79.970 48.240 ;
        RECT 85.170 48.180 85.490 48.240 ;
        RECT 70.445 48.040 74.335 48.180 ;
        RECT 70.445 47.995 71.095 48.040 ;
        RECT 71.830 47.980 72.150 48.040 ;
        RECT 73.745 47.995 74.335 48.040 ;
        RECT 74.680 48.040 85.490 48.180 ;
        RECT 64.010 47.840 64.330 47.900 ;
        RECT 64.485 47.840 64.775 47.885 ;
        RECT 64.010 47.700 64.775 47.840 ;
        RECT 64.010 47.640 64.330 47.700 ;
        RECT 64.485 47.655 64.775 47.700 ;
        RECT 67.250 47.840 67.540 47.885 ;
        RECT 69.085 47.840 69.375 47.885 ;
        RECT 72.665 47.840 72.955 47.885 ;
        RECT 67.250 47.700 72.955 47.840 ;
        RECT 67.250 47.655 67.540 47.700 ;
        RECT 69.085 47.655 69.375 47.700 ;
        RECT 72.665 47.655 72.955 47.700 ;
        RECT 73.745 47.680 74.035 47.995 ;
        RECT 66.770 47.300 67.090 47.560 ;
        RECT 68.150 47.500 68.470 47.560 ;
        RECT 74.680 47.500 74.820 48.040 ;
        RECT 79.650 47.980 79.970 48.040 ;
        RECT 85.170 47.980 85.490 48.040 ;
        RECT 87.025 48.180 87.315 48.225 ;
        RECT 87.470 48.180 87.790 48.240 ;
        RECT 87.025 48.040 87.790 48.180 ;
        RECT 87.025 47.995 87.315 48.040 ;
        RECT 87.470 47.980 87.790 48.040 ;
        RECT 88.940 47.900 89.080 48.380 ;
        RECT 93.540 48.380 96.440 48.520 ;
        RECT 93.540 48.240 93.680 48.380 ;
        RECT 91.150 48.180 91.470 48.240 ;
        RECT 93.450 48.180 93.770 48.240 ;
        RECT 91.150 48.040 93.770 48.180 ;
        RECT 91.150 47.980 91.470 48.040 ;
        RECT 76.430 47.840 76.750 47.900 ;
        RECT 77.825 47.840 78.115 47.885 ;
        RECT 76.430 47.700 78.115 47.840 ;
        RECT 76.430 47.640 76.750 47.700 ;
        RECT 77.825 47.655 78.115 47.700 ;
        RECT 78.285 47.840 78.575 47.885 ;
        RECT 83.345 47.840 83.635 47.885 ;
        RECT 78.285 47.700 83.635 47.840 ;
        RECT 78.285 47.655 78.575 47.700 ;
        RECT 83.345 47.655 83.635 47.700 ;
        RECT 68.150 47.360 74.820 47.500 ;
        RECT 75.050 47.500 75.370 47.560 ;
        RECT 78.360 47.500 78.500 47.655 ;
        RECT 88.390 47.640 88.710 47.900 ;
        RECT 88.850 47.640 89.170 47.900 ;
        RECT 89.310 47.640 89.630 47.900 ;
        RECT 92.160 47.885 92.300 48.040 ;
        RECT 93.450 47.980 93.770 48.040 ;
        RECT 93.910 48.180 94.230 48.240 ;
        RECT 94.385 48.180 94.675 48.225 ;
        RECT 93.910 48.040 94.675 48.180 ;
        RECT 93.910 47.980 94.230 48.040 ;
        RECT 94.385 47.995 94.675 48.040 ;
        RECT 90.245 47.840 90.535 47.885 ;
        RECT 90.705 47.840 90.995 47.885 ;
        RECT 90.245 47.700 90.995 47.840 ;
        RECT 90.245 47.655 90.535 47.700 ;
        RECT 90.705 47.655 90.995 47.700 ;
        RECT 91.625 47.655 91.915 47.885 ;
        RECT 92.085 47.655 92.375 47.885 ;
        RECT 92.545 47.840 92.835 47.885 ;
        RECT 92.990 47.840 93.310 47.900 ;
        RECT 94.830 47.840 95.150 47.900 ;
        RECT 96.300 47.885 96.440 48.380 ;
        RECT 98.600 48.380 100.580 48.520 ;
        RECT 98.600 48.180 98.740 48.380 ;
        RECT 96.760 48.040 98.740 48.180 ;
        RECT 98.970 48.180 99.290 48.240 ;
        RECT 99.905 48.180 100.195 48.225 ;
        RECT 98.970 48.040 100.195 48.180 ;
        RECT 100.440 48.180 100.580 48.380 ;
        RECT 104.950 48.180 105.270 48.240 ;
        RECT 100.440 48.040 106.100 48.180 ;
        RECT 96.760 47.885 96.900 48.040 ;
        RECT 98.970 47.980 99.290 48.040 ;
        RECT 99.905 47.995 100.195 48.040 ;
        RECT 104.950 47.980 105.270 48.040 ;
        RECT 95.765 47.840 96.055 47.885 ;
        RECT 92.545 47.700 96.055 47.840 ;
        RECT 92.545 47.655 92.835 47.700 ;
        RECT 75.050 47.360 78.500 47.500 ;
        RECT 68.150 47.300 68.470 47.360 ;
        RECT 75.050 47.300 75.370 47.360 ;
        RECT 78.730 47.300 79.050 47.560 ;
        RECT 79.190 47.500 79.510 47.560 ;
        RECT 86.105 47.500 86.395 47.545 ;
        RECT 79.190 47.360 86.395 47.500 ;
        RECT 79.190 47.300 79.510 47.360 ;
        RECT 86.105 47.315 86.395 47.360 ;
        RECT 87.470 47.500 87.790 47.560 ;
        RECT 90.320 47.500 90.460 47.655 ;
        RECT 87.470 47.360 90.460 47.500 ;
        RECT 91.700 47.500 91.840 47.655 ;
        RECT 92.990 47.640 93.310 47.700 ;
        RECT 94.830 47.640 95.150 47.700 ;
        RECT 95.765 47.655 96.055 47.700 ;
        RECT 96.225 47.655 96.515 47.885 ;
        RECT 96.685 47.655 96.975 47.885 ;
        RECT 97.605 47.655 97.895 47.885 ;
        RECT 98.510 47.840 98.830 47.900 ;
        RECT 105.960 47.885 106.100 48.040 ;
        RECT 100.365 47.840 100.655 47.885 ;
        RECT 102.665 47.840 102.955 47.885 ;
        RECT 98.510 47.700 102.955 47.840 ;
        RECT 95.290 47.500 95.610 47.560 ;
        RECT 97.680 47.500 97.820 47.655 ;
        RECT 98.510 47.640 98.830 47.700 ;
        RECT 100.365 47.655 100.655 47.700 ;
        RECT 102.665 47.655 102.955 47.700 ;
        RECT 105.885 47.655 106.175 47.885 ;
        RECT 106.345 47.655 106.635 47.885 ;
        RECT 91.700 47.360 95.610 47.500 ;
        RECT 87.470 47.300 87.790 47.360 ;
        RECT 95.290 47.300 95.610 47.360 ;
        RECT 96.300 47.360 97.820 47.500 ;
        RECT 56.650 47.020 63.780 47.160 ;
        RECT 67.655 47.160 67.945 47.205 ;
        RECT 69.545 47.160 69.835 47.205 ;
        RECT 72.665 47.160 72.955 47.205 ;
        RECT 67.655 47.020 72.955 47.160 ;
        RECT 56.650 46.960 56.970 47.020 ;
        RECT 61.265 46.975 61.555 47.020 ;
        RECT 67.655 46.975 67.945 47.020 ;
        RECT 69.545 46.975 69.835 47.020 ;
        RECT 72.665 46.975 72.955 47.020 ;
        RECT 75.525 47.160 75.815 47.205 ;
        RECT 79.280 47.160 79.420 47.300 ;
        RECT 75.525 47.020 79.420 47.160 ;
        RECT 92.530 47.160 92.850 47.220 ;
        RECT 93.925 47.160 94.215 47.205 ;
        RECT 96.300 47.160 96.440 47.360 ;
        RECT 98.985 47.315 99.275 47.545 ;
        RECT 92.530 47.020 94.215 47.160 ;
        RECT 75.525 46.975 75.815 47.020 ;
        RECT 92.530 46.960 92.850 47.020 ;
        RECT 93.925 46.975 94.215 47.020 ;
        RECT 94.460 47.020 96.440 47.160 ;
        RECT 22.700 46.680 29.280 46.820 ;
        RECT 51.130 46.820 51.450 46.880 ;
        RECT 55.270 46.820 55.590 46.880 ;
        RECT 64.930 46.820 65.250 46.880 ;
        RECT 51.130 46.680 65.250 46.820 ;
        RECT 24.910 46.620 25.230 46.680 ;
        RECT 26.750 46.620 27.070 46.680 ;
        RECT 51.130 46.620 51.450 46.680 ;
        RECT 55.270 46.620 55.590 46.680 ;
        RECT 64.930 46.620 65.250 46.680 ;
        RECT 66.770 46.820 67.090 46.880 ;
        RECT 69.070 46.820 69.390 46.880 ;
        RECT 66.770 46.680 69.390 46.820 ;
        RECT 66.770 46.620 67.090 46.680 ;
        RECT 69.070 46.620 69.390 46.680 ;
        RECT 78.730 46.820 79.050 46.880 ;
        RECT 86.550 46.820 86.870 46.880 ;
        RECT 78.730 46.680 86.870 46.820 ;
        RECT 78.730 46.620 79.050 46.680 ;
        RECT 86.550 46.620 86.870 46.680 ;
        RECT 92.070 46.820 92.390 46.880 ;
        RECT 94.460 46.820 94.600 47.020 ;
        RECT 92.070 46.680 94.600 46.820 ;
        RECT 94.830 46.820 95.150 46.880 ;
        RECT 99.060 46.820 99.200 47.315 ;
        RECT 102.205 47.160 102.495 47.205 ;
        RECT 106.420 47.160 106.560 47.655 ;
        RECT 102.205 47.020 106.560 47.160 ;
        RECT 102.205 46.975 102.495 47.020 ;
        RECT 94.830 46.680 99.200 46.820 ;
        RECT 106.790 46.820 107.110 46.880 ;
        RECT 107.265 46.820 107.555 46.865 ;
        RECT 106.790 46.680 107.555 46.820 ;
        RECT 92.070 46.620 92.390 46.680 ;
        RECT 94.830 46.620 95.150 46.680 ;
        RECT 106.790 46.620 107.110 46.680 ;
        RECT 107.265 46.635 107.555 46.680 ;
        RECT 5.520 46.000 118.680 46.480 ;
        RECT 28.145 45.800 28.435 45.845 ;
        RECT 30.890 45.800 31.210 45.860 ;
        RECT 28.145 45.660 31.210 45.800 ;
        RECT 28.145 45.615 28.435 45.660 ;
        RECT 30.890 45.600 31.210 45.660 ;
        RECT 31.365 45.800 31.655 45.845 ;
        RECT 32.270 45.800 32.590 45.860 ;
        RECT 31.365 45.660 32.590 45.800 ;
        RECT 31.365 45.615 31.655 45.660 ;
        RECT 32.270 45.600 32.590 45.660 ;
        RECT 58.030 45.800 58.350 45.860 ;
        RECT 64.010 45.800 64.330 45.860 ;
        RECT 58.030 45.660 64.330 45.800 ;
        RECT 58.030 45.600 58.350 45.660 ;
        RECT 64.010 45.600 64.330 45.660 ;
        RECT 64.930 45.800 65.250 45.860 ;
        RECT 68.150 45.800 68.470 45.860 ;
        RECT 79.665 45.800 79.955 45.845 ;
        RECT 64.930 45.660 68.470 45.800 ;
        RECT 64.930 45.600 65.250 45.660 ;
        RECT 68.150 45.600 68.470 45.660 ;
        RECT 68.700 45.660 79.955 45.800 ;
        RECT 62.645 45.460 62.935 45.505 ;
        RECT 67.690 45.460 68.010 45.520 ;
        RECT 48.230 45.320 68.010 45.460 ;
        RECT 22.150 44.920 22.470 45.180 ;
        RECT 27.210 45.120 27.530 45.180 ;
        RECT 48.230 45.120 48.370 45.320 ;
        RECT 62.645 45.275 62.935 45.320 ;
        RECT 67.690 45.260 68.010 45.320 ;
        RECT 26.840 44.980 48.370 45.120 ;
        RECT 52.510 45.120 52.830 45.180 ;
        RECT 53.445 45.120 53.735 45.165 ;
        RECT 52.510 44.980 53.735 45.120 ;
        RECT 16.170 44.580 16.490 44.840 ;
        RECT 23.530 44.780 23.850 44.840 ;
        RECT 24.910 44.780 25.230 44.840 ;
        RECT 23.530 44.640 25.230 44.780 ;
        RECT 23.530 44.580 23.850 44.640 ;
        RECT 24.910 44.580 25.230 44.640 ;
        RECT 25.845 44.595 26.135 44.825 ;
        RECT 11.110 44.440 11.430 44.500 ;
        RECT 23.990 44.440 24.310 44.500 ;
        RECT 25.920 44.440 26.060 44.595 ;
        RECT 26.290 44.580 26.610 44.840 ;
        RECT 26.840 44.825 26.980 44.980 ;
        RECT 27.210 44.920 27.530 44.980 ;
        RECT 26.765 44.595 27.055 44.825 ;
        RECT 29.985 44.780 30.275 44.825 ;
        RECT 30.890 44.780 31.210 44.840 ;
        RECT 32.820 44.825 32.960 44.980 ;
        RECT 52.510 44.920 52.830 44.980 ;
        RECT 53.445 44.935 53.735 44.980 ;
        RECT 53.890 45.120 54.210 45.180 ;
        RECT 53.890 44.980 55.960 45.120 ;
        RECT 53.890 44.920 54.210 44.980 ;
        RECT 29.985 44.640 31.210 44.780 ;
        RECT 29.985 44.595 30.275 44.640 ;
        RECT 30.890 44.580 31.210 44.640 ;
        RECT 32.745 44.595 33.035 44.825 ;
        RECT 33.205 44.595 33.495 44.825 ;
        RECT 11.110 44.300 19.160 44.440 ;
        RECT 11.110 44.240 11.430 44.300 ;
        RECT 14.330 44.100 14.650 44.160 ;
        RECT 19.020 44.145 19.160 44.300 ;
        RECT 23.990 44.300 26.060 44.440 ;
        RECT 26.380 44.440 26.520 44.580 ;
        RECT 33.280 44.440 33.420 44.595 ;
        RECT 33.650 44.580 33.970 44.840 ;
        RECT 34.570 44.580 34.890 44.840 ;
        RECT 43.770 44.780 44.090 44.840 ;
        RECT 47.465 44.780 47.755 44.825 ;
        RECT 43.770 44.640 47.755 44.780 ;
        RECT 43.770 44.580 44.090 44.640 ;
        RECT 47.465 44.595 47.755 44.640 ;
        RECT 48.830 44.780 49.150 44.840 ;
        RECT 49.765 44.780 50.055 44.825 ;
        RECT 50.210 44.780 50.530 44.840 ;
        RECT 48.830 44.640 50.530 44.780 ;
        RECT 48.830 44.580 49.150 44.640 ;
        RECT 49.765 44.595 50.055 44.640 ;
        RECT 50.210 44.580 50.530 44.640 ;
        RECT 50.685 44.595 50.975 44.825 ;
        RECT 46.990 44.440 47.310 44.500 ;
        RECT 50.760 44.440 50.900 44.595 ;
        RECT 51.130 44.580 51.450 44.840 ;
        RECT 51.605 44.595 51.895 44.825 ;
        RECT 54.810 44.780 55.130 44.840 ;
        RECT 52.600 44.640 55.130 44.780 ;
        RECT 26.380 44.300 45.380 44.440 ;
        RECT 23.990 44.240 24.310 44.300 ;
        RECT 15.265 44.100 15.555 44.145 ;
        RECT 14.330 43.960 15.555 44.100 ;
        RECT 14.330 43.900 14.650 43.960 ;
        RECT 15.265 43.915 15.555 43.960 ;
        RECT 18.945 43.915 19.235 44.145 ;
        RECT 20.770 43.900 21.090 44.160 ;
        RECT 21.230 43.900 21.550 44.160 ;
        RECT 30.905 44.100 31.195 44.145 ;
        RECT 33.190 44.100 33.510 44.160 ;
        RECT 30.905 43.960 33.510 44.100 ;
        RECT 30.905 43.915 31.195 43.960 ;
        RECT 33.190 43.900 33.510 43.960 ;
        RECT 42.390 44.100 42.710 44.160 ;
        RECT 44.705 44.100 44.995 44.145 ;
        RECT 42.390 43.960 44.995 44.100 ;
        RECT 45.240 44.100 45.380 44.300 ;
        RECT 46.990 44.300 50.900 44.440 ;
        RECT 51.680 44.440 51.820 44.595 ;
        RECT 52.600 44.440 52.740 44.640 ;
        RECT 54.810 44.580 55.130 44.640 ;
        RECT 55.270 44.580 55.590 44.840 ;
        RECT 55.820 44.825 55.960 44.980 ;
        RECT 57.660 44.980 61.020 45.120 ;
        RECT 55.745 44.595 56.035 44.825 ;
        RECT 56.650 44.580 56.970 44.840 ;
        RECT 57.660 44.825 57.800 44.980 ;
        RECT 57.585 44.595 57.875 44.825 ;
        RECT 58.030 44.580 58.350 44.840 ;
        RECT 58.950 44.580 59.270 44.840 ;
        RECT 59.425 44.780 59.715 44.825 ;
        RECT 60.330 44.780 60.650 44.840 ;
        RECT 59.425 44.640 60.650 44.780 ;
        RECT 60.880 44.780 61.020 44.980 ;
        RECT 61.690 44.780 61.980 44.825 ;
        RECT 63.550 44.780 63.870 44.840 ;
        RECT 60.880 44.640 63.870 44.780 ;
        RECT 59.425 44.595 59.715 44.640 ;
        RECT 60.330 44.580 60.650 44.640 ;
        RECT 61.690 44.595 61.980 44.640 ;
        RECT 63.550 44.580 63.870 44.640 ;
        RECT 64.010 44.580 64.330 44.840 ;
        RECT 68.700 44.825 68.840 45.660 ;
        RECT 79.665 45.615 79.955 45.660 ;
        RECT 82.870 45.800 83.190 45.860 ;
        RECT 83.345 45.800 83.635 45.845 ;
        RECT 82.870 45.660 83.635 45.800 ;
        RECT 82.870 45.600 83.190 45.660 ;
        RECT 83.345 45.615 83.635 45.660 ;
        RECT 90.230 45.800 90.550 45.860 ;
        RECT 91.625 45.800 91.915 45.845 ;
        RECT 98.510 45.800 98.830 45.860 ;
        RECT 90.230 45.660 91.915 45.800 ;
        RECT 90.230 45.600 90.550 45.660 ;
        RECT 91.625 45.615 91.915 45.660 ;
        RECT 94.000 45.660 98.830 45.800 ;
        RECT 71.335 45.460 71.625 45.505 ;
        RECT 73.225 45.460 73.515 45.505 ;
        RECT 76.345 45.460 76.635 45.505 ;
        RECT 71.335 45.320 76.635 45.460 ;
        RECT 71.335 45.275 71.625 45.320 ;
        RECT 73.225 45.275 73.515 45.320 ;
        RECT 76.345 45.275 76.635 45.320 ;
        RECT 81.950 45.460 82.270 45.520 ;
        RECT 81.950 45.320 86.780 45.460 ;
        RECT 81.950 45.260 82.270 45.320 ;
        RECT 69.070 45.120 69.390 45.180 ;
        RECT 70.465 45.120 70.755 45.165 ;
        RECT 73.670 45.120 73.990 45.180 ;
        RECT 69.070 44.980 73.990 45.120 ;
        RECT 69.070 44.920 69.390 44.980 ;
        RECT 70.465 44.935 70.755 44.980 ;
        RECT 73.670 44.920 73.990 44.980 ;
        RECT 78.360 44.980 84.020 45.120 ;
        RECT 68.625 44.595 68.915 44.825 ;
        RECT 70.930 44.780 71.220 44.825 ;
        RECT 72.765 44.780 73.055 44.825 ;
        RECT 76.345 44.780 76.635 44.825 ;
        RECT 70.930 44.640 76.635 44.780 ;
        RECT 70.930 44.595 71.220 44.640 ;
        RECT 72.765 44.595 73.055 44.640 ;
        RECT 76.345 44.595 76.635 44.640 ;
        RECT 51.680 44.300 52.740 44.440 ;
        RECT 52.985 44.440 53.275 44.485 ;
        RECT 53.430 44.440 53.750 44.500 ;
        RECT 52.985 44.300 53.750 44.440 ;
        RECT 46.990 44.240 47.310 44.300 ;
        RECT 50.670 44.100 50.990 44.160 ;
        RECT 45.240 43.960 50.990 44.100 ;
        RECT 42.390 43.900 42.710 43.960 ;
        RECT 44.705 43.915 44.995 43.960 ;
        RECT 50.670 43.900 50.990 43.960 ;
        RECT 51.130 44.100 51.450 44.160 ;
        RECT 51.680 44.100 51.820 44.300 ;
        RECT 52.985 44.255 53.275 44.300 ;
        RECT 53.430 44.240 53.750 44.300 ;
        RECT 62.720 44.300 71.600 44.440 ;
        RECT 51.130 43.960 51.820 44.100 ;
        RECT 51.130 43.900 51.450 43.960 ;
        RECT 59.870 43.900 60.190 44.160 ;
        RECT 60.805 44.100 61.095 44.145 ;
        RECT 61.250 44.100 61.570 44.160 ;
        RECT 62.720 44.100 62.860 44.300 ;
        RECT 60.805 43.960 62.860 44.100 ;
        RECT 69.545 44.100 69.835 44.145 ;
        RECT 70.910 44.100 71.230 44.160 ;
        RECT 69.545 43.960 71.230 44.100 ;
        RECT 71.460 44.100 71.600 44.300 ;
        RECT 71.830 44.240 72.150 44.500 ;
        RECT 74.125 44.440 74.775 44.485 ;
        RECT 76.890 44.440 77.210 44.500 ;
        RECT 77.425 44.485 77.715 44.800 ;
        RECT 77.425 44.440 78.015 44.485 ;
        RECT 74.125 44.300 78.015 44.440 ;
        RECT 74.125 44.255 74.775 44.300 ;
        RECT 76.890 44.240 77.210 44.300 ;
        RECT 77.725 44.255 78.015 44.300 ;
        RECT 78.360 44.100 78.500 44.980 ;
        RECT 83.880 44.840 84.020 44.980 ;
        RECT 82.410 44.580 82.730 44.840 ;
        RECT 83.790 44.780 84.110 44.840 ;
        RECT 84.725 44.780 85.015 44.825 ;
        RECT 83.790 44.640 85.015 44.780 ;
        RECT 83.790 44.580 84.110 44.640 ;
        RECT 84.725 44.595 85.015 44.640 ;
        RECT 85.170 44.580 85.490 44.840 ;
        RECT 86.640 44.825 86.780 45.320 ;
        RECT 94.000 45.165 94.140 45.660 ;
        RECT 98.510 45.600 98.830 45.660 ;
        RECT 104.950 45.600 105.270 45.860 ;
        RECT 97.095 45.460 97.385 45.505 ;
        RECT 98.985 45.460 99.275 45.505 ;
        RECT 102.105 45.460 102.395 45.505 ;
        RECT 97.095 45.320 102.395 45.460 ;
        RECT 97.095 45.275 97.385 45.320 ;
        RECT 98.985 45.275 99.275 45.320 ;
        RECT 102.105 45.275 102.395 45.320 ;
        RECT 93.925 44.935 94.215 45.165 ;
        RECT 94.830 44.920 95.150 45.180 ;
        RECT 96.210 44.920 96.530 45.180 ;
        RECT 97.590 44.920 97.910 45.180 ;
        RECT 102.650 45.120 102.970 45.180 ;
        RECT 102.650 44.980 106.560 45.120 ;
        RECT 102.650 44.920 102.970 44.980 ;
        RECT 85.645 44.595 85.935 44.825 ;
        RECT 86.565 44.780 86.855 44.825 ;
        RECT 87.470 44.780 87.790 44.840 ;
        RECT 86.565 44.640 87.790 44.780 ;
        RECT 86.565 44.595 86.855 44.640 ;
        RECT 80.570 44.440 80.890 44.500 ;
        RECT 85.720 44.440 85.860 44.595 ;
        RECT 87.470 44.580 87.790 44.640 ;
        RECT 89.310 44.780 89.630 44.840 ;
        RECT 106.420 44.825 106.560 44.980 ;
        RECT 89.785 44.780 90.075 44.825 ;
        RECT 89.310 44.640 90.075 44.780 ;
        RECT 89.310 44.580 89.630 44.640 ;
        RECT 89.785 44.595 90.075 44.640 ;
        RECT 96.690 44.780 96.980 44.825 ;
        RECT 98.525 44.780 98.815 44.825 ;
        RECT 102.105 44.780 102.395 44.825 ;
        RECT 96.690 44.640 102.395 44.780 ;
        RECT 96.690 44.595 96.980 44.640 ;
        RECT 98.525 44.595 98.815 44.640 ;
        RECT 102.105 44.595 102.395 44.640 ;
        RECT 89.860 44.440 90.000 44.595 ;
        RECT 103.185 44.485 103.475 44.800 ;
        RECT 106.345 44.780 106.635 44.825 ;
        RECT 106.805 44.780 107.095 44.825 ;
        RECT 106.345 44.640 107.095 44.780 ;
        RECT 106.345 44.595 106.635 44.640 ;
        RECT 106.805 44.595 107.095 44.640 ;
        RECT 80.570 44.300 85.860 44.440 ;
        RECT 86.640 44.300 90.000 44.440 ;
        RECT 99.885 44.440 100.535 44.485 ;
        RECT 103.185 44.440 103.775 44.485 ;
        RECT 105.885 44.440 106.175 44.485 ;
        RECT 99.885 44.300 106.175 44.440 ;
        RECT 80.570 44.240 80.890 44.300 ;
        RECT 71.460 43.960 78.500 44.100 ;
        RECT 79.190 44.100 79.510 44.160 ;
        RECT 86.640 44.100 86.780 44.300 ;
        RECT 99.885 44.255 100.535 44.300 ;
        RECT 103.485 44.255 103.775 44.300 ;
        RECT 105.885 44.255 106.175 44.300 ;
        RECT 79.190 43.960 86.780 44.100 ;
        RECT 60.805 43.915 61.095 43.960 ;
        RECT 61.250 43.900 61.570 43.960 ;
        RECT 69.545 43.915 69.835 43.960 ;
        RECT 70.910 43.900 71.230 43.960 ;
        RECT 79.190 43.900 79.510 43.960 ;
        RECT 87.010 43.900 87.330 44.160 ;
        RECT 93.450 43.900 93.770 44.160 ;
        RECT 105.410 44.100 105.730 44.160 ;
        RECT 107.265 44.100 107.555 44.145 ;
        RECT 105.410 43.960 107.555 44.100 ;
        RECT 105.410 43.900 105.730 43.960 ;
        RECT 107.265 43.915 107.555 43.960 ;
        RECT 5.520 43.280 118.680 43.760 ;
        RECT 14.790 43.080 15.110 43.140 ;
        RECT 36.870 43.080 37.190 43.140 ;
        RECT 40.565 43.080 40.855 43.125 ;
        RECT 13.040 42.940 32.040 43.080 ;
        RECT 11.110 42.200 11.430 42.460 ;
        RECT 13.040 42.445 13.180 42.940 ;
        RECT 14.790 42.880 15.110 42.940 ;
        RECT 14.330 42.540 14.650 42.800 ;
        RECT 16.625 42.740 17.275 42.785 ;
        RECT 20.225 42.740 20.515 42.785 ;
        RECT 22.625 42.740 22.915 42.785 ;
        RECT 16.625 42.600 22.915 42.740 ;
        RECT 16.625 42.555 17.275 42.600 ;
        RECT 19.925 42.555 20.515 42.600 ;
        RECT 22.625 42.555 22.915 42.600 ;
        RECT 12.505 42.215 12.795 42.445 ;
        RECT 12.965 42.215 13.255 42.445 ;
        RECT 13.430 42.400 13.720 42.445 ;
        RECT 15.265 42.400 15.555 42.445 ;
        RECT 18.845 42.400 19.135 42.445 ;
        RECT 13.430 42.260 19.135 42.400 ;
        RECT 13.430 42.215 13.720 42.260 ;
        RECT 15.265 42.215 15.555 42.260 ;
        RECT 18.845 42.215 19.135 42.260 ;
        RECT 19.925 42.240 20.215 42.555 ;
        RECT 30.890 42.540 31.210 42.800 ;
        RECT 23.085 42.400 23.375 42.445 ;
        RECT 21.320 42.260 23.375 42.400 ;
        RECT 12.580 42.060 12.720 42.215 ;
        RECT 17.090 42.060 17.410 42.120 ;
        RECT 21.320 42.060 21.460 42.260 ;
        RECT 23.085 42.215 23.375 42.260 ;
        RECT 23.990 42.200 24.310 42.460 ;
        RECT 31.900 42.445 32.040 42.940 ;
        RECT 36.870 42.940 43.080 43.080 ;
        RECT 36.870 42.880 37.190 42.940 ;
        RECT 40.565 42.895 40.855 42.940 ;
        RECT 33.190 42.540 33.510 42.800 ;
        RECT 35.485 42.740 36.135 42.785 ;
        RECT 39.085 42.740 39.375 42.785 ;
        RECT 41.485 42.740 41.775 42.785 ;
        RECT 35.485 42.600 41.775 42.740 ;
        RECT 42.940 42.740 43.080 42.940 ;
        RECT 43.770 42.880 44.090 43.140 ;
        RECT 45.610 42.880 45.930 43.140 ;
        RECT 49.290 43.080 49.610 43.140 ;
        RECT 49.765 43.080 50.055 43.125 ;
        RECT 49.290 42.940 50.055 43.080 ;
        RECT 49.290 42.880 49.610 42.940 ;
        RECT 49.765 42.895 50.055 42.940 ;
        RECT 50.210 43.080 50.530 43.140 ;
        RECT 54.350 43.080 54.670 43.140 ;
        RECT 62.185 43.080 62.475 43.125 ;
        RECT 50.210 42.940 54.120 43.080 ;
        RECT 50.210 42.880 50.530 42.940 ;
        RECT 45.700 42.740 45.840 42.880 ;
        RECT 42.940 42.600 45.840 42.740 ;
        RECT 46.085 42.740 46.375 42.785 ;
        RECT 46.530 42.740 46.850 42.800 ;
        RECT 53.445 42.740 53.735 42.785 ;
        RECT 46.085 42.600 53.735 42.740 ;
        RECT 35.485 42.555 36.135 42.600 ;
        RECT 38.785 42.555 39.375 42.600 ;
        RECT 41.485 42.555 41.775 42.600 ;
        RECT 46.085 42.555 46.375 42.600 ;
        RECT 31.825 42.215 32.115 42.445 ;
        RECT 32.290 42.400 32.580 42.445 ;
        RECT 34.125 42.400 34.415 42.445 ;
        RECT 37.705 42.400 37.995 42.445 ;
        RECT 32.290 42.260 37.995 42.400 ;
        RECT 32.290 42.215 32.580 42.260 ;
        RECT 34.125 42.215 34.415 42.260 ;
        RECT 37.705 42.215 37.995 42.260 ;
        RECT 38.785 42.240 39.075 42.555 ;
        RECT 46.530 42.540 46.850 42.600 ;
        RECT 53.445 42.555 53.735 42.600 ;
        RECT 41.930 42.200 42.250 42.460 ;
        RECT 42.390 42.200 42.710 42.460 ;
        RECT 51.130 42.200 51.450 42.460 ;
        RECT 51.590 42.200 51.910 42.460 ;
        RECT 52.065 42.215 52.355 42.445 ;
        RECT 52.985 42.400 53.275 42.445 ;
        RECT 53.980 42.400 54.120 42.940 ;
        RECT 54.350 42.940 62.475 43.080 ;
        RECT 54.350 42.880 54.670 42.940 ;
        RECT 62.185 42.895 62.475 42.940 ;
        RECT 66.770 42.880 67.090 43.140 ;
        RECT 75.050 42.880 75.370 43.140 ;
        RECT 76.905 43.080 77.195 43.125 ;
        RECT 82.410 43.080 82.730 43.140 ;
        RECT 76.905 42.940 82.730 43.080 ;
        RECT 76.905 42.895 77.195 42.940 ;
        RECT 82.410 42.880 82.730 42.940 ;
        RECT 85.185 43.080 85.475 43.125 ;
        RECT 87.010 43.080 87.330 43.140 ;
        RECT 85.185 42.940 87.330 43.080 ;
        RECT 85.185 42.895 85.475 42.940 ;
        RECT 87.010 42.880 87.330 42.940 ;
        RECT 88.390 43.080 88.710 43.140 ;
        RECT 88.390 42.940 89.540 43.080 ;
        RECT 88.390 42.880 88.710 42.940 ;
        RECT 59.870 42.740 60.190 42.800 ;
        RECT 63.565 42.740 63.855 42.785 ;
        RECT 70.925 42.740 71.215 42.785 ;
        RECT 59.870 42.600 71.215 42.740 ;
        RECT 59.870 42.540 60.190 42.600 ;
        RECT 63.565 42.555 63.855 42.600 ;
        RECT 70.925 42.555 71.215 42.600 ;
        RECT 74.605 42.740 74.895 42.785 ;
        RECT 79.190 42.740 79.510 42.800 ;
        RECT 74.605 42.600 79.510 42.740 ;
        RECT 74.605 42.555 74.895 42.600 ;
        RECT 79.190 42.540 79.510 42.600 ;
        RECT 56.650 42.400 56.970 42.460 ;
        RECT 52.985 42.260 56.970 42.400 ;
        RECT 52.985 42.215 53.275 42.260 ;
        RECT 12.580 41.920 21.460 42.060 ;
        RECT 21.705 42.060 21.995 42.105 ;
        RECT 24.080 42.060 24.220 42.200 ;
        RECT 21.705 41.920 24.220 42.060 ;
        RECT 24.910 42.060 25.230 42.120 ;
        RECT 27.210 42.060 27.530 42.120 ;
        RECT 24.910 41.920 27.530 42.060 ;
        RECT 17.090 41.860 17.410 41.920 ;
        RECT 21.705 41.875 21.995 41.920 ;
        RECT 24.910 41.860 25.230 41.920 ;
        RECT 27.210 41.860 27.530 41.920 ;
        RECT 28.130 41.860 28.450 42.120 ;
        RECT 47.005 42.060 47.295 42.105 ;
        RECT 47.910 42.060 48.230 42.120 ;
        RECT 47.005 41.920 48.230 42.060 ;
        RECT 52.140 42.060 52.280 42.215 ;
        RECT 56.650 42.200 56.970 42.260 ;
        RECT 58.950 42.200 59.270 42.460 ;
        RECT 61.265 42.400 61.555 42.445 ;
        RECT 61.710 42.400 62.030 42.460 ;
        RECT 61.265 42.260 62.030 42.400 ;
        RECT 61.265 42.215 61.555 42.260 ;
        RECT 61.710 42.200 62.030 42.260 ;
        RECT 64.470 42.200 64.790 42.460 ;
        RECT 67.230 42.200 67.550 42.460 ;
        RECT 87.470 42.200 87.790 42.460 ;
        RECT 88.405 42.215 88.695 42.445 ;
        RECT 53.430 42.060 53.750 42.120 ;
        RECT 56.205 42.060 56.495 42.105 ;
        RECT 52.140 41.920 56.495 42.060 ;
        RECT 47.005 41.875 47.295 41.920 ;
        RECT 47.910 41.860 48.230 41.920 ;
        RECT 53.430 41.860 53.750 41.920 ;
        RECT 56.205 41.875 56.495 41.920 ;
        RECT 57.110 42.060 57.430 42.120 ;
        RECT 59.425 42.060 59.715 42.105 ;
        RECT 57.110 41.920 59.715 42.060 ;
        RECT 57.110 41.860 57.430 41.920 ;
        RECT 59.425 41.875 59.715 41.920 ;
        RECT 59.870 41.860 60.190 42.120 ;
        RECT 60.330 41.860 60.650 42.120 ;
        RECT 72.305 42.060 72.595 42.105 ;
        RECT 74.145 42.060 74.435 42.105 ;
        RECT 78.730 42.060 79.050 42.120 ;
        RECT 72.305 41.920 79.050 42.060 ;
        RECT 72.305 41.875 72.595 41.920 ;
        RECT 74.145 41.875 74.435 41.920 ;
        RECT 78.730 41.860 79.050 41.920 ;
        RECT 80.570 42.060 80.890 42.120 ;
        RECT 81.965 42.060 82.255 42.105 ;
        RECT 80.570 41.920 82.255 42.060 ;
        RECT 80.570 41.860 80.890 41.920 ;
        RECT 81.965 41.875 82.255 41.920 ;
        RECT 85.630 41.860 85.950 42.120 ;
        RECT 86.090 41.860 86.410 42.120 ;
        RECT 86.550 42.060 86.870 42.120 ;
        RECT 88.480 42.060 88.620 42.215 ;
        RECT 88.850 42.200 89.170 42.460 ;
        RECT 89.400 42.445 89.540 42.940 ;
        RECT 90.690 42.880 91.010 43.140 ;
        RECT 92.070 43.080 92.390 43.140 ;
        RECT 91.700 42.940 92.390 43.080 ;
        RECT 91.700 42.445 91.840 42.940 ;
        RECT 92.070 42.880 92.390 42.940 ;
        RECT 92.530 42.880 92.850 43.140 ;
        RECT 92.990 43.080 93.310 43.140 ;
        RECT 96.210 43.080 96.530 43.140 ;
        RECT 92.990 42.940 93.680 43.080 ;
        RECT 92.990 42.880 93.310 42.940 ;
        RECT 92.620 42.740 92.760 42.880 ;
        RECT 92.620 42.600 93.220 42.740 ;
        RECT 89.325 42.215 89.615 42.445 ;
        RECT 91.625 42.215 91.915 42.445 ;
        RECT 92.070 42.400 92.390 42.460 ;
        RECT 93.080 42.445 93.220 42.600 ;
        RECT 93.540 42.445 93.680 42.940 ;
        RECT 96.210 42.940 107.940 43.080 ;
        RECT 96.210 42.880 96.530 42.940 ;
        RECT 94.845 42.740 95.135 42.785 ;
        RECT 98.050 42.740 98.370 42.800 ;
        RECT 94.845 42.600 98.370 42.740 ;
        RECT 94.845 42.555 95.135 42.600 ;
        RECT 98.050 42.540 98.370 42.600 ;
        RECT 98.970 42.540 99.290 42.800 ;
        RECT 100.925 42.740 101.215 42.785 ;
        RECT 104.165 42.740 104.815 42.785 ;
        RECT 105.410 42.740 105.730 42.800 ;
        RECT 100.925 42.600 105.730 42.740 ;
        RECT 100.925 42.555 101.515 42.600 ;
        RECT 104.165 42.555 104.815 42.600 ;
        RECT 92.545 42.400 92.835 42.445 ;
        RECT 92.070 42.260 92.835 42.400 ;
        RECT 92.070 42.200 92.390 42.260 ;
        RECT 92.545 42.215 92.835 42.260 ;
        RECT 93.005 42.215 93.295 42.445 ;
        RECT 93.465 42.215 93.755 42.445 ;
        RECT 95.750 42.400 96.070 42.460 ;
        RECT 95.750 42.260 99.660 42.400 ;
        RECT 95.750 42.200 96.070 42.260 ;
        RECT 99.520 42.105 99.660 42.260 ;
        RECT 101.225 42.240 101.515 42.555 ;
        RECT 105.410 42.540 105.730 42.600 ;
        RECT 106.790 42.540 107.110 42.800 ;
        RECT 107.800 42.740 107.940 42.940 ;
        RECT 107.800 42.600 108.400 42.740 ;
        RECT 108.260 42.445 108.400 42.600 ;
        RECT 102.305 42.400 102.595 42.445 ;
        RECT 105.885 42.400 106.175 42.445 ;
        RECT 107.720 42.400 108.010 42.445 ;
        RECT 102.305 42.260 108.010 42.400 ;
        RECT 102.305 42.215 102.595 42.260 ;
        RECT 105.885 42.215 106.175 42.260 ;
        RECT 107.720 42.215 108.010 42.260 ;
        RECT 108.185 42.215 108.475 42.445 ;
        RECT 86.550 41.920 88.620 42.060 ;
        RECT 86.550 41.860 86.870 41.920 ;
        RECT 99.445 41.875 99.735 42.105 ;
        RECT 12.045 41.720 12.335 41.765 ;
        RECT 13.835 41.720 14.125 41.765 ;
        RECT 15.725 41.720 16.015 41.765 ;
        RECT 18.845 41.720 19.135 41.765 ;
        RECT 12.045 41.580 13.640 41.720 ;
        RECT 12.045 41.535 12.335 41.580 ;
        RECT 8.350 41.380 8.670 41.440 ;
        RECT 10.205 41.380 10.495 41.425 ;
        RECT 8.350 41.240 10.495 41.380 ;
        RECT 13.500 41.380 13.640 41.580 ;
        RECT 13.835 41.580 19.135 41.720 ;
        RECT 13.835 41.535 14.125 41.580 ;
        RECT 15.725 41.535 16.015 41.580 ;
        RECT 18.845 41.535 19.135 41.580 ;
        RECT 32.695 41.720 32.985 41.765 ;
        RECT 34.585 41.720 34.875 41.765 ;
        RECT 37.705 41.720 37.995 41.765 ;
        RECT 32.695 41.580 37.995 41.720 ;
        RECT 32.695 41.535 32.985 41.580 ;
        RECT 34.585 41.535 34.875 41.580 ;
        RECT 37.705 41.535 37.995 41.580 ;
        RECT 47.450 41.720 47.770 41.780 ;
        RECT 53.890 41.720 54.210 41.780 ;
        RECT 65.390 41.720 65.710 41.780 ;
        RECT 47.450 41.580 54.210 41.720 ;
        RECT 47.450 41.520 47.770 41.580 ;
        RECT 53.890 41.520 54.210 41.580 ;
        RECT 54.440 41.580 65.710 41.720 ;
        RECT 15.250 41.380 15.570 41.440 ;
        RECT 13.500 41.240 15.570 41.380 ;
        RECT 8.350 41.180 8.670 41.240 ;
        RECT 10.205 41.195 10.495 41.240 ;
        RECT 15.250 41.180 15.570 41.240 ;
        RECT 27.210 41.180 27.530 41.440 ;
        RECT 43.310 41.180 43.630 41.440 ;
        RECT 50.670 41.380 50.990 41.440 ;
        RECT 54.440 41.380 54.580 41.580 ;
        RECT 65.390 41.520 65.710 41.580 ;
        RECT 76.430 41.720 76.750 41.780 ;
        RECT 79.205 41.720 79.495 41.765 ;
        RECT 76.430 41.580 79.495 41.720 ;
        RECT 76.430 41.520 76.750 41.580 ;
        RECT 79.205 41.535 79.495 41.580 ;
        RECT 102.305 41.720 102.595 41.765 ;
        RECT 105.425 41.720 105.715 41.765 ;
        RECT 107.315 41.720 107.605 41.765 ;
        RECT 102.305 41.580 107.605 41.720 ;
        RECT 102.305 41.535 102.595 41.580 ;
        RECT 105.425 41.535 105.715 41.580 ;
        RECT 107.315 41.535 107.605 41.580 ;
        RECT 50.670 41.240 54.580 41.380 ;
        RECT 82.870 41.380 83.190 41.440 ;
        RECT 83.345 41.380 83.635 41.425 ;
        RECT 82.870 41.240 83.635 41.380 ;
        RECT 50.670 41.180 50.990 41.240 ;
        RECT 82.870 41.180 83.190 41.240 ;
        RECT 83.345 41.195 83.635 41.240 ;
        RECT 86.090 41.380 86.410 41.440 ;
        RECT 87.470 41.380 87.790 41.440 ;
        RECT 86.090 41.240 87.790 41.380 ;
        RECT 86.090 41.180 86.410 41.240 ;
        RECT 87.470 41.180 87.790 41.240 ;
        RECT 5.520 40.560 118.680 41.040 ;
        RECT 16.170 40.360 16.490 40.420 ;
        RECT 18.945 40.360 19.235 40.405 ;
        RECT 16.170 40.220 19.235 40.360 ;
        RECT 16.170 40.160 16.490 40.220 ;
        RECT 18.945 40.175 19.235 40.220 ;
        RECT 28.130 40.360 28.450 40.420 ;
        RECT 33.665 40.360 33.955 40.405 ;
        RECT 47.910 40.360 48.230 40.420 ;
        RECT 28.130 40.220 33.955 40.360 ;
        RECT 28.130 40.160 28.450 40.220 ;
        RECT 33.665 40.175 33.955 40.220 ;
        RECT 36.500 40.220 48.230 40.360 ;
        RECT 9.235 40.020 9.525 40.065 ;
        RECT 11.125 40.020 11.415 40.065 ;
        RECT 14.245 40.020 14.535 40.065 ;
        RECT 9.235 39.880 14.535 40.020 ;
        RECT 9.235 39.835 9.525 39.880 ;
        RECT 11.125 39.835 11.415 39.880 ;
        RECT 14.245 39.835 14.535 39.880 ;
        RECT 17.105 40.020 17.395 40.065 ;
        RECT 22.610 40.020 22.930 40.080 ;
        RECT 34.570 40.020 34.890 40.080 ;
        RECT 17.105 39.880 22.930 40.020 ;
        RECT 17.105 39.835 17.395 39.880 ;
        RECT 22.610 39.820 22.930 39.880 ;
        RECT 24.080 39.880 34.890 40.020 ;
        RECT 8.365 39.680 8.655 39.725 ;
        RECT 14.790 39.680 15.110 39.740 ;
        RECT 8.365 39.540 15.110 39.680 ;
        RECT 8.365 39.495 8.655 39.540 ;
        RECT 14.790 39.480 15.110 39.540 ;
        RECT 22.150 39.480 22.470 39.740 ;
        RECT 8.830 39.340 9.120 39.385 ;
        RECT 10.665 39.340 10.955 39.385 ;
        RECT 14.245 39.340 14.535 39.385 ;
        RECT 8.830 39.200 14.535 39.340 ;
        RECT 8.830 39.155 9.120 39.200 ;
        RECT 10.665 39.155 10.955 39.200 ;
        RECT 14.245 39.155 14.535 39.200 ;
        RECT 15.250 39.360 15.570 39.400 ;
        RECT 15.250 39.140 15.615 39.360 ;
        RECT 20.785 39.340 21.075 39.385 ;
        RECT 21.230 39.340 21.550 39.400 ;
        RECT 20.785 39.200 21.550 39.340 ;
        RECT 20.785 39.155 21.075 39.200 ;
        RECT 21.230 39.140 21.550 39.200 ;
        RECT 23.085 39.340 23.375 39.385 ;
        RECT 23.530 39.340 23.850 39.400 ;
        RECT 24.080 39.385 24.220 39.880 ;
        RECT 34.570 39.820 34.890 39.880 ;
        RECT 26.305 39.680 26.595 39.725 ;
        RECT 28.590 39.680 28.910 39.740 ;
        RECT 24.540 39.540 25.600 39.680 ;
        RECT 24.540 39.385 24.680 39.540 ;
        RECT 23.085 39.200 23.850 39.340 ;
        RECT 23.085 39.155 23.375 39.200 ;
        RECT 23.530 39.140 23.850 39.200 ;
        RECT 24.005 39.155 24.295 39.385 ;
        RECT 24.465 39.155 24.755 39.385 ;
        RECT 24.910 39.140 25.230 39.400 ;
        RECT 25.460 39.340 25.600 39.540 ;
        RECT 26.305 39.540 28.910 39.680 ;
        RECT 26.305 39.495 26.595 39.540 ;
        RECT 28.590 39.480 28.910 39.540 ;
        RECT 29.985 39.680 30.275 39.725 ;
        RECT 35.030 39.680 35.350 39.740 ;
        RECT 36.500 39.725 36.640 40.220 ;
        RECT 47.910 40.160 48.230 40.220 ;
        RECT 53.430 40.160 53.750 40.420 ;
        RECT 54.825 40.360 55.115 40.405 ;
        RECT 58.030 40.360 58.350 40.420 ;
        RECT 54.825 40.220 58.350 40.360 ;
        RECT 54.825 40.175 55.115 40.220 ;
        RECT 58.030 40.160 58.350 40.220 ;
        RECT 63.550 40.360 63.870 40.420 ;
        RECT 66.325 40.360 66.615 40.405 ;
        RECT 63.550 40.220 66.615 40.360 ;
        RECT 63.550 40.160 63.870 40.220 ;
        RECT 66.325 40.175 66.615 40.220 ;
        RECT 73.225 40.360 73.515 40.405 ;
        RECT 76.890 40.360 77.210 40.420 ;
        RECT 73.225 40.220 77.210 40.360 ;
        RECT 73.225 40.175 73.515 40.220 ;
        RECT 76.890 40.160 77.210 40.220 ;
        RECT 84.725 40.360 85.015 40.405 ;
        RECT 85.630 40.360 85.950 40.420 ;
        RECT 87.010 40.360 87.330 40.420 ;
        RECT 84.725 40.220 87.330 40.360 ;
        RECT 84.725 40.175 85.015 40.220 ;
        RECT 85.630 40.160 85.950 40.220 ;
        RECT 87.010 40.160 87.330 40.220 ;
        RECT 92.085 40.360 92.375 40.405 ;
        RECT 93.450 40.360 93.770 40.420 ;
        RECT 92.085 40.220 93.770 40.360 ;
        RECT 92.085 40.175 92.375 40.220 ;
        RECT 93.450 40.160 93.770 40.220 ;
        RECT 43.310 40.020 43.630 40.080 ;
        RECT 45.575 40.020 45.865 40.065 ;
        RECT 47.465 40.020 47.755 40.065 ;
        RECT 50.585 40.020 50.875 40.065 ;
        RECT 43.310 39.880 45.380 40.020 ;
        RECT 43.310 39.820 43.630 39.880 ;
        RECT 36.425 39.680 36.715 39.725 ;
        RECT 29.985 39.540 36.715 39.680 ;
        RECT 29.985 39.495 30.275 39.540 ;
        RECT 35.030 39.480 35.350 39.540 ;
        RECT 36.425 39.495 36.715 39.540 ;
        RECT 39.170 39.680 39.490 39.740 ;
        RECT 44.705 39.680 44.995 39.725 ;
        RECT 39.170 39.540 44.995 39.680 ;
        RECT 45.240 39.680 45.380 39.880 ;
        RECT 45.575 39.880 50.875 40.020 ;
        RECT 45.575 39.835 45.865 39.880 ;
        RECT 47.465 39.835 47.755 39.880 ;
        RECT 50.585 39.835 50.875 39.880 ;
        RECT 57.110 40.020 57.430 40.080 ;
        RECT 60.330 40.020 60.650 40.080 ;
        RECT 102.205 40.020 102.495 40.065 ;
        RECT 57.110 39.880 65.620 40.020 ;
        RECT 57.110 39.820 57.430 39.880 ;
        RECT 60.330 39.820 60.650 39.880 ;
        RECT 46.085 39.680 46.375 39.725 ;
        RECT 45.240 39.540 46.375 39.680 ;
        RECT 39.170 39.480 39.490 39.540 ;
        RECT 44.705 39.495 44.995 39.540 ;
        RECT 46.085 39.495 46.375 39.540 ;
        RECT 55.745 39.680 56.035 39.725 ;
        RECT 55.745 39.540 58.260 39.680 ;
        RECT 55.745 39.495 56.035 39.540 ;
        RECT 26.750 39.340 27.070 39.400 ;
        RECT 25.460 39.200 27.070 39.340 ;
        RECT 26.750 39.140 27.070 39.200 ;
        RECT 27.210 39.140 27.530 39.400 ;
        RECT 29.065 39.340 29.355 39.385 ;
        RECT 33.650 39.340 33.970 39.400 ;
        RECT 29.065 39.200 33.970 39.340 ;
        RECT 29.065 39.155 29.355 39.200 ;
        RECT 33.650 39.140 33.970 39.200 ;
        RECT 35.965 39.340 36.255 39.385 ;
        RECT 36.870 39.340 37.190 39.400 ;
        RECT 35.965 39.200 37.190 39.340 ;
        RECT 35.965 39.155 36.255 39.200 ;
        RECT 36.870 39.140 37.190 39.200 ;
        RECT 41.930 39.340 42.250 39.400 ;
        RECT 42.865 39.340 43.155 39.385 ;
        RECT 41.930 39.200 43.155 39.340 ;
        RECT 41.930 39.140 42.250 39.200 ;
        RECT 42.865 39.155 43.155 39.200 ;
        RECT 45.170 39.340 45.460 39.385 ;
        RECT 47.005 39.340 47.295 39.385 ;
        RECT 50.585 39.340 50.875 39.385 ;
        RECT 45.170 39.200 50.875 39.340 ;
        RECT 45.170 39.155 45.460 39.200 ;
        RECT 47.005 39.155 47.295 39.200 ;
        RECT 50.585 39.155 50.875 39.200 ;
        RECT 8.350 39.000 8.670 39.060 ;
        RECT 15.325 39.045 15.615 39.140 ;
        RECT 9.745 39.000 10.035 39.045 ;
        RECT 8.350 38.860 10.035 39.000 ;
        RECT 8.350 38.800 8.670 38.860 ;
        RECT 9.745 38.815 10.035 38.860 ;
        RECT 12.025 39.000 12.675 39.045 ;
        RECT 15.325 39.000 15.915 39.045 ;
        RECT 27.300 39.000 27.440 39.140 ;
        RECT 51.665 39.045 51.955 39.360 ;
        RECT 56.190 39.140 56.510 39.400 ;
        RECT 56.665 39.155 56.955 39.385 ;
        RECT 28.605 39.000 28.895 39.045 ;
        RECT 48.365 39.000 49.015 39.045 ;
        RECT 51.665 39.000 52.255 39.045 ;
        RECT 12.025 38.860 15.915 39.000 ;
        RECT 12.025 38.815 12.675 38.860 ;
        RECT 15.625 38.815 15.915 38.860 ;
        RECT 21.320 38.860 28.895 39.000 ;
        RECT 21.320 38.705 21.460 38.860 ;
        RECT 28.605 38.815 28.895 38.860 ;
        RECT 46.620 38.860 52.255 39.000 ;
        RECT 21.245 38.475 21.535 38.705 ;
        RECT 26.765 38.660 27.055 38.705 ;
        RECT 27.210 38.660 27.530 38.720 ;
        RECT 26.765 38.520 27.530 38.660 ;
        RECT 26.765 38.475 27.055 38.520 ;
        RECT 27.210 38.460 27.530 38.520 ;
        RECT 35.490 38.460 35.810 38.720 ;
        RECT 43.325 38.660 43.615 38.705 ;
        RECT 46.620 38.660 46.760 38.860 ;
        RECT 48.365 38.815 49.015 38.860 ;
        RECT 51.965 38.815 52.255 38.860 ;
        RECT 43.325 38.520 46.760 38.660 ;
        RECT 56.740 38.660 56.880 39.155 ;
        RECT 57.110 39.140 57.430 39.400 ;
        RECT 58.120 39.385 58.260 39.540 ;
        RECT 59.410 39.480 59.730 39.740 ;
        RECT 60.420 39.680 60.560 39.820 ;
        RECT 65.480 39.725 65.620 39.880 ;
        RECT 102.205 39.880 106.560 40.020 ;
        RECT 102.205 39.835 102.495 39.880 ;
        RECT 64.485 39.680 64.775 39.725 ;
        RECT 60.420 39.540 61.020 39.680 ;
        RECT 58.045 39.340 58.335 39.385 ;
        RECT 58.045 39.200 59.640 39.340 ;
        RECT 58.045 39.155 58.335 39.200 ;
        RECT 59.500 39.060 59.640 39.200 ;
        RECT 60.330 39.140 60.650 39.400 ;
        RECT 60.880 39.385 61.020 39.540 ;
        RECT 62.260 39.540 64.775 39.680 ;
        RECT 60.805 39.155 61.095 39.385 ;
        RECT 61.250 39.340 61.570 39.400 ;
        RECT 62.260 39.385 62.400 39.540 ;
        RECT 64.485 39.495 64.775 39.540 ;
        RECT 65.405 39.495 65.695 39.725 ;
        RECT 82.870 39.680 83.190 39.740 ;
        RECT 89.310 39.680 89.630 39.740 ;
        RECT 81.580 39.540 83.190 39.680 ;
        RECT 62.185 39.340 62.475 39.385 ;
        RECT 61.250 39.200 62.475 39.340 ;
        RECT 61.250 39.140 61.570 39.200 ;
        RECT 62.185 39.155 62.475 39.200 ;
        RECT 64.025 39.155 64.315 39.385 ;
        RECT 59.410 38.800 59.730 39.060 ;
        RECT 58.950 38.660 59.270 38.720 ;
        RECT 60.330 38.660 60.650 38.720 ;
        RECT 61.250 38.660 61.570 38.720 ;
        RECT 56.740 38.520 61.570 38.660 ;
        RECT 43.325 38.475 43.615 38.520 ;
        RECT 58.950 38.460 59.270 38.520 ;
        RECT 60.330 38.460 60.650 38.520 ;
        RECT 61.250 38.460 61.570 38.520 ;
        RECT 61.710 38.660 62.030 38.720 ;
        RECT 64.100 38.660 64.240 39.155 ;
        RECT 64.930 39.140 65.250 39.400 ;
        RECT 72.290 39.340 72.610 39.400 ;
        RECT 72.765 39.340 73.055 39.385 ;
        RECT 72.290 39.200 73.055 39.340 ;
        RECT 72.290 39.140 72.610 39.200 ;
        RECT 72.765 39.155 73.055 39.200 ;
        RECT 73.670 39.340 73.990 39.400 ;
        RECT 81.580 39.385 81.720 39.540 ;
        RECT 82.870 39.480 83.190 39.540 ;
        RECT 83.420 39.540 89.630 39.680 ;
        RECT 83.420 39.385 83.560 39.540 ;
        RECT 89.310 39.480 89.630 39.540 ;
        RECT 94.830 39.680 95.150 39.740 ;
        RECT 106.420 39.725 106.560 39.880 ;
        RECT 98.985 39.680 99.275 39.725 ;
        RECT 94.830 39.540 99.275 39.680 ;
        RECT 94.830 39.480 95.150 39.540 ;
        RECT 98.985 39.495 99.275 39.540 ;
        RECT 106.345 39.495 106.635 39.725 ;
        RECT 77.365 39.340 77.655 39.385 ;
        RECT 73.670 39.200 77.655 39.340 ;
        RECT 73.670 39.140 73.990 39.200 ;
        RECT 77.365 39.155 77.655 39.200 ;
        RECT 81.505 39.155 81.795 39.385 ;
        RECT 81.965 39.155 82.255 39.385 ;
        RECT 83.345 39.155 83.635 39.385 ;
        RECT 86.550 39.340 86.870 39.400 ;
        RECT 87.485 39.340 87.775 39.385 ;
        RECT 86.550 39.200 87.775 39.340 ;
        RECT 82.040 39.000 82.180 39.155 ;
        RECT 86.550 39.140 86.870 39.200 ;
        RECT 87.485 39.155 87.775 39.200 ;
        RECT 88.850 39.340 89.170 39.400 ;
        RECT 91.165 39.340 91.455 39.385 ;
        RECT 88.850 39.200 91.455 39.340 ;
        RECT 88.850 39.140 89.170 39.200 ;
        RECT 91.165 39.155 91.455 39.200 ;
        RECT 95.290 39.140 95.610 39.400 ;
        RECT 97.130 39.340 97.450 39.400 ;
        RECT 99.905 39.340 100.195 39.385 ;
        RECT 103.110 39.340 103.430 39.400 ;
        RECT 105.425 39.340 105.715 39.385 ;
        RECT 97.130 39.200 105.715 39.340 ;
        RECT 97.130 39.140 97.450 39.200 ;
        RECT 99.905 39.155 100.195 39.200 ;
        RECT 103.110 39.140 103.430 39.200 ;
        RECT 105.425 39.155 105.715 39.200 ;
        RECT 109.565 39.340 109.855 39.385 ;
        RECT 110.945 39.340 111.235 39.385 ;
        RECT 109.565 39.200 111.235 39.340 ;
        RECT 109.565 39.155 109.855 39.200 ;
        RECT 110.945 39.155 111.235 39.200 ;
        RECT 88.405 39.000 88.695 39.045 ;
        RECT 82.040 38.860 88.695 39.000 ;
        RECT 88.405 38.815 88.695 38.860 ;
        RECT 98.970 39.000 99.290 39.060 ;
        RECT 100.365 39.000 100.655 39.045 ;
        RECT 98.970 38.860 100.655 39.000 ;
        RECT 98.970 38.800 99.290 38.860 ;
        RECT 100.365 38.815 100.655 38.860 ;
        RECT 61.710 38.520 64.240 38.660 ;
        RECT 75.050 38.660 75.370 38.720 ;
        RECT 80.585 38.660 80.875 38.705 ;
        RECT 75.050 38.520 80.875 38.660 ;
        RECT 61.710 38.460 62.030 38.520 ;
        RECT 75.050 38.460 75.370 38.520 ;
        RECT 80.585 38.475 80.875 38.520 ;
        RECT 82.870 38.460 83.190 38.720 ;
        RECT 84.265 38.660 84.555 38.705 ;
        RECT 87.930 38.660 88.250 38.720 ;
        RECT 84.265 38.520 88.250 38.660 ;
        RECT 84.265 38.475 84.555 38.520 ;
        RECT 87.930 38.460 88.250 38.520 ;
        RECT 102.650 38.460 102.970 38.720 ;
        RECT 110.010 38.460 110.330 38.720 ;
        RECT 5.520 37.840 118.680 38.320 ;
        RECT 19.405 37.640 19.695 37.685 ;
        RECT 21.230 37.640 21.550 37.700 ;
        RECT 19.405 37.500 21.550 37.640 ;
        RECT 19.405 37.455 19.695 37.500 ;
        RECT 21.230 37.440 21.550 37.500 ;
        RECT 35.490 37.440 35.810 37.700 ;
        RECT 46.530 37.440 46.850 37.700 ;
        RECT 46.990 37.440 47.310 37.700 ;
        RECT 58.490 37.640 58.810 37.700 ;
        RECT 61.725 37.640 62.015 37.685 ;
        RECT 58.490 37.500 62.015 37.640 ;
        RECT 58.490 37.440 58.810 37.500 ;
        RECT 61.725 37.455 62.015 37.500 ;
        RECT 82.425 37.640 82.715 37.685 ;
        RECT 86.550 37.640 86.870 37.700 ;
        RECT 82.425 37.500 86.870 37.640 ;
        RECT 82.425 37.455 82.715 37.500 ;
        RECT 86.550 37.440 86.870 37.500 ;
        RECT 87.010 37.440 87.330 37.700 ;
        RECT 88.850 37.440 89.170 37.700 ;
        RECT 89.310 37.440 89.630 37.700 ;
        RECT 91.165 37.640 91.455 37.685 ;
        RECT 102.650 37.640 102.970 37.700 ;
        RECT 91.165 37.500 102.970 37.640 ;
        RECT 91.165 37.455 91.455 37.500 ;
        RECT 102.650 37.440 102.970 37.500 ;
        RECT 103.110 37.640 103.430 37.700 ;
        RECT 106.805 37.640 107.095 37.685 ;
        RECT 103.110 37.500 107.095 37.640 ;
        RECT 103.110 37.440 103.430 37.500 ;
        RECT 106.805 37.455 107.095 37.500 ;
        RECT 20.770 37.300 21.090 37.360 ;
        RECT 23.085 37.300 23.375 37.345 ;
        RECT 20.770 37.160 23.375 37.300 ;
        RECT 20.770 37.100 21.090 37.160 ;
        RECT 23.085 37.115 23.375 37.160 ;
        RECT 30.445 37.300 30.735 37.345 ;
        RECT 57.110 37.300 57.430 37.360 ;
        RECT 58.045 37.300 58.335 37.345 ;
        RECT 60.330 37.300 60.650 37.360 ;
        RECT 60.805 37.300 61.095 37.345 ;
        RECT 30.445 37.160 34.340 37.300 ;
        RECT 30.445 37.115 30.735 37.160 ;
        RECT 22.610 36.760 22.930 37.020 ;
        RECT 27.210 36.760 27.530 37.020 ;
        RECT 34.200 37.005 34.340 37.160 ;
        RECT 57.110 37.160 58.720 37.300 ;
        RECT 57.110 37.100 57.430 37.160 ;
        RECT 58.045 37.115 58.335 37.160 ;
        RECT 58.580 37.020 58.720 37.160 ;
        RECT 60.330 37.160 61.095 37.300 ;
        RECT 60.330 37.100 60.650 37.160 ;
        RECT 60.805 37.115 61.095 37.160 ;
        RECT 75.050 37.100 75.370 37.360 ;
        RECT 77.345 37.300 77.995 37.345 ;
        RECT 80.945 37.300 81.235 37.345 ;
        RECT 83.805 37.300 84.095 37.345 ;
        RECT 95.290 37.300 95.610 37.360 ;
        RECT 77.345 37.160 84.095 37.300 ;
        RECT 77.345 37.115 77.995 37.160 ;
        RECT 80.645 37.115 81.235 37.160 ;
        RECT 83.805 37.115 84.095 37.160 ;
        RECT 86.640 37.160 95.610 37.300 ;
        RECT 32.745 36.775 33.035 37.005 ;
        RECT 34.125 36.775 34.415 37.005 ;
        RECT 23.990 36.620 24.310 36.680 ;
        RECT 25.845 36.620 26.135 36.665 ;
        RECT 27.670 36.620 27.990 36.680 ;
        RECT 23.990 36.480 27.990 36.620 ;
        RECT 23.990 36.420 24.310 36.480 ;
        RECT 25.845 36.435 26.135 36.480 ;
        RECT 27.670 36.420 27.990 36.480 ;
        RECT 32.820 36.280 32.960 36.775 ;
        RECT 58.490 36.760 58.810 37.020 ;
        RECT 74.150 36.960 74.440 37.005 ;
        RECT 75.985 36.960 76.275 37.005 ;
        RECT 79.565 36.960 79.855 37.005 ;
        RECT 74.150 36.820 79.855 36.960 ;
        RECT 74.150 36.775 74.440 36.820 ;
        RECT 75.985 36.775 76.275 36.820 ;
        RECT 79.565 36.775 79.855 36.820 ;
        RECT 80.645 36.800 80.935 37.115 ;
        RECT 86.640 37.005 86.780 37.160 ;
        RECT 95.290 37.100 95.610 37.160 ;
        RECT 101.725 37.300 102.375 37.345 ;
        RECT 104.490 37.300 104.810 37.360 ;
        RECT 105.325 37.300 105.615 37.345 ;
        RECT 101.725 37.160 105.615 37.300 ;
        RECT 101.725 37.115 102.375 37.160 ;
        RECT 104.490 37.100 104.810 37.160 ;
        RECT 105.025 37.115 105.615 37.160 ;
        RECT 84.265 36.960 84.555 37.005 ;
        RECT 81.120 36.820 85.860 36.960 ;
        RECT 33.650 36.620 33.970 36.680 ;
        RECT 38.265 36.620 38.555 36.665 ;
        RECT 33.650 36.480 38.555 36.620 ;
        RECT 33.650 36.420 33.970 36.480 ;
        RECT 38.265 36.435 38.555 36.480 ;
        RECT 47.910 36.420 48.230 36.680 ;
        RECT 59.410 36.620 59.730 36.680 ;
        RECT 60.345 36.620 60.635 36.665 ;
        RECT 64.930 36.620 65.250 36.680 ;
        RECT 59.410 36.480 65.250 36.620 ;
        RECT 59.410 36.420 59.730 36.480 ;
        RECT 60.345 36.435 60.635 36.480 ;
        RECT 64.930 36.420 65.250 36.480 ;
        RECT 73.670 36.420 73.990 36.680 ;
        RECT 81.120 36.620 81.260 36.820 ;
        RECT 84.265 36.775 84.555 36.820 ;
        RECT 74.220 36.480 81.260 36.620 ;
        RECT 41.930 36.280 42.250 36.340 ;
        RECT 32.820 36.140 42.250 36.280 ;
        RECT 41.930 36.080 42.250 36.140 ;
        RECT 56.650 36.280 56.970 36.340 ;
        RECT 58.045 36.280 58.335 36.325 ;
        RECT 61.710 36.280 62.030 36.340 ;
        RECT 56.650 36.140 62.030 36.280 ;
        RECT 56.650 36.080 56.970 36.140 ;
        RECT 58.045 36.095 58.335 36.140 ;
        RECT 61.710 36.080 62.030 36.140 ;
        RECT 72.290 36.280 72.610 36.340 ;
        RECT 74.220 36.280 74.360 36.480 ;
        RECT 72.290 36.140 74.360 36.280 ;
        RECT 74.555 36.280 74.845 36.325 ;
        RECT 76.445 36.280 76.735 36.325 ;
        RECT 79.565 36.280 79.855 36.325 ;
        RECT 74.555 36.140 79.855 36.280 ;
        RECT 72.290 36.080 72.610 36.140 ;
        RECT 74.555 36.095 74.845 36.140 ;
        RECT 76.445 36.095 76.735 36.140 ;
        RECT 79.565 36.095 79.855 36.140 ;
        RECT 32.285 35.940 32.575 35.985 ;
        RECT 32.730 35.940 33.050 36.000 ;
        RECT 32.285 35.800 33.050 35.940 ;
        RECT 32.285 35.755 32.575 35.800 ;
        RECT 32.730 35.740 33.050 35.800 ;
        RECT 33.190 35.740 33.510 36.000 ;
        RECT 43.770 35.940 44.090 36.000 ;
        RECT 44.705 35.940 44.995 35.985 ;
        RECT 43.770 35.800 44.995 35.940 ;
        RECT 85.720 35.940 85.860 36.820 ;
        RECT 86.565 36.775 86.855 37.005 ;
        RECT 87.470 36.960 87.790 37.020 ;
        RECT 94.385 36.960 94.675 37.005 ;
        RECT 96.670 36.960 96.990 37.020 ;
        RECT 87.100 36.820 92.760 36.960 ;
        RECT 86.105 36.620 86.395 36.665 ;
        RECT 87.100 36.620 87.240 36.820 ;
        RECT 87.470 36.760 87.790 36.820 ;
        RECT 86.105 36.480 87.240 36.620 ;
        RECT 86.105 36.435 86.395 36.480 ;
        RECT 86.640 36.340 86.780 36.480 ;
        RECT 91.610 36.420 91.930 36.680 ;
        RECT 92.620 36.665 92.760 36.820 ;
        RECT 94.385 36.820 96.990 36.960 ;
        RECT 94.385 36.775 94.675 36.820 ;
        RECT 96.670 36.760 96.990 36.820 ;
        RECT 98.530 36.960 98.820 37.005 ;
        RECT 100.365 36.960 100.655 37.005 ;
        RECT 103.945 36.960 104.235 37.005 ;
        RECT 98.530 36.820 104.235 36.960 ;
        RECT 98.530 36.775 98.820 36.820 ;
        RECT 100.365 36.775 100.655 36.820 ;
        RECT 103.945 36.775 104.235 36.820 ;
        RECT 105.025 36.800 105.315 37.115 ;
        RECT 92.545 36.620 92.835 36.665 ;
        RECT 94.830 36.620 95.150 36.680 ;
        RECT 92.545 36.480 95.150 36.620 ;
        RECT 92.545 36.435 92.835 36.480 ;
        RECT 94.830 36.420 95.150 36.480 ;
        RECT 98.065 36.435 98.355 36.665 ;
        RECT 99.445 36.620 99.735 36.665 ;
        RECT 110.010 36.620 110.330 36.680 ;
        RECT 99.445 36.480 110.330 36.620 ;
        RECT 99.445 36.435 99.735 36.480 ;
        RECT 86.550 36.080 86.870 36.340 ;
        RECT 88.390 36.280 88.710 36.340 ;
        RECT 98.140 36.280 98.280 36.435 ;
        RECT 110.010 36.420 110.330 36.480 ;
        RECT 88.390 36.140 98.280 36.280 ;
        RECT 98.935 36.280 99.225 36.325 ;
        RECT 100.825 36.280 101.115 36.325 ;
        RECT 103.945 36.280 104.235 36.325 ;
        RECT 98.935 36.140 104.235 36.280 ;
        RECT 88.390 36.080 88.710 36.140 ;
        RECT 98.935 36.095 99.225 36.140 ;
        RECT 100.825 36.095 101.115 36.140 ;
        RECT 103.945 36.095 104.235 36.140 ;
        RECT 87.010 35.940 87.330 36.000 ;
        RECT 85.720 35.800 87.330 35.940 ;
        RECT 43.770 35.740 44.090 35.800 ;
        RECT 44.705 35.755 44.995 35.800 ;
        RECT 87.010 35.740 87.330 35.800 ;
        RECT 93.910 35.740 94.230 36.000 ;
        RECT 5.520 35.120 118.680 35.600 ;
        RECT 27.620 34.920 27.910 34.965 ;
        RECT 33.190 34.920 33.510 34.980 ;
        RECT 27.620 34.780 33.510 34.920 ;
        RECT 27.620 34.735 27.910 34.780 ;
        RECT 33.190 34.720 33.510 34.780 ;
        RECT 33.650 34.920 33.970 34.980 ;
        RECT 35.045 34.920 35.335 34.965 ;
        RECT 33.650 34.780 35.335 34.920 ;
        RECT 33.650 34.720 33.970 34.780 ;
        RECT 35.045 34.735 35.335 34.780 ;
        RECT 82.870 34.920 83.190 34.980 ;
        RECT 87.850 34.920 88.140 34.965 ;
        RECT 82.870 34.780 88.140 34.920 ;
        RECT 82.870 34.720 83.190 34.780 ;
        RECT 87.850 34.735 88.140 34.780 ;
        RECT 95.290 34.720 95.610 34.980 ;
        RECT 27.175 34.580 27.465 34.625 ;
        RECT 29.065 34.580 29.355 34.625 ;
        RECT 32.185 34.580 32.475 34.625 ;
        RECT 27.175 34.440 32.475 34.580 ;
        RECT 27.175 34.395 27.465 34.440 ;
        RECT 29.065 34.395 29.355 34.440 ;
        RECT 32.185 34.395 32.475 34.440 ;
        RECT 73.670 34.580 73.990 34.640 ;
        RECT 83.790 34.580 84.110 34.640 ;
        RECT 87.435 34.580 87.725 34.625 ;
        RECT 89.325 34.580 89.615 34.625 ;
        RECT 92.445 34.580 92.735 34.625 ;
        RECT 73.670 34.440 86.780 34.580 ;
        RECT 73.670 34.380 73.990 34.440 ;
        RECT 83.790 34.380 84.110 34.440 ;
        RECT 14.790 34.240 15.110 34.300 ;
        RECT 26.305 34.240 26.595 34.285 ;
        RECT 14.790 34.100 26.595 34.240 ;
        RECT 14.790 34.040 15.110 34.100 ;
        RECT 26.305 34.055 26.595 34.100 ;
        RECT 41.930 34.240 42.250 34.300 ;
        RECT 42.850 34.240 43.170 34.300 ;
        RECT 60.790 34.240 61.110 34.300 ;
        RECT 67.230 34.240 67.550 34.300 ;
        RECT 68.625 34.240 68.915 34.285 ;
        RECT 70.910 34.240 71.230 34.300 ;
        RECT 41.930 34.100 45.380 34.240 ;
        RECT 41.930 34.040 42.250 34.100 ;
        RECT 42.850 34.040 43.170 34.100 ;
        RECT 19.850 33.700 20.170 33.960 ;
        RECT 23.070 33.700 23.390 33.960 ;
        RECT 26.770 33.900 27.060 33.945 ;
        RECT 28.605 33.900 28.895 33.945 ;
        RECT 32.185 33.900 32.475 33.945 ;
        RECT 26.770 33.760 32.475 33.900 ;
        RECT 26.770 33.715 27.060 33.760 ;
        RECT 28.605 33.715 28.895 33.760 ;
        RECT 32.185 33.715 32.475 33.760 ;
        RECT 29.965 33.560 30.615 33.605 ;
        RECT 32.730 33.560 33.050 33.620 ;
        RECT 33.265 33.605 33.555 33.920 ;
        RECT 43.770 33.700 44.090 33.960 ;
        RECT 45.240 33.945 45.380 34.100 ;
        RECT 60.790 34.100 71.230 34.240 ;
        RECT 60.790 34.040 61.110 34.100 ;
        RECT 67.230 34.040 67.550 34.100 ;
        RECT 68.625 34.055 68.915 34.100 ;
        RECT 70.910 34.040 71.230 34.100 ;
        RECT 75.985 34.240 76.275 34.285 ;
        RECT 86.090 34.240 86.410 34.300 ;
        RECT 86.640 34.285 86.780 34.440 ;
        RECT 87.435 34.440 92.735 34.580 ;
        RECT 87.435 34.395 87.725 34.440 ;
        RECT 89.325 34.395 89.615 34.440 ;
        RECT 92.445 34.395 92.735 34.440 ;
        RECT 75.985 34.100 86.410 34.240 ;
        RECT 75.985 34.055 76.275 34.100 ;
        RECT 86.090 34.040 86.410 34.100 ;
        RECT 86.565 34.240 86.855 34.285 ;
        RECT 88.390 34.240 88.710 34.300 ;
        RECT 86.565 34.100 88.710 34.240 ;
        RECT 86.565 34.055 86.855 34.100 ;
        RECT 88.390 34.040 88.710 34.100 ;
        RECT 96.670 34.040 96.990 34.300 ;
        RECT 103.125 34.240 103.415 34.285 ;
        RECT 104.490 34.240 104.810 34.300 ;
        RECT 103.125 34.100 104.810 34.240 ;
        RECT 103.125 34.055 103.415 34.100 ;
        RECT 104.490 34.040 104.810 34.100 ;
        RECT 45.165 33.715 45.455 33.945 ;
        RECT 71.845 33.900 72.135 33.945 ;
        RECT 75.525 33.900 75.815 33.945 ;
        RECT 76.430 33.900 76.750 33.960 ;
        RECT 71.845 33.760 73.440 33.900 ;
        RECT 71.845 33.715 72.135 33.760 ;
        RECT 33.265 33.560 33.855 33.605 ;
        RECT 29.965 33.420 33.855 33.560 ;
        RECT 29.965 33.375 30.615 33.420 ;
        RECT 32.730 33.360 33.050 33.420 ;
        RECT 33.565 33.375 33.855 33.420 ;
        RECT 16.630 33.220 16.950 33.280 ;
        RECT 18.945 33.220 19.235 33.265 ;
        RECT 16.630 33.080 19.235 33.220 ;
        RECT 16.630 33.020 16.950 33.080 ;
        RECT 18.945 33.035 19.235 33.080 ;
        RECT 25.845 33.220 26.135 33.265 ;
        RECT 26.750 33.220 27.070 33.280 ;
        RECT 25.845 33.080 27.070 33.220 ;
        RECT 25.845 33.035 26.135 33.080 ;
        RECT 26.750 33.020 27.070 33.080 ;
        RECT 42.390 33.220 42.710 33.280 ;
        RECT 42.865 33.220 43.155 33.265 ;
        RECT 42.390 33.080 43.155 33.220 ;
        RECT 42.390 33.020 42.710 33.080 ;
        RECT 42.865 33.035 43.155 33.080 ;
        RECT 45.150 33.220 45.470 33.280 ;
        RECT 45.625 33.220 45.915 33.265 ;
        RECT 45.150 33.080 45.915 33.220 ;
        RECT 45.150 33.020 45.470 33.080 ;
        RECT 45.625 33.035 45.915 33.080 ;
        RECT 59.870 33.220 60.190 33.280 ;
        RECT 65.865 33.220 66.155 33.265 ;
        RECT 59.870 33.080 66.155 33.220 ;
        RECT 59.870 33.020 60.190 33.080 ;
        RECT 65.865 33.035 66.155 33.080 ;
        RECT 72.750 33.020 73.070 33.280 ;
        RECT 73.300 33.265 73.440 33.760 ;
        RECT 75.525 33.760 76.750 33.900 ;
        RECT 75.525 33.715 75.815 33.760 ;
        RECT 76.430 33.700 76.750 33.760 ;
        RECT 77.350 33.700 77.670 33.960 ;
        RECT 87.030 33.900 87.320 33.945 ;
        RECT 88.865 33.900 89.155 33.945 ;
        RECT 92.445 33.900 92.735 33.945 ;
        RECT 87.030 33.760 92.735 33.900 ;
        RECT 87.030 33.715 87.320 33.760 ;
        RECT 88.865 33.715 89.155 33.760 ;
        RECT 92.445 33.715 92.735 33.760 ;
        RECT 93.525 33.605 93.815 33.920 ;
        RECT 96.760 33.900 96.900 34.040 ;
        RECT 97.145 33.900 97.435 33.945 ;
        RECT 102.665 33.900 102.955 33.945 ;
        RECT 96.760 33.760 102.955 33.900 ;
        RECT 97.145 33.715 97.435 33.760 ;
        RECT 102.665 33.715 102.955 33.760 ;
        RECT 90.225 33.560 90.875 33.605 ;
        RECT 93.525 33.560 94.115 33.605 ;
        RECT 96.685 33.560 96.975 33.605 ;
        RECT 90.225 33.420 96.975 33.560 ;
        RECT 90.225 33.375 90.875 33.420 ;
        RECT 93.825 33.375 94.115 33.420 ;
        RECT 96.685 33.375 96.975 33.420 ;
        RECT 73.225 33.035 73.515 33.265 ;
        RECT 75.050 33.020 75.370 33.280 ;
        RECT 5.520 32.400 118.680 32.880 ;
        RECT 19.850 32.200 20.170 32.260 ;
        RECT 24.465 32.200 24.755 32.245 ;
        RECT 19.850 32.060 24.755 32.200 ;
        RECT 19.850 32.000 20.170 32.060 ;
        RECT 24.465 32.015 24.755 32.060 ;
        RECT 31.825 32.015 32.115 32.245 ;
        RECT 46.990 32.200 47.310 32.260 ;
        RECT 49.535 32.200 49.825 32.245 ;
        RECT 46.990 32.060 49.825 32.200 ;
        RECT 16.630 31.660 16.950 31.920 ;
        RECT 18.925 31.860 19.575 31.905 ;
        RECT 22.525 31.860 22.815 31.905 ;
        RECT 23.530 31.860 23.850 31.920 ;
        RECT 18.925 31.720 23.850 31.860 ;
        RECT 18.925 31.675 19.575 31.720 ;
        RECT 22.225 31.675 22.815 31.720 ;
        RECT 13.870 31.320 14.190 31.580 ;
        RECT 14.790 31.520 15.110 31.580 ;
        RECT 15.265 31.520 15.555 31.565 ;
        RECT 14.790 31.380 15.555 31.520 ;
        RECT 14.790 31.320 15.110 31.380 ;
        RECT 15.265 31.335 15.555 31.380 ;
        RECT 15.730 31.520 16.020 31.565 ;
        RECT 17.565 31.520 17.855 31.565 ;
        RECT 21.145 31.520 21.435 31.565 ;
        RECT 15.730 31.380 21.435 31.520 ;
        RECT 15.730 31.335 16.020 31.380 ;
        RECT 17.565 31.335 17.855 31.380 ;
        RECT 21.145 31.335 21.435 31.380 ;
        RECT 22.225 31.360 22.515 31.675 ;
        RECT 23.530 31.660 23.850 31.720 ;
        RECT 26.305 31.520 26.595 31.565 ;
        RECT 30.905 31.520 31.195 31.565 ;
        RECT 31.900 31.520 32.040 32.015 ;
        RECT 46.990 32.000 47.310 32.060 ;
        RECT 49.535 32.015 49.825 32.060 ;
        RECT 55.745 32.200 56.035 32.245 ;
        RECT 56.650 32.200 56.970 32.260 ;
        RECT 55.745 32.060 56.970 32.200 ;
        RECT 55.745 32.015 56.035 32.060 ;
        RECT 56.650 32.000 56.970 32.060 ;
        RECT 61.725 32.015 62.015 32.245 ;
        RECT 63.090 32.200 63.410 32.260 ;
        RECT 66.770 32.200 67.090 32.260 ;
        RECT 63.090 32.060 67.090 32.200 ;
        RECT 41.490 31.860 41.780 31.905 ;
        RECT 43.350 31.860 43.640 31.905 ;
        RECT 41.490 31.720 43.640 31.860 ;
        RECT 41.490 31.675 41.780 31.720 ;
        RECT 43.350 31.675 43.640 31.720 ;
        RECT 44.270 31.860 44.560 31.905 ;
        RECT 45.150 31.860 45.470 31.920 ;
        RECT 47.530 31.860 47.820 31.905 ;
        RECT 44.270 31.720 47.820 31.860 ;
        RECT 44.270 31.675 44.560 31.720 ;
        RECT 26.305 31.380 30.660 31.520 ;
        RECT 26.305 31.335 26.595 31.380 ;
        RECT 23.070 31.180 23.390 31.240 ;
        RECT 24.005 31.180 24.295 31.225 ;
        RECT 26.750 31.180 27.070 31.240 ;
        RECT 23.070 31.040 24.295 31.180 ;
        RECT 23.070 30.980 23.390 31.040 ;
        RECT 24.005 30.995 24.295 31.040 ;
        RECT 24.540 31.040 27.070 31.180 ;
        RECT 16.135 30.840 16.425 30.885 ;
        RECT 18.025 30.840 18.315 30.885 ;
        RECT 21.145 30.840 21.435 30.885 ;
        RECT 16.135 30.700 21.435 30.840 ;
        RECT 16.135 30.655 16.425 30.700 ;
        RECT 18.025 30.655 18.315 30.700 ;
        RECT 21.145 30.655 21.435 30.700 ;
        RECT 14.805 30.500 15.095 30.545 ;
        RECT 15.250 30.500 15.570 30.560 ;
        RECT 14.805 30.360 15.570 30.500 ;
        RECT 14.805 30.315 15.095 30.360 ;
        RECT 15.250 30.300 15.570 30.360 ;
        RECT 20.310 30.500 20.630 30.560 ;
        RECT 24.540 30.500 24.680 31.040 ;
        RECT 26.750 30.980 27.070 31.040 ;
        RECT 27.685 30.995 27.975 31.225 ;
        RECT 30.520 31.180 30.660 31.380 ;
        RECT 30.905 31.380 32.040 31.520 ;
        RECT 33.665 31.520 33.955 31.565 ;
        RECT 33.665 31.380 36.180 31.520 ;
        RECT 30.905 31.335 31.195 31.380 ;
        RECT 33.665 31.335 33.955 31.380 ;
        RECT 31.810 31.180 32.130 31.240 ;
        RECT 34.125 31.180 34.415 31.225 ;
        RECT 30.520 31.040 34.415 31.180 ;
        RECT 24.910 30.840 25.230 30.900 ;
        RECT 27.760 30.840 27.900 30.995 ;
        RECT 31.810 30.980 32.130 31.040 ;
        RECT 34.125 30.995 34.415 31.040 ;
        RECT 35.030 30.980 35.350 31.240 ;
        RECT 35.120 30.840 35.260 30.980 ;
        RECT 24.910 30.700 35.260 30.840 ;
        RECT 36.040 30.840 36.180 31.380 ;
        RECT 36.410 31.320 36.730 31.580 ;
        RECT 40.105 31.520 40.395 31.565 ;
        RECT 41.930 31.520 42.250 31.580 ;
        RECT 40.105 31.380 42.250 31.520 ;
        RECT 40.105 31.335 40.395 31.380 ;
        RECT 41.930 31.320 42.250 31.380 ;
        RECT 42.390 31.320 42.710 31.580 ;
        RECT 43.425 31.520 43.640 31.675 ;
        RECT 45.150 31.660 45.470 31.720 ;
        RECT 47.530 31.675 47.820 31.720 ;
        RECT 56.205 31.860 56.495 31.905 ;
        RECT 59.410 31.860 59.730 31.920 ;
        RECT 56.205 31.720 59.730 31.860 ;
        RECT 61.800 31.860 61.940 32.015 ;
        RECT 63.090 32.000 63.410 32.060 ;
        RECT 66.770 32.000 67.090 32.060 ;
        RECT 70.910 32.000 71.230 32.260 ;
        RECT 75.050 32.200 75.370 32.260 ;
        RECT 85.645 32.200 85.935 32.245 ;
        RECT 75.050 32.060 85.935 32.200 ;
        RECT 75.050 32.000 75.370 32.060 ;
        RECT 85.645 32.015 85.935 32.060 ;
        RECT 63.565 31.860 63.855 31.905 ;
        RECT 61.800 31.720 63.855 31.860 ;
        RECT 56.205 31.675 56.495 31.720 ;
        RECT 59.410 31.660 59.730 31.720 ;
        RECT 63.565 31.675 63.855 31.720 ;
        RECT 65.845 31.860 66.495 31.905 ;
        RECT 67.230 31.860 67.550 31.920 ;
        RECT 69.445 31.860 69.735 31.905 ;
        RECT 65.845 31.720 69.735 31.860 ;
        RECT 65.845 31.675 66.495 31.720 ;
        RECT 67.230 31.660 67.550 31.720 ;
        RECT 69.145 31.675 69.735 31.720 ;
        RECT 72.750 31.860 73.070 31.920 ;
        RECT 73.225 31.860 73.515 31.905 ;
        RECT 72.750 31.720 73.515 31.860 ;
        RECT 45.670 31.520 45.960 31.565 ;
        RECT 43.425 31.380 45.960 31.520 ;
        RECT 45.670 31.335 45.960 31.380 ;
        RECT 56.665 31.520 56.955 31.565 ;
        RECT 58.490 31.520 58.810 31.580 ;
        RECT 56.665 31.380 58.810 31.520 ;
        RECT 56.665 31.335 56.955 31.380 ;
        RECT 58.490 31.320 58.810 31.380 ;
        RECT 59.870 31.320 60.190 31.580 ;
        RECT 62.650 31.520 62.940 31.565 ;
        RECT 64.485 31.520 64.775 31.565 ;
        RECT 68.065 31.520 68.355 31.565 ;
        RECT 62.650 31.380 68.355 31.520 ;
        RECT 62.650 31.335 62.940 31.380 ;
        RECT 64.485 31.335 64.775 31.380 ;
        RECT 68.065 31.335 68.355 31.380 ;
        RECT 69.145 31.360 69.435 31.675 ;
        RECT 72.750 31.660 73.070 31.720 ;
        RECT 73.225 31.675 73.515 31.720 ;
        RECT 75.505 31.860 76.155 31.905 ;
        RECT 79.105 31.860 79.395 31.905 ;
        RECT 75.505 31.720 79.395 31.860 ;
        RECT 75.505 31.675 76.155 31.720 ;
        RECT 78.805 31.675 79.395 31.720 ;
        RECT 83.790 31.860 84.110 31.920 ;
        RECT 88.410 31.860 88.700 31.905 ;
        RECT 90.270 31.860 90.560 31.905 ;
        RECT 83.790 31.720 87.700 31.860 ;
        RECT 78.805 31.580 79.095 31.675 ;
        RECT 83.790 31.660 84.110 31.720 ;
        RECT 72.310 31.520 72.600 31.565 ;
        RECT 74.145 31.520 74.435 31.565 ;
        RECT 77.725 31.520 78.015 31.565 ;
        RECT 72.310 31.380 78.015 31.520 ;
        RECT 72.310 31.335 72.600 31.380 ;
        RECT 74.145 31.335 74.435 31.380 ;
        RECT 77.725 31.335 78.015 31.380 ;
        RECT 78.730 31.360 79.095 31.580 ;
        RECT 87.560 31.565 87.700 31.720 ;
        RECT 88.410 31.720 90.560 31.860 ;
        RECT 88.410 31.675 88.700 31.720 ;
        RECT 90.270 31.675 90.560 31.720 ;
        RECT 91.190 31.860 91.480 31.905 ;
        RECT 93.910 31.860 94.230 31.920 ;
        RECT 94.450 31.860 94.740 31.905 ;
        RECT 91.190 31.720 94.740 31.860 ;
        RECT 91.190 31.675 91.480 31.720 ;
        RECT 81.045 31.520 81.335 31.565 ;
        RECT 85.185 31.520 85.475 31.565 ;
        RECT 81.045 31.380 83.560 31.520 ;
        RECT 78.730 31.320 79.050 31.360 ;
        RECT 81.045 31.335 81.335 31.380 ;
        RECT 36.500 31.180 36.640 31.320 ;
        RECT 39.170 31.180 39.490 31.240 ;
        RECT 40.565 31.180 40.855 31.225 ;
        RECT 36.500 31.040 40.855 31.180 ;
        RECT 39.170 30.980 39.490 31.040 ;
        RECT 40.565 30.995 40.855 31.040 ;
        RECT 52.970 31.180 53.290 31.240 ;
        RECT 54.825 31.180 55.115 31.225 ;
        RECT 52.970 31.040 55.115 31.180 ;
        RECT 52.970 30.980 53.290 31.040 ;
        RECT 54.825 30.995 55.115 31.040 ;
        RECT 59.425 31.180 59.715 31.225 ;
        RECT 61.710 31.180 62.030 31.240 ;
        RECT 59.425 31.040 62.030 31.180 ;
        RECT 59.425 30.995 59.715 31.040 ;
        RECT 41.030 30.840 41.320 30.885 ;
        RECT 42.890 30.840 43.180 30.885 ;
        RECT 45.670 30.840 45.960 30.885 ;
        RECT 36.040 30.700 39.860 30.840 ;
        RECT 24.910 30.640 25.230 30.700 ;
        RECT 20.310 30.360 24.680 30.500 ;
        RECT 28.590 30.500 28.910 30.560 ;
        RECT 29.985 30.500 30.275 30.545 ;
        RECT 28.590 30.360 30.275 30.500 ;
        RECT 20.310 30.300 20.630 30.360 ;
        RECT 28.590 30.300 28.910 30.360 ;
        RECT 29.985 30.315 30.275 30.360 ;
        RECT 39.170 30.300 39.490 30.560 ;
        RECT 39.720 30.500 39.860 30.700 ;
        RECT 41.030 30.700 45.960 30.840 ;
        RECT 41.030 30.655 41.320 30.700 ;
        RECT 42.890 30.655 43.180 30.700 ;
        RECT 45.670 30.655 45.960 30.700 ;
        RECT 56.205 30.840 56.495 30.885 ;
        RECT 59.500 30.840 59.640 30.995 ;
        RECT 61.710 30.980 62.030 31.040 ;
        RECT 62.185 31.180 62.475 31.225 ;
        RECT 71.845 31.180 72.135 31.225 ;
        RECT 73.670 31.180 73.990 31.240 ;
        RECT 62.185 31.040 73.990 31.180 ;
        RECT 62.185 30.995 62.475 31.040 ;
        RECT 69.160 30.900 69.300 31.040 ;
        RECT 71.845 30.995 72.135 31.040 ;
        RECT 73.670 30.980 73.990 31.040 ;
        RECT 80.570 30.980 80.890 31.240 ;
        RECT 56.205 30.700 59.640 30.840 ;
        RECT 63.055 30.840 63.345 30.885 ;
        RECT 64.945 30.840 65.235 30.885 ;
        RECT 68.065 30.840 68.355 30.885 ;
        RECT 63.055 30.700 68.355 30.840 ;
        RECT 56.205 30.655 56.495 30.700 ;
        RECT 63.055 30.655 63.345 30.700 ;
        RECT 64.945 30.655 65.235 30.700 ;
        RECT 68.065 30.655 68.355 30.700 ;
        RECT 69.070 30.640 69.390 30.900 ;
        RECT 83.420 30.885 83.560 31.380 ;
        RECT 85.185 31.380 87.240 31.520 ;
        RECT 85.185 31.335 85.475 31.380 ;
        RECT 86.550 30.980 86.870 31.240 ;
        RECT 87.100 31.180 87.240 31.380 ;
        RECT 87.485 31.335 87.775 31.565 ;
        RECT 87.930 31.520 88.250 31.580 ;
        RECT 89.325 31.520 89.615 31.565 ;
        RECT 87.930 31.380 89.615 31.520 ;
        RECT 90.345 31.520 90.560 31.675 ;
        RECT 93.910 31.660 94.230 31.720 ;
        RECT 94.450 31.675 94.740 31.720 ;
        RECT 92.590 31.520 92.880 31.565 ;
        RECT 90.345 31.380 92.880 31.520 ;
        RECT 87.930 31.320 88.250 31.380 ;
        RECT 89.325 31.335 89.615 31.380 ;
        RECT 92.590 31.335 92.880 31.380 ;
        RECT 91.610 31.180 91.930 31.240 ;
        RECT 96.455 31.180 96.745 31.225 ;
        RECT 87.100 31.040 96.745 31.180 ;
        RECT 91.610 30.980 91.930 31.040 ;
        RECT 96.455 30.995 96.745 31.040 ;
        RECT 72.715 30.840 73.005 30.885 ;
        RECT 74.605 30.840 74.895 30.885 ;
        RECT 77.725 30.840 78.015 30.885 ;
        RECT 72.715 30.700 78.015 30.840 ;
        RECT 72.715 30.655 73.005 30.700 ;
        RECT 74.605 30.655 74.895 30.700 ;
        RECT 77.725 30.655 78.015 30.700 ;
        RECT 83.345 30.655 83.635 30.885 ;
        RECT 87.950 30.840 88.240 30.885 ;
        RECT 89.810 30.840 90.100 30.885 ;
        RECT 92.590 30.840 92.880 30.885 ;
        RECT 87.950 30.700 92.880 30.840 ;
        RECT 87.950 30.655 88.240 30.700 ;
        RECT 89.810 30.655 90.100 30.700 ;
        RECT 92.590 30.655 92.880 30.700 ;
        RECT 47.450 30.500 47.770 30.560 ;
        RECT 39.720 30.360 47.770 30.500 ;
        RECT 47.450 30.300 47.770 30.360 ;
        RECT 81.965 30.500 82.255 30.545 ;
        RECT 82.410 30.500 82.730 30.560 ;
        RECT 81.965 30.360 82.730 30.500 ;
        RECT 81.965 30.315 82.255 30.360 ;
        RECT 82.410 30.300 82.730 30.360 ;
        RECT 5.520 29.680 118.680 30.160 ;
        RECT 13.870 29.480 14.190 29.540 ;
        RECT 18.945 29.480 19.235 29.525 ;
        RECT 13.870 29.340 19.235 29.480 ;
        RECT 13.870 29.280 14.190 29.340 ;
        RECT 18.945 29.295 19.235 29.340 ;
        RECT 23.530 29.280 23.850 29.540 ;
        RECT 41.930 29.480 42.250 29.540 ;
        RECT 44.705 29.480 44.995 29.525 ;
        RECT 41.930 29.340 44.995 29.480 ;
        RECT 41.930 29.280 42.250 29.340 ;
        RECT 44.705 29.295 44.995 29.340 ;
        RECT 59.885 29.480 60.175 29.525 ;
        RECT 60.330 29.480 60.650 29.540 ;
        RECT 59.885 29.340 60.650 29.480 ;
        RECT 59.885 29.295 60.175 29.340 ;
        RECT 60.330 29.280 60.650 29.340 ;
        RECT 62.630 29.280 62.950 29.540 ;
        RECT 67.230 29.280 67.550 29.540 ;
        RECT 78.730 29.480 79.050 29.540 ;
        RECT 84.725 29.480 85.015 29.525 ;
        RECT 78.730 29.340 85.015 29.480 ;
        RECT 78.730 29.280 79.050 29.340 ;
        RECT 84.725 29.295 85.015 29.340 ;
        RECT 20.770 29.140 21.090 29.200 ;
        RECT 20.770 29.000 21.460 29.140 ;
        RECT 20.770 28.940 21.090 29.000 ;
        RECT 21.320 28.845 21.460 29.000 ;
        RECT 60.805 28.955 61.095 29.185 ;
        RECT 77.925 29.140 78.215 29.185 ;
        RECT 81.045 29.140 81.335 29.185 ;
        RECT 82.935 29.140 83.225 29.185 ;
        RECT 77.925 29.000 83.225 29.140 ;
        RECT 77.925 28.955 78.215 29.000 ;
        RECT 81.045 28.955 81.335 29.000 ;
        RECT 82.935 28.955 83.225 29.000 ;
        RECT 21.245 28.615 21.535 28.845 ;
        RECT 22.150 28.800 22.470 28.860 ;
        RECT 24.910 28.800 25.230 28.860 ;
        RECT 22.150 28.660 25.230 28.800 ;
        RECT 22.150 28.600 22.470 28.660 ;
        RECT 24.910 28.600 25.230 28.660 ;
        RECT 47.910 28.600 48.230 28.860 ;
        RECT 60.880 28.800 61.020 28.955 ;
        RECT 62.645 28.800 62.935 28.845 ;
        RECT 60.880 28.660 62.935 28.800 ;
        RECT 62.645 28.615 62.935 28.660 ;
        RECT 82.410 28.600 82.730 28.860 ;
        RECT 83.790 28.600 84.110 28.860 ;
        RECT 17.090 28.460 17.410 28.520 ;
        RECT 24.005 28.460 24.295 28.505 ;
        RECT 17.090 28.320 38.020 28.460 ;
        RECT 17.090 28.260 17.410 28.320 ;
        RECT 24.005 28.275 24.295 28.320 ;
        RECT 14.790 28.120 15.110 28.180 ;
        RECT 27.210 28.120 27.530 28.180 ;
        RECT 29.525 28.120 29.815 28.165 ;
        RECT 36.410 28.120 36.730 28.180 ;
        RECT 14.790 27.980 36.730 28.120 ;
        RECT 37.880 28.120 38.020 28.320 ;
        RECT 38.250 28.260 38.570 28.520 ;
        RECT 39.645 28.275 39.935 28.505 ;
        RECT 39.720 28.120 39.860 28.275 ;
        RECT 42.850 28.260 43.170 28.520 ;
        RECT 46.545 28.460 46.835 28.505 ;
        RECT 46.990 28.460 47.310 28.520 ;
        RECT 46.545 28.320 47.310 28.460 ;
        RECT 46.545 28.275 46.835 28.320 ;
        RECT 46.990 28.260 47.310 28.320 ;
        RECT 56.650 28.460 56.970 28.520 ;
        RECT 58.045 28.460 58.335 28.505 ;
        RECT 56.650 28.320 58.335 28.460 ;
        RECT 56.650 28.260 56.970 28.320 ;
        RECT 58.045 28.275 58.335 28.320 ;
        RECT 46.070 28.120 46.390 28.180 ;
        RECT 58.120 28.120 58.260 28.275 ;
        RECT 59.870 28.260 60.190 28.520 ;
        RECT 64.010 28.260 64.330 28.520 ;
        RECT 66.770 28.260 67.090 28.520 ;
        RECT 60.330 28.120 60.650 28.180 ;
        RECT 66.860 28.120 67.000 28.260 ;
        RECT 76.845 28.165 77.135 28.480 ;
        RECT 77.925 28.460 78.215 28.505 ;
        RECT 81.505 28.460 81.795 28.505 ;
        RECT 83.340 28.460 83.630 28.505 ;
        RECT 77.925 28.320 83.630 28.460 ;
        RECT 77.925 28.275 78.215 28.320 ;
        RECT 81.505 28.275 81.795 28.320 ;
        RECT 83.340 28.275 83.630 28.320 ;
        RECT 84.265 28.460 84.555 28.505 ;
        RECT 87.010 28.460 87.330 28.520 ;
        RECT 84.265 28.320 87.330 28.460 ;
        RECT 84.265 28.275 84.555 28.320 ;
        RECT 37.880 27.980 48.140 28.120 ;
        RECT 58.120 27.980 60.650 28.120 ;
        RECT 14.790 27.920 15.110 27.980 ;
        RECT 27.210 27.920 27.530 27.980 ;
        RECT 29.525 27.935 29.815 27.980 ;
        RECT 36.410 27.920 36.730 27.980 ;
        RECT 46.070 27.920 46.390 27.980 ;
        RECT 17.550 27.580 17.870 27.840 ;
        RECT 20.310 27.780 20.630 27.840 ;
        RECT 20.785 27.780 21.075 27.825 ;
        RECT 20.310 27.640 21.075 27.780 ;
        RECT 20.310 27.580 20.630 27.640 ;
        RECT 20.785 27.595 21.075 27.640 ;
        RECT 35.030 27.780 35.350 27.840 ;
        RECT 39.185 27.780 39.475 27.825 ;
        RECT 35.030 27.640 39.475 27.780 ;
        RECT 35.030 27.580 35.350 27.640 ;
        RECT 39.185 27.595 39.475 27.640 ;
        RECT 42.850 27.780 43.170 27.840 ;
        RECT 43.325 27.780 43.615 27.825 ;
        RECT 42.850 27.640 43.615 27.780 ;
        RECT 42.850 27.580 43.170 27.640 ;
        RECT 43.325 27.595 43.615 27.640 ;
        RECT 47.005 27.780 47.295 27.825 ;
        RECT 47.450 27.780 47.770 27.840 ;
        RECT 47.005 27.640 47.770 27.780 ;
        RECT 48.000 27.780 48.140 27.980 ;
        RECT 60.330 27.920 60.650 27.980 ;
        RECT 60.880 27.980 67.000 28.120 ;
        RECT 76.545 28.120 77.135 28.165 ;
        RECT 79.650 28.165 79.970 28.180 ;
        RECT 79.650 28.120 80.435 28.165 ;
        RECT 76.545 27.980 80.435 28.120 ;
        RECT 60.880 27.780 61.020 27.980 ;
        RECT 76.545 27.935 76.835 27.980 ;
        RECT 79.650 27.935 80.435 27.980 ;
        RECT 83.790 28.120 84.110 28.180 ;
        RECT 84.340 28.120 84.480 28.275 ;
        RECT 87.010 28.260 87.330 28.320 ;
        RECT 83.790 27.980 84.480 28.120 ;
        RECT 79.650 27.920 79.970 27.935 ;
        RECT 83.790 27.920 84.110 27.980 ;
        RECT 48.000 27.640 61.020 27.780 ;
        RECT 47.005 27.595 47.295 27.640 ;
        RECT 47.450 27.580 47.770 27.640 ;
        RECT 61.250 27.580 61.570 27.840 ;
        RECT 75.065 27.780 75.355 27.825 ;
        RECT 82.410 27.780 82.730 27.840 ;
        RECT 75.065 27.640 82.730 27.780 ;
        RECT 75.065 27.595 75.355 27.640 ;
        RECT 82.410 27.580 82.730 27.640 ;
        RECT 5.520 26.960 118.680 27.440 ;
        RECT 22.625 26.760 22.915 26.805 ;
        RECT 23.990 26.760 24.310 26.820 ;
        RECT 22.625 26.620 24.310 26.760 ;
        RECT 22.625 26.575 22.915 26.620 ;
        RECT 23.990 26.560 24.310 26.620 ;
        RECT 31.810 26.560 32.130 26.820 ;
        RECT 47.450 26.805 47.770 26.820 ;
        RECT 47.235 26.575 47.770 26.805 ;
        RECT 61.725 26.760 62.015 26.805 ;
        RECT 63.185 26.760 63.475 26.805 ;
        RECT 61.725 26.620 63.475 26.760 ;
        RECT 61.725 26.575 62.015 26.620 ;
        RECT 63.185 26.575 63.475 26.620 ;
        RECT 75.050 26.760 75.370 26.820 ;
        RECT 75.525 26.760 75.815 26.805 ;
        RECT 75.050 26.620 75.815 26.760 ;
        RECT 47.450 26.560 47.770 26.575 ;
        RECT 75.050 26.560 75.370 26.620 ;
        RECT 75.525 26.575 75.815 26.620 ;
        RECT 79.650 26.560 79.970 26.820 ;
        RECT 14.790 26.420 15.110 26.480 ;
        RECT 13.960 26.280 15.110 26.420 ;
        RECT 13.960 26.125 14.100 26.280 ;
        RECT 14.790 26.220 15.110 26.280 ;
        RECT 15.250 26.220 15.570 26.480 ;
        RECT 17.550 26.465 17.870 26.480 ;
        RECT 17.545 26.420 18.195 26.465 ;
        RECT 21.145 26.420 21.435 26.465 ;
        RECT 17.545 26.280 21.435 26.420 ;
        RECT 17.545 26.235 18.195 26.280 ;
        RECT 20.845 26.235 21.435 26.280 ;
        RECT 39.190 26.420 39.480 26.465 ;
        RECT 41.050 26.420 41.340 26.465 ;
        RECT 39.190 26.280 41.340 26.420 ;
        RECT 39.190 26.235 39.480 26.280 ;
        RECT 41.050 26.235 41.340 26.280 ;
        RECT 41.970 26.420 42.260 26.465 ;
        RECT 42.850 26.420 43.170 26.480 ;
        RECT 45.230 26.420 45.520 26.465 ;
        RECT 41.970 26.280 45.520 26.420 ;
        RECT 41.970 26.235 42.260 26.280 ;
        RECT 17.550 26.220 17.870 26.235 ;
        RECT 13.885 25.895 14.175 26.125 ;
        RECT 14.350 26.080 14.640 26.125 ;
        RECT 16.185 26.080 16.475 26.125 ;
        RECT 19.765 26.080 20.055 26.125 ;
        RECT 14.350 25.940 20.055 26.080 ;
        RECT 14.350 25.895 14.640 25.940 ;
        RECT 16.185 25.895 16.475 25.940 ;
        RECT 19.765 25.895 20.055 25.940 ;
        RECT 20.845 25.920 21.135 26.235 ;
        RECT 34.570 25.880 34.890 26.140 ;
        RECT 36.410 26.080 36.730 26.140 ;
        RECT 38.265 26.080 38.555 26.125 ;
        RECT 36.410 25.940 38.555 26.080 ;
        RECT 41.125 26.080 41.340 26.235 ;
        RECT 42.850 26.220 43.170 26.280 ;
        RECT 45.230 26.235 45.520 26.280 ;
        RECT 57.570 26.420 57.890 26.480 ;
        RECT 61.250 26.420 61.570 26.480 ;
        RECT 62.185 26.420 62.475 26.465 ;
        RECT 57.570 26.280 62.475 26.420 ;
        RECT 57.570 26.220 57.890 26.280 ;
        RECT 61.250 26.220 61.570 26.280 ;
        RECT 62.185 26.235 62.475 26.280 ;
        RECT 43.370 26.080 43.660 26.125 ;
        RECT 41.125 25.940 43.660 26.080 ;
        RECT 36.410 25.880 36.730 25.940 ;
        RECT 38.265 25.895 38.555 25.940 ;
        RECT 43.370 25.895 43.660 25.940 ;
        RECT 58.490 26.080 58.810 26.140 ;
        RECT 59.425 26.080 59.715 26.125 ;
        RECT 64.010 26.080 64.330 26.140 ;
        RECT 58.490 25.940 64.330 26.080 ;
        RECT 58.490 25.880 58.810 25.940 ;
        RECT 59.425 25.895 59.715 25.940 ;
        RECT 64.010 25.880 64.330 25.940 ;
        RECT 79.205 26.080 79.495 26.125 ;
        RECT 83.790 26.080 84.110 26.140 ;
        RECT 79.205 25.940 84.110 26.080 ;
        RECT 79.205 25.895 79.495 25.940 ;
        RECT 83.790 25.880 84.110 25.940 ;
        RECT 39.170 25.740 39.490 25.800 ;
        RECT 40.105 25.740 40.395 25.785 ;
        RECT 59.870 25.740 60.190 25.800 ;
        RECT 39.170 25.600 40.395 25.740 ;
        RECT 39.170 25.540 39.490 25.600 ;
        RECT 40.105 25.555 40.395 25.600 ;
        RECT 59.500 25.600 60.190 25.740 ;
        RECT 14.755 25.400 15.045 25.445 ;
        RECT 16.645 25.400 16.935 25.445 ;
        RECT 19.765 25.400 20.055 25.445 ;
        RECT 14.755 25.260 20.055 25.400 ;
        RECT 14.755 25.215 15.045 25.260 ;
        RECT 16.645 25.215 16.935 25.260 ;
        RECT 19.765 25.215 20.055 25.260 ;
        RECT 38.730 25.400 39.020 25.445 ;
        RECT 40.590 25.400 40.880 25.445 ;
        RECT 43.370 25.400 43.660 25.445 ;
        RECT 38.730 25.260 43.660 25.400 ;
        RECT 38.730 25.215 39.020 25.260 ;
        RECT 40.590 25.215 40.880 25.260 ;
        RECT 43.370 25.215 43.660 25.260 ;
        RECT 52.970 25.400 53.290 25.460 ;
        RECT 59.500 25.400 59.640 25.600 ;
        RECT 59.870 25.540 60.190 25.600 ;
        RECT 60.330 25.540 60.650 25.800 ;
        RECT 60.805 25.740 61.095 25.785 ;
        RECT 62.630 25.740 62.950 25.800 ;
        RECT 60.805 25.600 62.950 25.740 ;
        RECT 60.805 25.555 61.095 25.600 ;
        RECT 52.970 25.260 59.640 25.400 ;
        RECT 52.970 25.200 53.290 25.260 ;
        RECT 59.410 25.060 59.730 25.120 ;
        RECT 60.880 25.060 61.020 25.555 ;
        RECT 62.630 25.540 62.950 25.600 ;
        RECT 78.745 25.740 79.035 25.785 ;
        RECT 82.410 25.740 82.730 25.800 ;
        RECT 78.745 25.600 82.730 25.740 ;
        RECT 78.745 25.555 79.035 25.600 ;
        RECT 82.410 25.540 82.730 25.600 ;
        RECT 59.410 24.920 61.020 25.060 ;
        RECT 59.410 24.860 59.730 24.920 ;
        RECT 63.090 24.860 63.410 25.120 ;
        RECT 64.025 25.060 64.315 25.105 ;
        RECT 64.470 25.060 64.790 25.120 ;
        RECT 64.025 24.920 64.790 25.060 ;
        RECT 64.025 24.875 64.315 24.920 ;
        RECT 64.470 24.860 64.790 24.920 ;
        RECT 5.520 24.240 118.680 24.720 ;
        RECT 34.570 24.040 34.890 24.100 ;
        RECT 35.965 24.040 36.255 24.085 ;
        RECT 34.570 23.900 36.255 24.040 ;
        RECT 34.570 23.840 34.890 23.900 ;
        RECT 35.965 23.855 36.255 23.900 ;
        RECT 52.050 24.040 52.370 24.100 ;
        RECT 60.330 24.040 60.650 24.100 ;
        RECT 52.050 23.900 60.650 24.040 ;
        RECT 52.050 23.840 52.370 23.900 ;
        RECT 60.330 23.840 60.650 23.900 ;
        RECT 62.185 24.040 62.475 24.085 ;
        RECT 68.150 24.040 68.470 24.100 ;
        RECT 62.185 23.900 68.470 24.040 ;
        RECT 62.185 23.855 62.475 23.900 ;
        RECT 68.150 23.840 68.470 23.900 ;
        RECT 28.095 23.700 28.385 23.745 ;
        RECT 29.985 23.700 30.275 23.745 ;
        RECT 33.105 23.700 33.395 23.745 ;
        RECT 28.095 23.560 33.395 23.700 ;
        RECT 28.095 23.515 28.385 23.560 ;
        RECT 29.985 23.515 30.275 23.560 ;
        RECT 33.105 23.515 33.395 23.560 ;
        RECT 58.505 23.700 58.795 23.745 ;
        RECT 59.410 23.700 59.730 23.760 ;
        RECT 58.505 23.560 59.730 23.700 ;
        RECT 58.505 23.515 58.795 23.560 ;
        RECT 59.410 23.500 59.730 23.560 ;
        RECT 59.870 23.700 60.190 23.760 ;
        RECT 64.025 23.700 64.315 23.745 ;
        RECT 59.870 23.560 64.315 23.700 ;
        RECT 59.870 23.500 60.190 23.560 ;
        RECT 64.025 23.515 64.315 23.560 ;
        RECT 27.210 23.160 27.530 23.420 ;
        RECT 28.590 23.160 28.910 23.420 ;
        RECT 57.110 23.360 57.430 23.420 ;
        RECT 50.300 23.220 57.430 23.360 ;
        RECT 27.690 23.020 27.980 23.065 ;
        RECT 29.525 23.020 29.815 23.065 ;
        RECT 33.105 23.020 33.395 23.065 ;
        RECT 27.690 22.880 33.395 23.020 ;
        RECT 27.690 22.835 27.980 22.880 ;
        RECT 29.525 22.835 29.815 22.880 ;
        RECT 33.105 22.835 33.395 22.880 ;
        RECT 34.185 22.725 34.475 23.040 ;
        RECT 46.070 23.020 46.390 23.080 ;
        RECT 50.300 23.065 50.440 23.220 ;
        RECT 57.110 23.160 57.430 23.220 ;
        RECT 46.545 23.020 46.835 23.065 ;
        RECT 46.070 22.880 46.835 23.020 ;
        RECT 46.070 22.820 46.390 22.880 ;
        RECT 46.545 22.835 46.835 22.880 ;
        RECT 48.845 22.835 49.135 23.065 ;
        RECT 50.225 22.835 50.515 23.065 ;
        RECT 50.685 22.835 50.975 23.065 ;
        RECT 51.605 23.020 51.895 23.065 ;
        RECT 52.970 23.020 53.290 23.080 ;
        RECT 51.605 22.880 53.290 23.020 ;
        RECT 51.605 22.835 51.895 22.880 ;
        RECT 30.885 22.680 31.535 22.725 ;
        RECT 34.185 22.680 34.775 22.725 ;
        RECT 35.030 22.680 35.350 22.740 ;
        RECT 30.885 22.540 35.350 22.680 ;
        RECT 48.920 22.680 49.060 22.835 ;
        RECT 50.760 22.680 50.900 22.835 ;
        RECT 52.970 22.820 53.290 22.880 ;
        RECT 53.890 23.020 54.210 23.080 ;
        RECT 54.365 23.020 54.655 23.065 ;
        RECT 61.250 23.020 61.570 23.080 ;
        RECT 53.890 22.880 61.570 23.020 ;
        RECT 53.890 22.820 54.210 22.880 ;
        RECT 54.365 22.835 54.655 22.880 ;
        RECT 61.250 22.820 61.570 22.880 ;
        RECT 64.470 22.820 64.790 23.080 ;
        RECT 52.050 22.680 52.370 22.740 ;
        RECT 48.920 22.540 52.370 22.680 ;
        RECT 30.885 22.495 31.535 22.540 ;
        RECT 34.485 22.495 34.775 22.540 ;
        RECT 35.030 22.480 35.350 22.540 ;
        RECT 52.050 22.480 52.370 22.540 ;
        RECT 58.490 22.480 58.810 22.740 ;
        RECT 63.105 22.680 63.395 22.725 ;
        RECT 62.030 22.540 63.395 22.680 ;
        RECT 47.005 22.340 47.295 22.385 ;
        RECT 47.450 22.340 47.770 22.400 ;
        RECT 47.005 22.200 47.770 22.340 ;
        RECT 47.005 22.155 47.295 22.200 ;
        RECT 47.450 22.140 47.770 22.200 ;
        RECT 48.370 22.140 48.690 22.400 ;
        RECT 49.290 22.140 49.610 22.400 ;
        RECT 51.605 22.340 51.895 22.385 ;
        RECT 53.430 22.340 53.750 22.400 ;
        RECT 51.605 22.200 53.750 22.340 ;
        RECT 51.605 22.155 51.895 22.200 ;
        RECT 53.430 22.140 53.750 22.200 ;
        RECT 53.905 22.340 54.195 22.385 ;
        RECT 56.650 22.340 56.970 22.400 ;
        RECT 53.905 22.200 56.970 22.340 ;
        RECT 53.905 22.155 54.195 22.200 ;
        RECT 56.650 22.140 56.970 22.200 ;
        RECT 57.585 22.340 57.875 22.385 ;
        RECT 58.030 22.340 58.350 22.400 ;
        RECT 57.585 22.200 58.350 22.340 ;
        RECT 57.585 22.155 57.875 22.200 ;
        RECT 58.030 22.140 58.350 22.200 ;
        RECT 58.950 22.340 59.270 22.400 ;
        RECT 60.805 22.340 61.095 22.385 ;
        RECT 62.030 22.340 62.170 22.540 ;
        RECT 63.105 22.495 63.395 22.540 ;
        RECT 58.950 22.200 62.170 22.340 ;
        RECT 65.405 22.340 65.695 22.385 ;
        RECT 71.830 22.340 72.150 22.400 ;
        RECT 65.405 22.200 72.150 22.340 ;
        RECT 58.950 22.140 59.270 22.200 ;
        RECT 60.805 22.155 61.095 22.200 ;
        RECT 65.405 22.155 65.695 22.200 ;
        RECT 71.830 22.140 72.150 22.200 ;
        RECT 5.520 21.520 118.680 22.000 ;
        RECT 56.205 21.320 56.495 21.365 ;
        RECT 57.110 21.320 57.430 21.380 ;
        RECT 56.205 21.180 57.430 21.320 ;
        RECT 56.205 21.135 56.495 21.180 ;
        RECT 57.110 21.120 57.430 21.180 ;
        RECT 58.505 21.320 58.795 21.365 ;
        RECT 60.330 21.320 60.650 21.380 ;
        RECT 58.505 21.180 60.650 21.320 ;
        RECT 58.505 21.135 58.795 21.180 ;
        RECT 60.330 21.120 60.650 21.180 ;
        RECT 61.250 21.120 61.570 21.380 ;
        RECT 47.450 20.980 47.770 21.040 ;
        RECT 48.365 20.980 49.015 21.025 ;
        RECT 51.965 20.980 52.255 21.025 ;
        RECT 47.450 20.840 52.255 20.980 ;
        RECT 47.450 20.780 47.770 20.840 ;
        RECT 48.365 20.795 49.015 20.840 ;
        RECT 51.665 20.795 52.255 20.840 ;
        RECT 53.430 20.980 53.750 21.040 ;
        RECT 54.365 20.980 54.655 21.025 ;
        RECT 53.430 20.840 54.655 20.980 ;
        RECT 36.410 20.640 36.730 20.700 ;
        RECT 44.690 20.640 45.010 20.700 ;
        RECT 36.410 20.500 45.010 20.640 ;
        RECT 36.410 20.440 36.730 20.500 ;
        RECT 44.690 20.440 45.010 20.500 ;
        RECT 45.170 20.640 45.460 20.685 ;
        RECT 47.005 20.640 47.295 20.685 ;
        RECT 50.585 20.640 50.875 20.685 ;
        RECT 45.170 20.500 50.875 20.640 ;
        RECT 45.170 20.455 45.460 20.500 ;
        RECT 47.005 20.455 47.295 20.500 ;
        RECT 50.585 20.455 50.875 20.500 ;
        RECT 51.665 20.480 51.955 20.795 ;
        RECT 53.430 20.780 53.750 20.840 ;
        RECT 54.365 20.795 54.655 20.840 ;
        RECT 55.445 20.980 55.735 21.025 ;
        RECT 57.570 20.980 57.890 21.040 ;
        RECT 55.445 20.840 57.890 20.980 ;
        RECT 55.445 20.795 55.735 20.840 ;
        RECT 57.570 20.780 57.890 20.840 ;
        RECT 58.030 20.780 58.350 21.040 ;
        RECT 65.965 20.980 66.255 21.025 ;
        RECT 68.150 20.980 68.470 21.040 ;
        RECT 69.205 20.980 69.855 21.025 ;
        RECT 65.965 20.840 69.855 20.980 ;
        RECT 65.965 20.795 66.555 20.840 ;
        RECT 58.950 20.640 59.270 20.700 ;
        RECT 61.850 20.640 62.140 20.685 ;
        RECT 58.950 20.500 62.140 20.640 ;
        RECT 58.950 20.440 59.270 20.500 ;
        RECT 61.850 20.455 62.140 20.500 ;
        RECT 66.265 20.480 66.555 20.795 ;
        RECT 68.150 20.780 68.470 20.840 ;
        RECT 69.205 20.795 69.855 20.840 ;
        RECT 67.345 20.640 67.635 20.685 ;
        RECT 70.925 20.640 71.215 20.685 ;
        RECT 72.760 20.640 73.050 20.685 ;
        RECT 67.345 20.500 73.050 20.640 ;
        RECT 67.345 20.455 67.635 20.500 ;
        RECT 70.925 20.455 71.215 20.500 ;
        RECT 72.760 20.455 73.050 20.500 ;
        RECT 46.085 20.300 46.375 20.345 ;
        RECT 48.370 20.300 48.690 20.360 ;
        RECT 46.085 20.160 48.690 20.300 ;
        RECT 46.085 20.115 46.375 20.160 ;
        RECT 48.370 20.100 48.690 20.160 ;
        RECT 53.445 20.300 53.735 20.345 ;
        RECT 53.890 20.300 54.210 20.360 ;
        RECT 53.445 20.160 54.210 20.300 ;
        RECT 53.445 20.115 53.735 20.160 ;
        RECT 53.890 20.100 54.210 20.160 ;
        RECT 58.490 20.300 58.810 20.360 ;
        RECT 59.425 20.300 59.715 20.345 ;
        RECT 58.490 20.160 59.715 20.300 ;
        RECT 58.490 20.100 58.810 20.160 ;
        RECT 59.425 20.115 59.715 20.160 ;
        RECT 59.870 20.300 60.190 20.360 ;
        RECT 60.805 20.300 61.095 20.345 ;
        RECT 59.870 20.160 61.095 20.300 ;
        RECT 45.575 19.960 45.865 20.005 ;
        RECT 47.465 19.960 47.755 20.005 ;
        RECT 50.585 19.960 50.875 20.005 ;
        RECT 56.650 19.960 56.970 20.020 ;
        RECT 45.575 19.820 50.875 19.960 ;
        RECT 45.575 19.775 45.865 19.820 ;
        RECT 47.465 19.775 47.755 19.820 ;
        RECT 50.585 19.775 50.875 19.820 ;
        RECT 55.360 19.820 56.970 19.960 ;
        RECT 59.500 19.960 59.640 20.115 ;
        RECT 59.870 20.100 60.190 20.160 ;
        RECT 60.805 20.115 61.095 20.160 ;
        RECT 63.105 20.115 63.395 20.345 ;
        RECT 63.180 19.960 63.320 20.115 ;
        RECT 71.830 20.100 72.150 20.360 ;
        RECT 73.225 20.300 73.515 20.345 ;
        RECT 72.840 20.160 73.515 20.300 ;
        RECT 59.500 19.820 63.320 19.960 ;
        RECT 67.345 19.960 67.635 20.005 ;
        RECT 70.465 19.960 70.755 20.005 ;
        RECT 72.355 19.960 72.645 20.005 ;
        RECT 67.345 19.820 72.645 19.960 ;
        RECT 55.360 19.665 55.500 19.820 ;
        RECT 56.650 19.760 56.970 19.820 ;
        RECT 67.345 19.775 67.635 19.820 ;
        RECT 70.465 19.775 70.755 19.820 ;
        RECT 72.355 19.775 72.645 19.820 ;
        RECT 55.285 19.435 55.575 19.665 ;
        RECT 62.645 19.620 62.935 19.665 ;
        RECT 66.310 19.620 66.630 19.680 ;
        RECT 62.645 19.480 66.630 19.620 ;
        RECT 62.645 19.435 62.935 19.480 ;
        RECT 66.310 19.420 66.630 19.480 ;
        RECT 69.070 19.620 69.390 19.680 ;
        RECT 72.840 19.620 72.980 20.160 ;
        RECT 73.225 20.115 73.515 20.160 ;
        RECT 69.070 19.480 72.980 19.620 ;
        RECT 69.070 19.420 69.390 19.480 ;
        RECT 5.520 18.800 118.680 19.280 ;
        RECT 55.285 18.600 55.575 18.645 ;
        RECT 58.950 18.600 59.270 18.660 ;
        RECT 55.285 18.460 59.270 18.600 ;
        RECT 55.285 18.415 55.575 18.460 ;
        RECT 58.950 18.400 59.270 18.460 ;
        RECT 59.870 18.600 60.190 18.660 ;
        RECT 64.485 18.600 64.775 18.645 ;
        RECT 59.870 18.460 64.775 18.600 ;
        RECT 59.870 18.400 60.190 18.460 ;
        RECT 64.485 18.415 64.775 18.460 ;
        RECT 67.705 18.600 67.995 18.645 ;
        RECT 68.150 18.600 68.470 18.660 ;
        RECT 67.705 18.460 68.470 18.600 ;
        RECT 67.705 18.415 67.995 18.460 ;
        RECT 68.150 18.400 68.470 18.460 ;
        RECT 47.415 18.260 47.705 18.305 ;
        RECT 49.305 18.260 49.595 18.305 ;
        RECT 52.425 18.260 52.715 18.305 ;
        RECT 47.415 18.120 52.715 18.260 ;
        RECT 47.415 18.075 47.705 18.120 ;
        RECT 49.305 18.075 49.595 18.120 ;
        RECT 52.425 18.075 52.715 18.120 ;
        RECT 56.615 18.260 56.905 18.305 ;
        RECT 58.505 18.260 58.795 18.305 ;
        RECT 61.625 18.260 61.915 18.305 ;
        RECT 56.615 18.120 61.915 18.260 ;
        RECT 56.615 18.075 56.905 18.120 ;
        RECT 58.505 18.075 58.795 18.120 ;
        RECT 61.625 18.075 61.915 18.120 ;
        RECT 44.690 17.920 45.010 17.980 ;
        RECT 46.545 17.920 46.835 17.965 ;
        RECT 44.690 17.780 46.835 17.920 ;
        RECT 44.690 17.720 45.010 17.780 ;
        RECT 46.545 17.735 46.835 17.780 ;
        RECT 55.745 17.920 56.035 17.965 ;
        RECT 69.070 17.920 69.390 17.980 ;
        RECT 55.745 17.780 69.390 17.920 ;
        RECT 55.745 17.735 56.035 17.780 ;
        RECT 69.070 17.720 69.390 17.780 ;
        RECT 47.010 17.580 47.300 17.625 ;
        RECT 48.845 17.580 49.135 17.625 ;
        RECT 52.425 17.580 52.715 17.625 ;
        RECT 47.010 17.440 52.715 17.580 ;
        RECT 47.010 17.395 47.300 17.440 ;
        RECT 48.845 17.395 49.135 17.440 ;
        RECT 52.425 17.395 52.715 17.440 ;
        RECT 47.925 17.240 48.215 17.285 ;
        RECT 49.290 17.240 49.610 17.300 ;
        RECT 53.505 17.285 53.795 17.600 ;
        RECT 56.210 17.580 56.500 17.625 ;
        RECT 58.045 17.580 58.335 17.625 ;
        RECT 61.625 17.580 61.915 17.625 ;
        RECT 56.210 17.440 61.915 17.580 ;
        RECT 56.210 17.395 56.500 17.440 ;
        RECT 58.045 17.395 58.335 17.440 ;
        RECT 61.625 17.395 61.915 17.440 ;
        RECT 47.925 17.100 49.610 17.240 ;
        RECT 47.925 17.055 48.215 17.100 ;
        RECT 49.290 17.040 49.610 17.100 ;
        RECT 50.205 17.240 50.855 17.285 ;
        RECT 53.505 17.240 54.095 17.285 ;
        RECT 50.205 17.100 56.880 17.240 ;
        RECT 50.205 17.055 50.855 17.100 ;
        RECT 53.805 17.055 54.095 17.100 ;
        RECT 56.740 16.900 56.880 17.100 ;
        RECT 57.110 17.040 57.430 17.300 ;
        RECT 62.705 17.285 62.995 17.600 ;
        RECT 65.865 17.580 66.155 17.625 ;
        RECT 66.770 17.580 67.090 17.640 ;
        RECT 67.245 17.580 67.535 17.625 ;
        RECT 65.865 17.440 67.535 17.580 ;
        RECT 65.865 17.395 66.155 17.440 ;
        RECT 66.770 17.380 67.090 17.440 ;
        RECT 67.245 17.395 67.535 17.440 ;
        RECT 59.405 17.240 60.055 17.285 ;
        RECT 62.705 17.240 63.295 17.285 ;
        RECT 65.405 17.240 65.695 17.285 ;
        RECT 59.405 17.100 65.695 17.240 ;
        RECT 59.405 17.055 60.055 17.100 ;
        RECT 63.005 17.055 63.295 17.100 ;
        RECT 65.405 17.055 65.695 17.100 ;
        RECT 58.950 16.900 59.270 16.960 ;
        RECT 56.740 16.760 59.270 16.900 ;
        RECT 58.950 16.700 59.270 16.760 ;
        RECT 5.520 16.080 118.680 16.560 ;
        RECT 55.745 15.880 56.035 15.925 ;
        RECT 57.110 15.880 57.430 15.940 ;
        RECT 55.745 15.740 57.430 15.880 ;
        RECT 55.745 15.695 56.035 15.740 ;
        RECT 57.110 15.680 57.430 15.740 ;
        RECT 58.950 15.880 59.270 15.940 ;
        RECT 59.885 15.880 60.175 15.925 ;
        RECT 58.950 15.740 60.175 15.880 ;
        RECT 58.950 15.680 59.270 15.740 ;
        RECT 59.885 15.695 60.175 15.740 ;
        RECT 53.905 15.015 54.195 15.245 ;
        RECT 58.965 15.200 59.255 15.245 ;
        RECT 59.870 15.200 60.190 15.260 ;
        RECT 58.965 15.060 60.190 15.200 ;
        RECT 58.965 15.015 59.255 15.060 ;
        RECT 53.430 14.660 53.750 14.920 ;
        RECT 53.980 14.520 54.120 15.015 ;
        RECT 59.870 15.000 60.190 15.060 ;
        RECT 60.345 15.200 60.635 15.245 ;
        RECT 66.770 15.200 67.090 15.260 ;
        RECT 60.345 15.060 67.090 15.200 ;
        RECT 60.345 15.015 60.635 15.060 ;
        RECT 66.770 15.000 67.090 15.060 ;
        RECT 58.045 14.520 58.335 14.565 ;
        RECT 59.410 14.520 59.730 14.580 ;
        RECT 53.980 14.380 59.730 14.520 ;
        RECT 58.045 14.335 58.335 14.380 ;
        RECT 59.410 14.320 59.730 14.380 ;
        RECT 5.520 13.360 118.680 13.840 ;
        RECT 5.520 10.640 118.680 11.120 ;
      LAYER met2 ;
        RECT 39.260 133.550 41.030 133.690 ;
        RECT 46.160 133.550 47.010 133.690 ;
        RECT 77.190 133.550 78.500 133.690 ;
        RECT 5.220 113.550 5.360 133.000 ;
        RECT 11.200 123.490 11.340 133.000 ;
        RECT 11.200 123.350 12.260 123.490 ;
        RECT 9.580 122.215 11.460 122.585 ;
        RECT 7.000 118.330 7.260 118.650 ;
        RECT 7.060 116.125 7.200 118.330 ;
        RECT 9.580 116.775 11.460 117.145 ;
        RECT 6.990 115.755 7.270 116.125 ;
        RECT 12.120 115.930 12.260 123.350 ;
        RECT 13.440 120.710 13.700 121.030 ;
        RECT 12.980 120.030 13.240 120.350 ;
        RECT 12.060 115.610 12.320 115.930 ;
        RECT 13.040 115.250 13.180 120.030 ;
        RECT 12.980 114.930 13.240 115.250 ;
        RECT 13.500 113.800 13.640 120.710 ;
        RECT 16.660 118.670 16.920 118.990 ;
        RECT 15.740 114.930 16.000 115.250 ;
        RECT 13.900 113.800 14.160 113.890 ;
        RECT 13.500 113.660 14.160 113.800 ;
        RECT 5.160 113.230 5.420 113.550 ;
        RECT 12.980 113.230 13.240 113.550 ;
        RECT 9.580 111.335 11.460 111.705 ;
        RECT 13.040 110.490 13.180 113.230 ;
        RECT 12.980 110.170 13.240 110.490 ;
        RECT 13.500 110.150 13.640 113.660 ;
        RECT 13.900 113.570 14.160 113.660 ;
        RECT 13.900 112.550 14.160 112.870 ;
        RECT 11.140 109.830 11.400 110.150 ;
        RECT 13.440 109.830 13.700 110.150 ;
        RECT 11.200 108.450 11.340 109.830 ;
        RECT 13.960 109.810 14.100 112.550 ;
        RECT 13.900 109.490 14.160 109.810 ;
        RECT 15.800 109.470 15.940 114.930 ;
        RECT 16.720 113.890 16.860 118.670 ;
        RECT 17.180 118.310 17.320 133.000 ;
        RECT 23.160 124.170 23.300 133.000 ;
        RECT 23.160 124.030 24.220 124.170 ;
        RECT 17.120 117.990 17.380 118.310 ;
        RECT 18.960 117.990 19.220 118.310 ;
        RECT 20.800 117.990 21.060 118.310 ;
        RECT 22.180 117.990 22.440 118.310 ;
        RECT 19.020 113.890 19.160 117.990 ;
        RECT 20.860 115.930 21.000 117.990 ;
        RECT 20.800 115.610 21.060 115.930 ;
        RECT 20.860 115.330 21.000 115.610 ;
        RECT 20.860 115.190 21.460 115.330 ;
        RECT 16.660 113.570 16.920 113.890 ;
        RECT 18.960 113.570 19.220 113.890 ;
        RECT 21.320 112.530 21.460 115.190 ;
        RECT 21.720 114.930 21.980 115.250 ;
        RECT 21.780 113.890 21.920 114.930 ;
        RECT 21.720 113.570 21.980 113.890 ;
        RECT 21.720 112.890 21.980 113.210 ;
        RECT 21.260 112.210 21.520 112.530 ;
        RECT 21.320 109.470 21.460 112.210 ;
        RECT 15.740 109.150 16.000 109.470 ;
        RECT 21.260 109.150 21.520 109.470 ;
        RECT 11.140 108.130 11.400 108.450 ;
        RECT 20.340 107.110 20.600 107.430 ;
        RECT 19.880 106.770 20.140 107.090 ;
        RECT 17.580 106.430 17.840 106.750 ;
        RECT 9.580 105.895 11.460 106.265 ;
        RECT 17.640 104.710 17.780 106.430 ;
        RECT 17.580 104.390 17.840 104.710 ;
        RECT 14.820 104.050 15.080 104.370 ;
        RECT 12.520 102.010 12.780 102.330 ;
        RECT 14.360 102.240 14.620 102.330 ;
        RECT 14.880 102.240 15.020 104.050 ;
        RECT 16.660 103.710 16.920 104.030 ;
        RECT 19.420 103.710 19.680 104.030 ;
        RECT 16.720 102.330 16.860 103.710 ;
        RECT 19.480 102.670 19.620 103.710 ;
        RECT 19.420 102.350 19.680 102.670 ;
        RECT 14.360 102.100 15.020 102.240 ;
        RECT 14.360 102.010 14.620 102.100 ;
        RECT 11.600 100.990 11.860 101.310 ;
        RECT 9.580 100.455 11.460 100.825 ;
        RECT 11.660 99.610 11.800 100.990 ;
        RECT 12.580 100.290 12.720 102.010 ;
        RECT 13.900 100.990 14.160 101.310 ;
        RECT 12.520 99.970 12.780 100.290 ;
        RECT 11.600 99.290 11.860 99.610 ;
        RECT 8.380 98.950 8.640 99.270 ;
        RECT 8.440 96.890 8.580 98.950 ;
        RECT 13.960 98.930 14.100 100.990 ;
        RECT 13.900 98.610 14.160 98.930 ;
        RECT 14.360 96.910 14.620 97.230 ;
        RECT 8.380 96.570 8.640 96.890 ;
        RECT 8.440 83.970 8.580 96.570 ;
        RECT 12.520 96.230 12.780 96.550 ;
        RECT 9.580 95.015 11.460 95.385 ;
        RECT 12.580 94.850 12.720 96.230 ;
        RECT 14.420 94.850 14.560 96.910 ;
        RECT 12.520 94.530 12.780 94.850 ;
        RECT 14.360 94.530 14.620 94.850 ;
        RECT 14.880 93.830 15.020 102.100 ;
        RECT 16.660 102.010 16.920 102.330 ;
        RECT 19.420 99.520 19.680 99.610 ;
        RECT 19.940 99.520 20.080 106.770 ;
        RECT 19.420 99.380 20.080 99.520 ;
        RECT 19.420 99.290 19.680 99.380 ;
        RECT 19.480 96.550 19.620 99.290 ;
        RECT 20.400 99.270 20.540 107.110 ;
        RECT 21.320 104.710 21.460 109.150 ;
        RECT 21.260 104.390 21.520 104.710 ;
        RECT 21.320 103.010 21.460 104.390 ;
        RECT 21.260 102.690 21.520 103.010 ;
        RECT 20.340 98.950 20.600 99.270 ;
        RECT 19.880 98.610 20.140 98.930 ;
        RECT 19.940 97.570 20.080 98.610 ;
        RECT 19.880 97.250 20.140 97.570 ;
        RECT 19.420 96.230 19.680 96.550 ;
        RECT 18.040 95.550 18.300 95.870 ;
        RECT 18.100 94.170 18.240 95.550 ;
        RECT 18.040 93.850 18.300 94.170 ;
        RECT 19.940 93.830 20.080 97.250 ;
        RECT 20.400 96.800 20.540 98.950 ;
        RECT 20.400 96.660 21.000 96.800 ;
        RECT 14.820 93.510 15.080 93.830 ;
        RECT 19.880 93.510 20.140 93.830 ;
        RECT 14.880 90.770 15.020 93.510 ;
        RECT 20.860 91.450 21.000 96.660 ;
        RECT 21.780 93.570 21.920 112.890 ;
        RECT 22.240 112.530 22.380 117.990 ;
        RECT 23.560 114.930 23.820 115.250 ;
        RECT 23.620 113.890 23.760 114.930 ;
        RECT 24.080 114.910 24.220 124.030 ;
        RECT 24.580 119.495 26.460 119.865 ;
        RECT 29.140 118.990 29.280 133.000 ;
        RECT 35.120 121.370 35.260 133.000 ;
        RECT 33.680 121.050 33.940 121.370 ;
        RECT 35.060 121.050 35.320 121.370 ;
        RECT 33.220 120.370 33.480 120.690 ;
        RECT 28.620 118.670 28.880 118.990 ;
        RECT 29.080 118.670 29.340 118.990 ;
        RECT 28.680 116.610 28.820 118.670 ;
        RECT 28.620 116.290 28.880 116.610 ;
        RECT 30.460 115.270 30.720 115.590 ;
        RECT 24.020 114.590 24.280 114.910 ;
        RECT 24.580 114.055 26.460 114.425 ;
        RECT 23.560 113.570 23.820 113.890 ;
        RECT 30.520 113.550 30.660 115.270 ;
        RECT 33.280 113.890 33.420 120.370 ;
        RECT 33.740 118.310 33.880 121.050 ;
        RECT 35.520 120.370 35.780 120.690 ;
        RECT 33.680 117.990 33.940 118.310 ;
        RECT 33.740 115.930 33.880 117.990 ;
        RECT 35.580 116.610 35.720 120.370 ;
        RECT 35.520 116.290 35.780 116.610 ;
        RECT 33.680 115.610 33.940 115.930 ;
        RECT 35.060 114.930 35.320 115.250 ;
        RECT 35.120 113.890 35.260 114.930 ;
        RECT 39.260 114.910 39.400 133.550 ;
        RECT 39.580 122.215 41.460 122.585 ;
        RECT 46.160 118.990 46.300 133.550 ;
        RECT 45.180 118.670 45.440 118.990 ;
        RECT 46.100 118.670 46.360 118.990 ;
        RECT 44.720 117.990 44.980 118.310 ;
        RECT 39.580 116.775 41.460 117.145 ;
        RECT 44.780 116.610 44.920 117.990 ;
        RECT 44.720 116.290 44.980 116.610 ;
        RECT 40.120 114.930 40.380 115.250 ;
        RECT 39.200 114.590 39.460 114.910 ;
        RECT 40.180 113.890 40.320 114.930 ;
        RECT 45.240 113.890 45.380 118.670 ;
        RECT 46.560 117.990 46.820 118.310 ;
        RECT 46.620 115.930 46.760 117.990 ;
        RECT 53.060 115.930 53.200 133.000 ;
        RECT 54.580 119.495 56.460 119.865 ;
        RECT 59.040 118.990 59.180 133.000 ;
        RECT 58.980 118.670 59.240 118.990 ;
        RECT 53.460 118.330 53.720 118.650 ;
        RECT 46.560 115.610 46.820 115.930 ;
        RECT 53.000 115.610 53.260 115.930 ;
        RECT 46.100 115.270 46.360 115.590 ;
        RECT 33.220 113.570 33.480 113.890 ;
        RECT 35.060 113.570 35.320 113.890 ;
        RECT 40.120 113.570 40.380 113.890 ;
        RECT 45.180 113.570 45.440 113.890 ;
        RECT 30.460 113.230 30.720 113.550 ;
        RECT 22.640 112.890 22.900 113.210 ;
        RECT 29.540 112.890 29.800 113.210 ;
        RECT 33.220 112.890 33.480 113.210 ;
        RECT 38.280 112.890 38.540 113.210 ;
        RECT 22.180 112.210 22.440 112.530 ;
        RECT 21.320 93.430 21.920 93.570 ;
        RECT 22.180 93.510 22.440 93.830 ;
        RECT 20.800 91.130 21.060 91.450 ;
        RECT 14.820 90.450 15.080 90.770 ;
        RECT 9.580 89.575 11.460 89.945 ;
        RECT 12.060 87.390 12.320 87.710 ;
        RECT 12.120 86.010 12.260 87.390 ;
        RECT 12.060 85.690 12.320 86.010 ;
        RECT 11.600 85.350 11.860 85.670 ;
        RECT 8.840 84.670 9.100 84.990 ;
        RECT 8.380 83.650 8.640 83.970 ;
        RECT 7.000 82.970 7.260 83.290 ;
        RECT 7.060 75.130 7.200 82.970 ;
        RECT 8.900 82.950 9.040 84.670 ;
        RECT 9.580 84.135 11.460 84.505 ;
        RECT 11.660 83.970 11.800 85.350 ;
        RECT 13.440 84.670 13.700 84.990 ;
        RECT 11.600 83.650 11.860 83.970 ;
        RECT 12.980 83.310 13.240 83.630 ;
        RECT 8.840 82.630 9.100 82.950 ;
        RECT 12.520 82.290 12.780 82.610 ;
        RECT 12.580 81.250 12.720 82.290 ;
        RECT 12.520 80.930 12.780 81.250 ;
        RECT 13.040 80.650 13.180 83.310 ;
        RECT 13.500 81.250 13.640 84.670 ;
        RECT 13.440 80.930 13.700 81.250 ;
        RECT 13.040 80.570 13.640 80.650 ;
        RECT 13.040 80.510 13.700 80.570 ;
        RECT 13.440 80.250 13.700 80.510 ;
        RECT 9.580 78.695 11.460 79.065 ;
        RECT 13.500 77.510 13.640 80.250 ;
        RECT 13.440 77.190 13.700 77.510 ;
        RECT 9.300 76.510 9.560 76.830 ;
        RECT 12.980 76.510 13.240 76.830 ;
        RECT 9.360 75.130 9.500 76.510 ;
        RECT 13.040 75.470 13.180 76.510 ;
        RECT 12.980 75.150 13.240 75.470 ;
        RECT 7.000 74.810 7.260 75.130 ;
        RECT 9.300 74.810 9.560 75.130 ;
        RECT 7.060 72.410 7.200 74.810 ;
        RECT 9.580 73.255 11.460 73.625 ;
        RECT 7.000 72.090 7.260 72.410 ;
        RECT 9.760 71.410 10.020 71.730 ;
        RECT 9.820 70.370 9.960 71.410 ;
        RECT 9.760 70.050 10.020 70.370 ;
        RECT 13.500 69.690 13.640 77.190 ;
        RECT 14.880 74.700 15.020 90.450 ;
        RECT 19.880 88.070 20.140 88.390 ;
        RECT 19.940 86.690 20.080 88.070 ;
        RECT 20.800 87.730 21.060 88.050 ;
        RECT 19.880 86.370 20.140 86.690 ;
        RECT 17.120 86.030 17.380 86.350 ;
        RECT 17.180 82.950 17.320 86.030 ;
        RECT 20.340 85.690 20.600 86.010 ;
        RECT 19.880 85.010 20.140 85.330 ;
        RECT 17.120 82.630 17.380 82.950 ;
        RECT 15.740 82.290 16.000 82.610 ;
        RECT 15.800 81.250 15.940 82.290 ;
        RECT 15.740 80.930 16.000 81.250 ;
        RECT 15.280 80.250 15.540 80.570 ;
        RECT 15.340 77.850 15.480 80.250 ;
        RECT 19.940 80.230 20.080 85.010 ;
        RECT 20.400 83.630 20.540 85.690 ;
        RECT 20.340 83.310 20.600 83.630 ;
        RECT 20.340 82.630 20.600 82.950 ;
        RECT 19.880 79.910 20.140 80.230 ;
        RECT 15.280 77.530 15.540 77.850 ;
        RECT 19.420 77.760 19.680 77.850 ;
        RECT 19.940 77.760 20.080 79.910 ;
        RECT 20.400 78.610 20.540 82.630 ;
        RECT 20.860 82.610 21.000 87.730 ;
        RECT 20.800 82.290 21.060 82.610 ;
        RECT 21.320 79.550 21.460 93.430 ;
        RECT 21.720 92.830 21.980 93.150 ;
        RECT 21.780 89.410 21.920 92.830 ;
        RECT 22.240 91.450 22.380 93.510 ;
        RECT 22.180 91.130 22.440 91.450 ;
        RECT 22.700 89.410 22.840 112.890 ;
        RECT 28.620 110.170 28.880 110.490 ;
        RECT 24.580 108.615 26.460 108.985 ;
        RECT 23.560 107.450 23.820 107.770 ;
        RECT 24.020 107.450 24.280 107.770 ;
        RECT 23.100 106.430 23.360 106.750 ;
        RECT 23.160 104.710 23.300 106.430 ;
        RECT 23.100 104.390 23.360 104.710 ;
        RECT 23.620 101.990 23.760 107.450 ;
        RECT 24.080 103.010 24.220 107.450 ;
        RECT 27.240 104.050 27.500 104.370 ;
        RECT 24.580 103.175 26.460 103.545 ;
        RECT 27.300 103.010 27.440 104.050 ;
        RECT 24.020 102.690 24.280 103.010 ;
        RECT 27.240 102.690 27.500 103.010 ;
        RECT 26.780 102.350 27.040 102.670 ;
        RECT 23.560 101.670 23.820 101.990 ;
        RECT 23.620 94.170 23.760 101.670 ;
        RECT 24.580 97.735 26.460 98.105 ;
        RECT 23.560 93.850 23.820 94.170 ;
        RECT 26.840 93.830 26.980 102.350 ;
        RECT 27.700 101.670 27.960 101.990 ;
        RECT 27.760 99.610 27.900 101.670 ;
        RECT 27.700 99.290 27.960 99.610 ;
        RECT 27.700 96.570 27.960 96.890 ;
        RECT 27.760 94.170 27.900 96.570 ;
        RECT 27.700 93.850 27.960 94.170 ;
        RECT 26.780 93.510 27.040 93.830 ;
        RECT 26.780 92.830 27.040 93.150 ;
        RECT 28.160 92.830 28.420 93.150 ;
        RECT 24.580 92.295 26.460 92.665 ;
        RECT 23.100 90.110 23.360 90.430 ;
        RECT 21.720 89.090 21.980 89.410 ;
        RECT 22.640 89.090 22.900 89.410 ;
        RECT 21.720 88.070 21.980 88.390 ;
        RECT 22.180 88.070 22.440 88.390 ;
        RECT 21.260 79.230 21.520 79.550 ;
        RECT 20.400 78.470 21.460 78.610 ;
        RECT 19.420 77.620 20.080 77.760 ;
        RECT 19.420 77.530 19.680 77.620 ;
        RECT 15.340 75.470 15.480 77.530 ;
        RECT 15.740 76.510 16.000 76.830 ;
        RECT 15.800 75.810 15.940 76.510 ;
        RECT 15.740 75.490 16.000 75.810 ;
        RECT 18.960 75.490 19.220 75.810 ;
        RECT 15.280 75.150 15.540 75.470 ;
        RECT 14.880 74.560 15.480 74.700 ;
        RECT 14.820 71.410 15.080 71.730 ;
        RECT 15.340 71.640 15.480 74.560 ;
        RECT 17.120 73.790 17.380 74.110 ;
        RECT 16.200 71.640 16.460 71.730 ;
        RECT 15.340 71.500 16.460 71.640 ;
        RECT 14.880 70.370 15.020 71.410 ;
        RECT 14.820 70.050 15.080 70.370 ;
        RECT 13.440 69.370 13.700 69.690 ;
        RECT 9.580 67.815 11.460 68.185 ;
        RECT 15.340 66.970 15.480 71.500 ;
        RECT 16.200 71.410 16.460 71.500 ;
        RECT 17.180 70.030 17.320 73.790 ;
        RECT 19.020 73.090 19.160 75.490 ;
        RECT 19.940 74.790 20.080 77.620 ;
        RECT 21.320 77.510 21.460 78.470 ;
        RECT 20.340 77.420 20.600 77.510 ;
        RECT 20.340 77.280 21.000 77.420 ;
        RECT 20.340 77.190 20.600 77.280 ;
        RECT 20.860 75.130 21.000 77.280 ;
        RECT 21.260 77.190 21.520 77.510 ;
        RECT 20.800 74.810 21.060 75.130 ;
        RECT 19.880 74.470 20.140 74.790 ;
        RECT 18.960 72.770 19.220 73.090 ;
        RECT 21.320 72.750 21.460 77.190 ;
        RECT 21.260 72.430 21.520 72.750 ;
        RECT 20.800 70.050 21.060 70.370 ;
        RECT 17.120 69.710 17.380 70.030 ;
        RECT 16.660 69.030 16.920 69.350 ;
        RECT 15.280 66.650 15.540 66.970 ;
        RECT 16.200 63.590 16.460 63.910 ;
        RECT 12.060 62.910 12.320 63.230 ;
        RECT 9.580 62.375 11.460 62.745 ;
        RECT 12.120 61.190 12.260 62.910 ;
        RECT 16.260 62.210 16.400 63.590 ;
        RECT 16.200 61.890 16.460 62.210 ;
        RECT 12.060 60.870 12.320 61.190 ;
        RECT 13.900 60.870 14.160 61.190 ;
        RECT 9.300 60.530 9.560 60.850 ;
        RECT 9.360 58.810 9.500 60.530 ;
        RECT 11.600 60.190 11.860 60.510 ;
        RECT 13.440 60.190 13.700 60.510 ;
        RECT 9.300 58.490 9.560 58.810 ;
        RECT 8.380 58.150 8.640 58.470 ;
        RECT 8.440 55.750 8.580 58.150 ;
        RECT 9.580 56.935 11.460 57.305 ;
        RECT 11.660 56.770 11.800 60.190 ;
        RECT 11.600 56.450 11.860 56.770 ;
        RECT 8.380 55.430 8.640 55.750 ;
        RECT 5.160 53.050 5.420 53.370 ;
        RECT 5.220 50.845 5.360 53.050 ;
        RECT 5.150 50.475 5.430 50.845 ;
        RECT 8.440 50.650 8.580 55.430 ;
        RECT 13.500 55.410 13.640 60.190 ;
        RECT 13.440 55.090 13.700 55.410 ;
        RECT 11.600 52.030 11.860 52.350 ;
        RECT 9.580 51.495 11.460 51.865 ;
        RECT 11.660 50.650 11.800 52.030 ;
        RECT 8.380 50.330 8.640 50.650 ;
        RECT 11.600 50.330 11.860 50.650 ;
        RECT 13.960 49.630 14.100 60.870 ;
        RECT 16.720 60.510 16.860 69.030 ;
        RECT 18.500 68.690 18.760 69.010 ;
        RECT 15.740 60.190 16.000 60.510 ;
        RECT 16.660 60.190 16.920 60.510 ;
        RECT 15.800 53.030 15.940 60.190 ;
        RECT 18.560 53.370 18.700 68.690 ;
        RECT 19.880 66.310 20.140 66.630 ;
        RECT 18.960 60.870 19.220 61.190 ;
        RECT 19.020 56.770 19.160 60.870 ;
        RECT 19.420 58.830 19.680 59.150 ;
        RECT 18.960 56.450 19.220 56.770 ;
        RECT 18.500 53.050 18.760 53.370 ;
        RECT 15.740 52.710 16.000 53.030 ;
        RECT 15.800 51.330 15.940 52.710 ;
        RECT 15.740 51.010 16.000 51.330 ;
        RECT 18.560 50.990 18.700 53.050 ;
        RECT 19.480 51.330 19.620 58.830 ;
        RECT 19.940 58.810 20.080 66.310 ;
        RECT 20.860 64.590 21.000 70.050 ;
        RECT 21.260 65.630 21.520 65.950 ;
        RECT 20.800 64.270 21.060 64.590 ;
        RECT 20.860 63.650 21.000 64.270 ;
        RECT 21.320 64.250 21.460 65.630 ;
        RECT 21.260 63.930 21.520 64.250 ;
        RECT 20.860 63.510 21.460 63.650 ;
        RECT 20.800 62.910 21.060 63.230 ;
        RECT 20.340 61.210 20.600 61.530 ;
        RECT 20.400 58.810 20.540 61.210 ;
        RECT 19.880 58.490 20.140 58.810 ;
        RECT 20.340 58.490 20.600 58.810 ;
        RECT 19.940 57.790 20.080 58.490 ;
        RECT 19.880 57.470 20.140 57.790 ;
        RECT 19.940 54.050 20.080 57.470 ;
        RECT 19.880 53.730 20.140 54.050 ;
        RECT 20.400 53.030 20.540 58.490 ;
        RECT 20.860 56.430 21.000 62.910 ;
        RECT 21.320 59.150 21.460 63.510 ;
        RECT 21.260 58.830 21.520 59.150 ;
        RECT 20.800 56.110 21.060 56.430 ;
        RECT 20.860 55.750 21.000 56.110 ;
        RECT 21.260 55.770 21.520 56.090 ;
        RECT 20.800 55.430 21.060 55.750 ;
        RECT 21.320 53.370 21.460 55.770 ;
        RECT 21.260 53.050 21.520 53.370 ;
        RECT 20.340 52.710 20.600 53.030 ;
        RECT 21.780 51.330 21.920 88.070 ;
        RECT 22.240 67.650 22.380 88.070 ;
        RECT 22.640 87.730 22.900 88.050 ;
        RECT 22.700 82.610 22.840 87.730 ;
        RECT 22.640 82.290 22.900 82.610 ;
        RECT 22.700 78.530 22.840 82.290 ;
        RECT 23.160 78.530 23.300 90.110 ;
        RECT 23.560 88.070 23.820 88.390 ;
        RECT 24.020 88.070 24.280 88.390 ;
        RECT 24.940 88.245 25.200 88.390 ;
        RECT 23.620 82.950 23.760 88.070 ;
        RECT 24.080 86.350 24.220 88.070 ;
        RECT 24.930 87.875 25.210 88.245 ;
        RECT 24.580 86.855 26.460 87.225 ;
        RECT 24.020 86.030 24.280 86.350 ;
        RECT 23.560 82.630 23.820 82.950 ;
        RECT 22.640 78.210 22.900 78.530 ;
        RECT 23.100 78.210 23.360 78.530 ;
        RECT 23.620 77.930 23.760 82.630 ;
        RECT 24.580 81.415 26.460 81.785 ;
        RECT 24.020 79.230 24.280 79.550 ;
        RECT 24.080 78.190 24.220 79.230 ;
        RECT 22.640 77.530 22.900 77.850 ;
        RECT 23.160 77.790 23.760 77.930 ;
        RECT 24.020 77.870 24.280 78.190 ;
        RECT 22.180 67.330 22.440 67.650 ;
        RECT 22.180 65.970 22.440 66.290 ;
        RECT 22.240 62.210 22.380 65.970 ;
        RECT 22.180 61.890 22.440 62.210 ;
        RECT 22.700 61.610 22.840 77.530 ;
        RECT 23.160 75.130 23.300 77.790 ;
        RECT 23.560 77.190 23.820 77.510 ;
        RECT 24.020 77.190 24.280 77.510 ;
        RECT 23.620 75.810 23.760 77.190 ;
        RECT 23.560 75.490 23.820 75.810 ;
        RECT 23.100 74.810 23.360 75.130 ;
        RECT 23.160 72.070 23.300 74.810 ;
        RECT 23.100 71.750 23.360 72.070 ;
        RECT 23.560 69.370 23.820 69.690 ;
        RECT 23.100 69.030 23.360 69.350 ;
        RECT 23.160 68.670 23.300 69.030 ;
        RECT 23.100 68.350 23.360 68.670 ;
        RECT 23.160 64.250 23.300 68.350 ;
        RECT 23.620 66.630 23.760 69.370 ;
        RECT 23.560 66.310 23.820 66.630 ;
        RECT 23.620 64.250 23.760 66.310 ;
        RECT 24.080 64.930 24.220 77.190 ;
        RECT 24.580 75.975 26.460 76.345 ;
        RECT 24.940 75.490 25.200 75.810 ;
        RECT 25.000 75.130 25.140 75.490 ;
        RECT 24.940 74.810 25.200 75.130 ;
        RECT 25.000 72.070 25.140 74.810 ;
        RECT 25.400 74.470 25.660 74.790 ;
        RECT 25.460 72.410 25.600 74.470 ;
        RECT 26.840 74.110 26.980 92.830 ;
        RECT 28.220 89.410 28.360 92.830 ;
        RECT 28.160 89.090 28.420 89.410 ;
        RECT 27.700 84.670 27.960 84.990 ;
        RECT 27.760 83.290 27.900 84.670 ;
        RECT 27.700 82.970 27.960 83.290 ;
        RECT 27.700 74.810 27.960 75.130 ;
        RECT 26.780 73.790 27.040 74.110 ;
        RECT 25.400 72.090 25.660 72.410 ;
        RECT 24.940 71.750 25.200 72.070 ;
        RECT 25.460 71.925 25.600 72.090 ;
        RECT 25.390 71.555 25.670 71.925 ;
        RECT 24.580 70.535 26.460 70.905 ;
        RECT 27.760 70.370 27.900 74.810 ;
        RECT 28.680 74.110 28.820 110.170 ;
        RECT 29.600 89.410 29.740 112.890 ;
        RECT 31.380 108.130 31.640 108.450 ;
        RECT 30.460 103.710 30.720 104.030 ;
        RECT 30.520 102.670 30.660 103.710 ;
        RECT 30.460 102.350 30.720 102.670 ;
        RECT 30.000 94.190 30.260 94.510 ;
        RECT 29.540 89.090 29.800 89.410 ;
        RECT 29.080 88.070 29.340 88.390 ;
        RECT 28.620 73.790 28.880 74.110 ;
        RECT 28.160 71.070 28.420 71.390 ;
        RECT 24.480 70.050 24.740 70.370 ;
        RECT 27.700 70.050 27.960 70.370 ;
        RECT 24.540 69.690 24.680 70.050 ;
        RECT 28.220 70.030 28.360 71.070 ;
        RECT 28.160 69.710 28.420 70.030 ;
        RECT 24.480 69.370 24.740 69.690 ;
        RECT 25.400 69.600 25.660 69.690 ;
        RECT 25.000 69.460 25.660 69.600 ;
        RECT 24.540 65.950 24.680 69.370 ;
        RECT 25.000 69.010 25.140 69.460 ;
        RECT 25.400 69.370 25.660 69.460 ;
        RECT 26.320 69.370 26.580 69.690 ;
        RECT 24.940 68.690 25.200 69.010 ;
        RECT 26.380 67.650 26.520 69.370 ;
        RECT 28.620 69.030 28.880 69.350 ;
        RECT 27.700 68.690 27.960 69.010 ;
        RECT 26.320 67.330 26.580 67.650 ;
        RECT 27.760 66.630 27.900 68.690 ;
        RECT 27.700 66.310 27.960 66.630 ;
        RECT 24.480 65.630 24.740 65.950 ;
        RECT 24.580 65.095 26.460 65.465 ;
        RECT 24.020 64.610 24.280 64.930 ;
        RECT 23.100 63.930 23.360 64.250 ;
        RECT 23.560 63.930 23.820 64.250 ;
        RECT 24.020 63.930 24.280 64.250 ;
        RECT 27.700 63.930 27.960 64.250 ;
        RECT 23.560 63.250 23.820 63.570 ;
        RECT 22.240 61.470 22.840 61.610 ;
        RECT 22.240 56.430 22.380 61.470 ;
        RECT 22.640 60.870 22.900 61.190 ;
        RECT 22.700 58.470 22.840 60.870 ;
        RECT 23.100 60.190 23.360 60.510 ;
        RECT 23.160 59.490 23.300 60.190 ;
        RECT 23.100 59.170 23.360 59.490 ;
        RECT 22.640 58.150 22.900 58.470 ;
        RECT 23.620 57.530 23.760 63.250 ;
        RECT 24.080 58.130 24.220 63.930 ;
        RECT 27.240 61.210 27.500 61.530 ;
        RECT 26.780 60.190 27.040 60.510 ;
        RECT 24.580 59.655 26.460 60.025 ;
        RECT 26.840 59.150 26.980 60.190 ;
        RECT 26.780 58.830 27.040 59.150 ;
        RECT 24.020 57.810 24.280 58.130 ;
        RECT 23.160 57.390 23.760 57.530 ;
        RECT 22.180 56.110 22.440 56.430 ;
        RECT 22.180 55.430 22.440 55.750 ;
        RECT 22.240 54.050 22.380 55.430 ;
        RECT 22.640 54.750 22.900 55.070 ;
        RECT 22.180 53.730 22.440 54.050 ;
        RECT 22.700 53.710 22.840 54.750 ;
        RECT 22.640 53.390 22.900 53.710 ;
        RECT 23.160 53.030 23.300 57.390 ;
        RECT 24.020 56.110 24.280 56.430 ;
        RECT 23.100 52.710 23.360 53.030 ;
        RECT 19.420 51.010 19.680 51.330 ;
        RECT 21.720 51.010 21.980 51.330 ;
        RECT 18.500 50.670 18.760 50.990 ;
        RECT 23.100 49.990 23.360 50.310 ;
        RECT 23.560 49.990 23.820 50.310 ;
        RECT 14.820 49.650 15.080 49.970 ;
        RECT 22.640 49.650 22.900 49.970 ;
        RECT 13.900 49.310 14.160 49.630 ;
        RECT 13.960 47.930 14.100 49.310 ;
        RECT 14.880 48.610 15.020 49.650 ;
        RECT 14.820 48.290 15.080 48.610 ;
        RECT 13.900 47.610 14.160 47.930 ;
        RECT 9.580 46.055 11.460 46.425 ;
        RECT 22.180 44.890 22.440 45.210 ;
        RECT 16.200 44.550 16.460 44.870 ;
        RECT 11.140 44.210 11.400 44.530 ;
        RECT 11.200 42.490 11.340 44.210 ;
        RECT 14.360 43.870 14.620 44.190 ;
        RECT 14.420 42.830 14.560 43.870 ;
        RECT 14.820 42.850 15.080 43.170 ;
        RECT 14.360 42.510 14.620 42.830 ;
        RECT 11.140 42.170 11.400 42.490 ;
        RECT 8.380 41.150 8.640 41.470 ;
        RECT 8.440 39.090 8.580 41.150 ;
        RECT 9.580 40.615 11.460 40.985 ;
        RECT 14.880 39.770 15.020 42.850 ;
        RECT 15.280 41.150 15.540 41.470 ;
        RECT 14.820 39.450 15.080 39.770 ;
        RECT 8.380 38.770 8.640 39.090 ;
        RECT 9.580 35.175 11.460 35.545 ;
        RECT 14.880 34.330 15.020 39.450 ;
        RECT 15.340 39.430 15.480 41.150 ;
        RECT 16.260 40.450 16.400 44.550 ;
        RECT 20.800 43.870 21.060 44.190 ;
        RECT 21.260 43.870 21.520 44.190 ;
        RECT 17.120 41.830 17.380 42.150 ;
        RECT 16.200 40.130 16.460 40.450 ;
        RECT 15.280 39.110 15.540 39.430 ;
        RECT 14.820 34.010 15.080 34.330 ;
        RECT 14.880 31.610 15.020 34.010 ;
        RECT 16.660 32.990 16.920 33.310 ;
        RECT 16.720 31.950 16.860 32.990 ;
        RECT 16.660 31.630 16.920 31.950 ;
        RECT 13.900 31.290 14.160 31.610 ;
        RECT 14.820 31.290 15.080 31.610 ;
        RECT 9.580 29.735 11.460 30.105 ;
        RECT 13.960 29.570 14.100 31.290 ;
        RECT 13.900 29.250 14.160 29.570 ;
        RECT 14.880 28.210 15.020 31.290 ;
        RECT 15.280 30.270 15.540 30.590 ;
        RECT 14.820 27.890 15.080 28.210 ;
        RECT 14.880 26.510 15.020 27.890 ;
        RECT 15.340 26.510 15.480 30.270 ;
        RECT 17.180 28.550 17.320 41.830 ;
        RECT 20.860 37.390 21.000 43.870 ;
        RECT 21.320 39.430 21.460 43.870 ;
        RECT 22.240 39.770 22.380 44.890 ;
        RECT 22.700 40.110 22.840 49.650 ;
        RECT 23.160 48.610 23.300 49.990 ;
        RECT 23.100 48.290 23.360 48.610 ;
        RECT 23.620 47.930 23.760 49.990 ;
        RECT 23.100 47.610 23.360 47.930 ;
        RECT 23.560 47.610 23.820 47.930 ;
        RECT 22.640 39.790 22.900 40.110 ;
        RECT 22.180 39.450 22.440 39.770 ;
        RECT 21.260 39.110 21.520 39.430 ;
        RECT 21.320 37.730 21.460 39.110 ;
        RECT 21.260 37.410 21.520 37.730 ;
        RECT 20.800 37.070 21.060 37.390 ;
        RECT 19.880 33.670 20.140 33.990 ;
        RECT 19.940 32.290 20.080 33.670 ;
        RECT 19.880 31.970 20.140 32.290 ;
        RECT 20.340 30.270 20.600 30.590 ;
        RECT 17.120 28.230 17.380 28.550 ;
        RECT 20.400 27.870 20.540 30.270 ;
        RECT 20.860 29.230 21.000 37.070 ;
        RECT 20.800 28.910 21.060 29.230 ;
        RECT 22.240 28.890 22.380 39.450 ;
        RECT 22.700 37.050 22.840 39.790 ;
        RECT 22.640 36.730 22.900 37.050 ;
        RECT 23.160 33.990 23.300 47.610 ;
        RECT 24.080 47.250 24.220 56.110 ;
        RECT 27.300 56.090 27.440 61.210 ;
        RECT 27.760 59.490 27.900 63.930 ;
        RECT 28.160 62.910 28.420 63.230 ;
        RECT 27.700 59.170 27.960 59.490 ;
        RECT 28.220 56.090 28.360 62.910 ;
        RECT 27.240 55.770 27.500 56.090 ;
        RECT 28.160 55.770 28.420 56.090 ;
        RECT 24.580 54.215 26.460 54.585 ;
        RECT 25.860 53.390 26.120 53.710 ;
        RECT 25.920 51.330 26.060 53.390 ;
        RECT 25.860 51.010 26.120 51.330 ;
        RECT 27.300 50.650 27.440 55.770 ;
        RECT 27.240 50.330 27.500 50.650 ;
        RECT 26.780 49.650 27.040 49.970 ;
        RECT 24.580 48.775 26.460 49.145 ;
        RECT 26.320 47.270 26.580 47.590 ;
        RECT 24.020 46.930 24.280 47.250 ;
        RECT 24.940 46.590 25.200 46.910 ;
        RECT 25.000 44.870 25.140 46.590 ;
        RECT 26.380 44.870 26.520 47.270 ;
        RECT 26.840 46.910 26.980 49.650 ;
        RECT 28.680 48.270 28.820 69.030 ;
        RECT 29.140 67.650 29.280 88.070 ;
        RECT 30.060 75.210 30.200 94.190 ;
        RECT 30.460 90.450 30.720 90.770 ;
        RECT 30.520 88.390 30.660 90.450 ;
        RECT 30.920 88.410 31.180 88.730 ;
        RECT 30.460 88.070 30.720 88.390 ;
        RECT 30.460 87.390 30.720 87.710 ;
        RECT 30.520 82.610 30.660 87.390 ;
        RECT 30.460 82.290 30.720 82.610 ;
        RECT 30.060 75.070 30.660 75.210 ;
        RECT 30.000 74.470 30.260 74.790 ;
        RECT 29.540 73.790 29.800 74.110 ;
        RECT 29.600 71.730 29.740 73.790 ;
        RECT 29.540 71.410 29.800 71.730 ;
        RECT 30.060 71.130 30.200 74.470 ;
        RECT 29.600 70.990 30.200 71.130 ;
        RECT 29.080 67.330 29.340 67.650 ;
        RECT 28.620 47.950 28.880 48.270 ;
        RECT 27.240 47.610 27.500 47.930 ;
        RECT 28.160 47.840 28.420 47.930 ;
        RECT 27.760 47.700 28.420 47.840 ;
        RECT 26.780 46.590 27.040 46.910 ;
        RECT 27.300 45.210 27.440 47.610 ;
        RECT 27.240 44.890 27.500 45.210 ;
        RECT 23.560 44.550 23.820 44.870 ;
        RECT 24.940 44.550 25.200 44.870 ;
        RECT 26.320 44.780 26.580 44.870 ;
        RECT 26.320 44.640 26.980 44.780 ;
        RECT 26.320 44.550 26.580 44.640 ;
        RECT 23.620 39.430 23.760 44.550 ;
        RECT 24.020 44.210 24.280 44.530 ;
        RECT 24.080 42.490 24.220 44.210 ;
        RECT 24.580 43.335 26.460 43.705 ;
        RECT 24.020 42.170 24.280 42.490 ;
        RECT 24.940 41.830 25.200 42.150 ;
        RECT 25.000 39.430 25.140 41.830 ;
        RECT 26.840 39.430 26.980 44.640 ;
        RECT 27.300 42.150 27.440 44.890 ;
        RECT 27.240 41.830 27.500 42.150 ;
        RECT 27.240 41.150 27.500 41.470 ;
        RECT 27.300 39.430 27.440 41.150 ;
        RECT 23.560 39.110 23.820 39.430 ;
        RECT 24.940 39.110 25.200 39.430 ;
        RECT 26.780 39.110 27.040 39.430 ;
        RECT 27.240 39.110 27.500 39.430 ;
        RECT 27.240 38.430 27.500 38.750 ;
        RECT 24.580 37.895 26.460 38.265 ;
        RECT 27.300 37.050 27.440 38.430 ;
        RECT 27.240 36.730 27.500 37.050 ;
        RECT 27.760 36.710 27.900 47.700 ;
        RECT 28.160 47.610 28.420 47.700 ;
        RECT 28.160 41.830 28.420 42.150 ;
        RECT 28.220 40.450 28.360 41.830 ;
        RECT 28.160 40.130 28.420 40.450 ;
        RECT 29.600 39.850 29.740 70.990 ;
        RECT 30.000 68.580 30.260 68.670 ;
        RECT 30.520 68.580 30.660 75.070 ;
        RECT 30.000 68.440 30.660 68.580 ;
        RECT 30.000 68.350 30.260 68.440 ;
        RECT 30.460 66.990 30.720 67.310 ;
        RECT 30.000 65.970 30.260 66.290 ;
        RECT 30.060 62.170 30.200 65.970 ;
        RECT 30.520 65.950 30.660 66.990 ;
        RECT 30.460 65.630 30.720 65.950 ;
        RECT 30.060 62.030 30.660 62.170 ;
        RECT 30.520 61.190 30.660 62.030 ;
        RECT 30.460 60.870 30.720 61.190 ;
        RECT 30.520 54.050 30.660 60.870 ;
        RECT 30.460 53.730 30.720 54.050 ;
        RECT 30.980 45.890 31.120 88.410 ;
        RECT 31.440 70.370 31.580 108.130 ;
        RECT 31.840 107.450 32.100 107.770 ;
        RECT 31.900 103.010 32.040 107.450 ;
        RECT 32.760 106.430 33.020 106.750 ;
        RECT 32.820 105.050 32.960 106.430 ;
        RECT 32.760 104.730 33.020 105.050 ;
        RECT 31.840 102.690 32.100 103.010 ;
        RECT 32.760 102.010 33.020 102.330 ;
        RECT 32.820 99.270 32.960 102.010 ;
        RECT 32.760 98.950 33.020 99.270 ;
        RECT 31.840 96.570 32.100 96.890 ;
        RECT 32.760 96.570 33.020 96.890 ;
        RECT 31.900 89.410 32.040 96.570 ;
        RECT 32.820 93.830 32.960 96.570 ;
        RECT 32.760 93.510 33.020 93.830 ;
        RECT 32.820 90.770 32.960 93.510 ;
        RECT 32.760 90.450 33.020 90.770 ;
        RECT 33.280 89.410 33.420 112.890 ;
        RECT 33.680 102.010 33.940 102.330 ;
        RECT 33.740 96.890 33.880 102.010 ;
        RECT 33.680 96.570 33.940 96.890 ;
        RECT 34.600 96.230 34.860 96.550 ;
        RECT 34.140 95.550 34.400 95.870 ;
        RECT 34.200 94.170 34.340 95.550 ;
        RECT 34.140 93.850 34.400 94.170 ;
        RECT 34.660 93.150 34.800 96.230 ;
        RECT 37.360 93.170 37.620 93.490 ;
        RECT 34.600 92.830 34.860 93.150 ;
        RECT 37.420 93.005 37.560 93.170 ;
        RECT 34.660 91.450 34.800 92.830 ;
        RECT 37.350 92.635 37.630 93.005 ;
        RECT 37.820 92.830 38.080 93.150 ;
        RECT 34.600 91.130 34.860 91.450 ;
        RECT 31.840 89.090 32.100 89.410 ;
        RECT 33.220 89.090 33.480 89.410 ;
        RECT 32.300 88.410 32.560 88.730 ;
        RECT 31.840 87.730 32.100 88.050 ;
        RECT 31.900 86.690 32.040 87.730 ;
        RECT 31.840 86.370 32.100 86.690 ;
        RECT 31.380 70.050 31.640 70.370 ;
        RECT 31.840 58.490 32.100 58.810 ;
        RECT 31.900 58.325 32.040 58.490 ;
        RECT 31.830 57.955 32.110 58.325 ;
        RECT 32.360 45.890 32.500 88.410 ;
        RECT 34.660 88.390 34.800 91.130 ;
        RECT 37.880 88.730 38.020 92.830 ;
        RECT 38.340 89.410 38.480 112.890 ;
        RECT 39.580 111.335 41.460 111.705 ;
        RECT 40.120 109.490 40.380 109.810 ;
        RECT 40.180 109.325 40.320 109.490 ;
        RECT 40.110 108.955 40.390 109.325 ;
        RECT 41.960 107.790 42.220 108.110 ;
        RECT 39.200 106.430 39.460 106.750 ;
        RECT 39.260 105.050 39.400 106.430 ;
        RECT 39.580 105.895 41.460 106.265 ;
        RECT 42.020 105.730 42.160 107.790 ;
        RECT 44.720 107.110 44.980 107.430 ;
        RECT 44.780 105.730 44.920 107.110 ;
        RECT 41.960 105.410 42.220 105.730 ;
        RECT 44.720 105.410 44.980 105.730 ;
        RECT 39.200 104.730 39.460 105.050 ;
        RECT 39.260 103.010 39.400 104.730 ;
        RECT 45.640 104.390 45.900 104.710 ;
        RECT 39.660 103.710 39.920 104.030 ;
        RECT 39.200 102.690 39.460 103.010 ;
        RECT 39.260 94.250 39.400 102.690 ;
        RECT 39.720 102.330 39.860 103.710 ;
        RECT 45.700 103.010 45.840 104.390 ;
        RECT 45.640 102.690 45.900 103.010 ;
        RECT 39.660 102.010 39.920 102.330 ;
        RECT 39.580 100.455 41.460 100.825 ;
        RECT 41.960 98.950 42.220 99.270 ;
        RECT 39.660 98.270 39.920 98.590 ;
        RECT 39.720 97.230 39.860 98.270 ;
        RECT 39.660 96.910 39.920 97.230 ;
        RECT 39.580 95.015 41.460 95.385 ;
        RECT 41.500 94.250 41.760 94.510 ;
        RECT 39.260 94.190 41.760 94.250 ;
        RECT 39.260 94.110 41.700 94.190 ;
        RECT 39.200 93.510 39.460 93.830 ;
        RECT 38.280 89.090 38.540 89.410 ;
        RECT 37.820 88.410 38.080 88.730 ;
        RECT 33.220 88.070 33.480 88.390 ;
        RECT 32.760 87.390 33.020 87.710 ;
        RECT 32.820 86.010 32.960 87.390 ;
        RECT 32.760 85.690 33.020 86.010 ;
        RECT 33.280 67.650 33.420 88.070 ;
        RECT 33.670 87.875 33.950 88.245 ;
        RECT 34.600 88.070 34.860 88.390 ;
        RECT 35.060 88.070 35.320 88.390 ;
        RECT 33.740 86.010 33.880 87.875 ;
        RECT 34.660 86.350 34.800 88.070 ;
        RECT 34.600 86.030 34.860 86.350 ;
        RECT 33.680 85.690 33.940 86.010 ;
        RECT 34.140 85.690 34.400 86.010 ;
        RECT 33.740 71.925 33.880 85.690 ;
        RECT 34.200 83.290 34.340 85.690 ;
        RECT 34.660 83.970 34.800 86.030 ;
        RECT 35.120 86.010 35.260 88.070 ;
        RECT 39.260 86.690 39.400 93.510 ;
        RECT 42.020 91.450 42.160 98.950 ;
        RECT 44.720 96.230 44.980 96.550 ;
        RECT 44.780 93.150 44.920 96.230 ;
        RECT 44.720 92.830 44.980 93.150 ;
        RECT 41.960 91.130 42.220 91.450 ;
        RECT 44.720 91.130 44.980 91.450 ;
        RECT 42.420 90.110 42.680 90.430 ;
        RECT 39.580 89.575 41.460 89.945 ;
        RECT 41.500 88.410 41.760 88.730 ;
        RECT 39.200 86.370 39.460 86.690 ;
        RECT 40.120 86.370 40.380 86.690 ;
        RECT 38.740 86.030 39.000 86.350 ;
        RECT 35.060 85.690 35.320 86.010 ;
        RECT 34.600 83.650 34.860 83.970 ;
        RECT 38.800 83.630 38.940 86.030 ;
        RECT 39.660 85.920 39.920 86.010 ;
        RECT 40.180 85.920 40.320 86.370 ;
        RECT 39.660 85.780 40.320 85.920 ;
        RECT 39.660 85.690 39.920 85.780 ;
        RECT 41.560 85.670 41.700 88.410 ;
        RECT 42.480 88.050 42.620 90.110 ;
        RECT 44.780 88.390 44.920 91.130 ;
        RECT 44.720 88.070 44.980 88.390 ;
        RECT 42.420 87.730 42.680 88.050 ;
        RECT 44.720 87.390 44.980 87.710 ;
        RECT 44.780 86.350 44.920 87.390 ;
        RECT 44.720 86.030 44.980 86.350 ;
        RECT 41.500 85.350 41.760 85.670 ;
        RECT 41.960 85.350 42.220 85.670 ;
        RECT 39.580 84.135 41.460 84.505 ;
        RECT 42.020 83.970 42.160 85.350 ;
        RECT 46.160 85.330 46.300 115.270 ;
        RECT 46.620 107.430 46.760 115.610 ;
        RECT 49.320 114.930 49.580 115.250 ;
        RECT 51.160 114.930 51.420 115.250 ;
        RECT 49.380 113.890 49.520 114.930 ;
        RECT 49.320 113.570 49.580 113.890 ;
        RECT 51.220 110.490 51.360 114.930 ;
        RECT 53.520 113.890 53.660 118.330 ;
        RECT 57.140 117.990 57.400 118.310 ;
        RECT 59.440 117.990 59.700 118.310 ;
        RECT 53.920 117.310 54.180 117.630 ;
        RECT 53.460 113.570 53.720 113.890 ;
        RECT 53.980 113.210 54.120 117.310 ;
        RECT 57.200 116.610 57.340 117.990 ;
        RECT 59.500 117.630 59.640 117.990 ;
        RECT 59.440 117.310 59.700 117.630 ;
        RECT 57.140 116.290 57.400 116.610 ;
        RECT 59.500 115.930 59.640 117.310 ;
        RECT 59.440 115.610 59.700 115.930 ;
        RECT 64.500 115.840 64.760 115.930 ;
        RECT 65.020 115.840 65.160 133.000 ;
        RECT 71.000 123.490 71.140 133.000 ;
        RECT 71.000 123.350 72.060 123.490 ;
        RECT 69.580 122.215 71.460 122.585 ;
        RECT 71.920 118.990 72.060 123.350 ;
        RECT 78.360 118.990 78.500 133.550 ;
        RECT 94.000 133.550 94.850 133.690 ;
        RECT 101.110 133.550 102.880 133.690 ;
        RECT 113.070 133.550 114.380 133.690 ;
        RECT 68.640 118.670 68.900 118.990 ;
        RECT 71.860 118.670 72.120 118.990 ;
        RECT 76.460 118.670 76.720 118.990 ;
        RECT 78.300 118.670 78.560 118.990 ;
        RECT 68.700 116.270 68.840 118.670 ;
        RECT 69.100 117.990 69.360 118.310 ;
        RECT 75.080 117.990 75.340 118.310 ;
        RECT 76.520 118.050 76.660 118.670 ;
        RECT 80.600 118.330 80.860 118.650 ;
        RECT 69.160 116.610 69.300 117.990 ;
        RECT 69.580 116.775 71.460 117.145 ;
        RECT 69.100 116.290 69.360 116.610 ;
        RECT 68.640 115.950 68.900 116.270 ;
        RECT 64.500 115.700 65.160 115.840 ;
        RECT 64.500 115.610 64.760 115.700 ;
        RECT 58.060 115.270 58.320 115.590 ;
        RECT 54.580 114.055 56.460 114.425 ;
        RECT 57.140 113.230 57.400 113.550 ;
        RECT 53.920 112.890 54.180 113.210 ;
        RECT 54.840 112.890 55.100 113.210 ;
        RECT 51.620 112.550 51.880 112.870 ;
        RECT 51.160 110.170 51.420 110.490 ;
        RECT 51.680 110.150 51.820 112.550 ;
        RECT 54.900 110.150 55.040 112.890 ;
        RECT 51.620 109.830 51.880 110.150 ;
        RECT 54.840 109.830 55.100 110.150 ;
        RECT 54.580 108.615 56.460 108.985 ;
        RECT 50.240 107.790 50.500 108.110 ;
        RECT 46.560 107.110 46.820 107.430 ;
        RECT 47.480 107.110 47.740 107.430 ;
        RECT 48.400 107.110 48.660 107.430 ;
        RECT 47.540 105.050 47.680 107.110 ;
        RECT 47.480 104.730 47.740 105.050 ;
        RECT 48.460 103.010 48.600 107.110 ;
        RECT 49.320 105.070 49.580 105.390 ;
        RECT 48.860 103.710 49.120 104.030 ;
        RECT 48.400 102.690 48.660 103.010 ;
        RECT 48.920 102.330 49.060 103.710 ;
        RECT 48.860 102.010 49.120 102.330 ;
        RECT 49.380 101.990 49.520 105.070 ;
        RECT 49.780 104.050 50.040 104.370 ;
        RECT 49.840 102.330 49.980 104.050 ;
        RECT 50.300 103.010 50.440 107.790 ;
        RECT 53.460 106.430 53.720 106.750 ;
        RECT 53.520 105.050 53.660 106.430 ;
        RECT 53.460 104.730 53.720 105.050 ;
        RECT 52.080 104.390 52.340 104.710 ;
        RECT 52.140 103.010 52.280 104.390 ;
        RECT 50.240 102.690 50.500 103.010 ;
        RECT 52.080 102.690 52.340 103.010 ;
        RECT 53.520 102.670 53.660 104.730 ;
        RECT 53.920 103.710 54.180 104.030 ;
        RECT 53.980 103.010 54.120 103.710 ;
        RECT 54.580 103.175 56.460 103.545 ;
        RECT 53.920 102.690 54.180 103.010 ;
        RECT 53.460 102.580 53.720 102.670 ;
        RECT 53.060 102.440 53.720 102.580 ;
        RECT 49.780 102.010 50.040 102.330 ;
        RECT 49.320 101.670 49.580 101.990 ;
        RECT 49.840 99.270 49.980 102.010 ;
        RECT 49.320 98.950 49.580 99.270 ;
        RECT 49.780 98.950 50.040 99.270 ;
        RECT 47.480 98.270 47.740 98.590 ;
        RECT 47.540 96.890 47.680 98.270 ;
        RECT 47.480 96.570 47.740 96.890 ;
        RECT 48.400 96.230 48.660 96.550 ;
        RECT 48.460 94.850 48.600 96.230 ;
        RECT 49.380 94.850 49.520 98.950 ;
        RECT 50.240 98.270 50.500 98.590 ;
        RECT 50.300 97.230 50.440 98.270 ;
        RECT 50.240 96.910 50.500 97.230 ;
        RECT 52.540 95.550 52.800 95.870 ;
        RECT 48.400 94.530 48.660 94.850 ;
        RECT 49.320 94.530 49.580 94.850 ;
        RECT 51.160 94.530 51.420 94.850 ;
        RECT 49.780 92.830 50.040 93.150 ;
        RECT 49.840 89.410 49.980 92.830 ;
        RECT 49.780 89.090 50.040 89.410 ;
        RECT 46.560 88.410 46.820 88.730 ;
        RECT 49.320 88.410 49.580 88.730 ;
        RECT 46.620 85.670 46.760 88.410 ;
        RECT 47.940 87.730 48.200 88.050 ;
        RECT 48.000 86.690 48.140 87.730 ;
        RECT 47.940 86.370 48.200 86.690 ;
        RECT 48.860 86.030 49.120 86.350 ;
        RECT 46.560 85.350 46.820 85.670 ;
        RECT 46.100 85.010 46.360 85.330 ;
        RECT 41.960 83.650 42.220 83.970 ;
        RECT 38.740 83.310 39.000 83.630 ;
        RECT 34.140 82.970 34.400 83.290 ;
        RECT 36.440 77.190 36.700 77.510 ;
        RECT 35.980 76.510 36.240 76.830 ;
        RECT 36.040 75.810 36.180 76.510 ;
        RECT 35.980 75.490 36.240 75.810 ;
        RECT 36.500 74.110 36.640 77.190 ;
        RECT 38.800 75.130 38.940 83.310 ;
        RECT 46.620 82.950 46.760 85.350 ;
        RECT 47.940 84.670 48.200 84.990 ;
        RECT 48.400 84.670 48.660 84.990 ;
        RECT 48.000 83.290 48.140 84.670 ;
        RECT 47.940 82.970 48.200 83.290 ;
        RECT 46.560 82.630 46.820 82.950 ;
        RECT 39.580 78.695 41.460 79.065 ;
        RECT 48.000 77.850 48.140 82.970 ;
        RECT 48.460 82.270 48.600 84.670 ;
        RECT 48.400 81.950 48.660 82.270 ;
        RECT 47.940 77.530 48.200 77.850 ;
        RECT 41.960 76.510 42.220 76.830 ;
        RECT 47.020 76.510 47.280 76.830 ;
        RECT 39.200 75.150 39.460 75.470 ;
        RECT 37.820 74.810 38.080 75.130 ;
        RECT 38.740 74.810 39.000 75.130 ;
        RECT 36.440 73.790 36.700 74.110 ;
        RECT 37.360 73.790 37.620 74.110 ;
        RECT 36.500 73.090 36.640 73.790 ;
        RECT 36.440 72.770 36.700 73.090 ;
        RECT 33.670 71.555 33.950 71.925 ;
        RECT 37.420 71.730 37.560 73.790 ;
        RECT 37.360 71.410 37.620 71.730 ;
        RECT 34.140 68.350 34.400 68.670 ;
        RECT 33.220 67.330 33.480 67.650 ;
        RECT 34.200 66.630 34.340 68.350 ;
        RECT 34.140 66.310 34.400 66.630 ;
        RECT 34.600 66.310 34.860 66.630 ;
        RECT 32.760 62.910 33.020 63.230 ;
        RECT 32.820 55.410 32.960 62.910 ;
        RECT 34.660 59.150 34.800 66.310 ;
        RECT 37.880 64.590 38.020 74.810 ;
        RECT 38.800 72.750 38.940 74.810 ;
        RECT 39.260 72.750 39.400 75.150 ;
        RECT 42.020 74.790 42.160 76.510 ;
        RECT 47.080 75.810 47.220 76.510 ;
        RECT 47.020 75.490 47.280 75.810 ;
        RECT 42.420 75.150 42.680 75.470 ;
        RECT 41.960 74.470 42.220 74.790 ;
        RECT 39.580 73.255 41.460 73.625 ;
        RECT 42.480 73.090 42.620 75.150 ;
        RECT 46.560 74.470 46.820 74.790 ;
        RECT 42.420 72.770 42.680 73.090 ;
        RECT 38.740 72.430 39.000 72.750 ;
        RECT 39.200 72.430 39.460 72.750 ;
        RECT 45.170 71.555 45.450 71.925 ;
        RECT 39.200 71.070 39.460 71.390 ;
        RECT 39.660 71.070 39.920 71.390 ;
        RECT 39.260 70.370 39.400 71.070 ;
        RECT 39.200 70.050 39.460 70.370 ;
        RECT 39.200 69.260 39.460 69.350 ;
        RECT 39.720 69.260 39.860 71.070 ;
        RECT 45.240 70.030 45.380 71.555 ;
        RECT 46.620 71.390 46.760 74.470 ;
        RECT 47.080 72.070 47.220 75.490 ;
        RECT 48.000 74.110 48.140 77.530 ;
        RECT 48.460 77.510 48.600 81.950 ;
        RECT 48.400 77.190 48.660 77.510 ;
        RECT 47.940 73.790 48.200 74.110 ;
        RECT 48.000 72.410 48.140 73.790 ;
        RECT 47.940 72.090 48.200 72.410 ;
        RECT 47.020 71.750 47.280 72.070 ;
        RECT 46.560 71.070 46.820 71.390 ;
        RECT 46.620 70.370 46.760 71.070 ;
        RECT 46.560 70.050 46.820 70.370 ;
        RECT 45.180 69.710 45.440 70.030 ;
        RECT 39.200 69.120 39.860 69.260 ;
        RECT 39.200 69.030 39.460 69.120 ;
        RECT 41.040 69.030 41.300 69.350 ;
        RECT 41.100 68.580 41.240 69.030 ;
        RECT 41.100 68.440 42.160 68.580 ;
        RECT 39.580 67.815 41.460 68.185 ;
        RECT 37.820 64.270 38.080 64.590 ;
        RECT 42.020 64.250 42.160 68.440 ;
        RECT 48.400 66.310 48.660 66.630 ;
        RECT 36.440 63.930 36.700 64.250 ;
        RECT 41.960 63.930 42.220 64.250 ;
        RECT 35.980 62.910 36.240 63.230 ;
        RECT 36.040 61.530 36.180 62.910 ;
        RECT 35.980 61.210 36.240 61.530 ;
        RECT 35.520 60.870 35.780 61.190 ;
        RECT 35.580 59.490 35.720 60.870 ;
        RECT 35.520 59.170 35.780 59.490 ;
        RECT 34.600 58.830 34.860 59.150 ;
        RECT 34.660 56.090 34.800 58.830 ;
        RECT 36.500 56.770 36.640 63.930 ;
        RECT 38.740 62.910 39.000 63.230 ;
        RECT 38.800 60.850 38.940 62.910 ;
        RECT 39.580 62.375 41.460 62.745 ;
        RECT 38.740 60.530 39.000 60.850 ;
        RECT 38.280 60.190 38.540 60.510 ;
        RECT 36.440 56.450 36.700 56.770 ;
        RECT 38.340 56.090 38.480 60.190 ;
        RECT 42.020 59.490 42.160 63.930 ;
        RECT 44.260 63.590 44.520 63.910 ;
        RECT 44.720 63.590 44.980 63.910 ;
        RECT 48.460 63.765 48.600 66.310 ;
        RECT 44.320 61.870 44.460 63.590 ;
        RECT 44.780 62.210 44.920 63.590 ;
        RECT 48.390 63.395 48.670 63.765 ;
        RECT 44.720 61.890 44.980 62.210 ;
        RECT 44.260 61.550 44.520 61.870 ;
        RECT 41.960 59.170 42.220 59.490 ;
        RECT 39.200 58.150 39.460 58.470 ;
        RECT 39.260 56.090 39.400 58.150 ;
        RECT 39.580 56.935 41.460 57.305 ;
        RECT 41.040 56.450 41.300 56.770 ;
        RECT 41.100 56.090 41.240 56.450 ;
        RECT 42.020 56.090 42.160 59.170 ;
        RECT 34.600 55.770 34.860 56.090 ;
        RECT 38.280 55.770 38.540 56.090 ;
        RECT 39.200 55.770 39.460 56.090 ;
        RECT 41.040 55.770 41.300 56.090 ;
        RECT 41.960 55.770 42.220 56.090 ;
        RECT 32.760 55.090 33.020 55.410 ;
        RECT 41.100 53.030 41.240 55.770 ;
        RECT 42.020 53.370 42.160 55.770 ;
        RECT 44.320 55.750 44.460 61.550 ;
        RECT 45.180 57.470 45.440 57.790 ;
        RECT 44.260 55.430 44.520 55.750 ;
        RECT 45.240 53.370 45.380 57.470 ;
        RECT 48.920 56.170 49.060 86.030 ;
        RECT 49.380 59.570 49.520 88.410 ;
        RECT 49.780 85.690 50.040 86.010 ;
        RECT 49.840 83.290 49.980 85.690 ;
        RECT 50.700 85.010 50.960 85.330 ;
        RECT 50.760 83.290 50.900 85.010 ;
        RECT 49.780 82.970 50.040 83.290 ;
        RECT 50.700 83.200 50.960 83.290 ;
        RECT 50.300 83.060 50.960 83.200 ;
        RECT 49.840 75.130 49.980 82.970 ;
        RECT 50.300 75.470 50.440 83.060 ;
        RECT 50.700 82.970 50.960 83.060 ;
        RECT 50.700 75.490 50.960 75.810 ;
        RECT 50.240 75.150 50.500 75.470 ;
        RECT 50.760 75.130 50.900 75.490 ;
        RECT 49.780 74.810 50.040 75.130 ;
        RECT 50.700 74.810 50.960 75.130 ;
        RECT 49.840 74.450 49.980 74.810 ;
        RECT 49.780 74.130 50.040 74.450 ;
        RECT 51.220 73.090 51.360 94.530 ;
        RECT 52.600 94.170 52.740 95.550 ;
        RECT 52.540 93.850 52.800 94.170 ;
        RECT 52.540 93.170 52.800 93.490 ;
        RECT 52.600 88.810 52.740 93.170 ;
        RECT 53.060 91.450 53.200 102.440 ;
        RECT 53.460 102.350 53.720 102.440 ;
        RECT 53.460 101.670 53.720 101.990 ;
        RECT 53.520 96.550 53.660 101.670 ;
        RECT 53.460 96.230 53.720 96.550 ;
        RECT 53.980 95.870 54.120 102.690 ;
        RECT 54.580 97.735 56.460 98.105 ;
        RECT 53.920 95.550 54.180 95.870 ;
        RECT 54.380 95.550 54.640 95.870 ;
        RECT 53.980 94.510 54.120 95.550 ;
        RECT 53.920 94.190 54.180 94.510 ;
        RECT 54.440 94.170 54.580 95.550 ;
        RECT 54.380 93.850 54.640 94.170 ;
        RECT 54.580 92.295 56.460 92.665 ;
        RECT 53.000 91.130 53.260 91.450 ;
        RECT 53.000 90.110 53.260 90.430 ;
        RECT 52.140 88.670 52.740 88.810 ;
        RECT 51.620 85.690 51.880 86.010 ;
        RECT 51.680 82.270 51.820 85.690 ;
        RECT 51.620 81.950 51.880 82.270 ;
        RECT 52.140 78.530 52.280 88.670 ;
        RECT 52.540 88.070 52.800 88.390 ;
        RECT 52.080 78.210 52.340 78.530 ;
        RECT 51.620 77.190 51.880 77.510 ;
        RECT 51.160 72.770 51.420 73.090 ;
        RECT 50.700 66.990 50.960 67.310 ;
        RECT 50.760 66.630 50.900 66.990 ;
        RECT 50.240 66.310 50.500 66.630 ;
        RECT 50.700 66.310 50.960 66.630 ;
        RECT 51.160 66.310 51.420 66.630 ;
        RECT 49.780 64.270 50.040 64.590 ;
        RECT 49.840 62.210 49.980 64.270 ;
        RECT 49.780 61.890 50.040 62.210 ;
        RECT 50.300 60.510 50.440 66.310 ;
        RECT 50.760 64.590 50.900 66.310 ;
        RECT 50.700 64.270 50.960 64.590 ;
        RECT 51.220 64.250 51.360 66.310 ;
        RECT 51.160 63.930 51.420 64.250 ;
        RECT 51.680 63.085 51.820 77.190 ;
        RECT 52.080 76.510 52.340 76.830 ;
        RECT 52.140 67.050 52.280 76.510 ;
        RECT 52.600 67.650 52.740 88.070 ;
        RECT 53.060 84.990 53.200 90.110 ;
        RECT 53.920 87.730 54.180 88.050 ;
        RECT 53.980 86.690 54.120 87.730 ;
        RECT 54.580 86.855 56.460 87.225 ;
        RECT 53.920 86.370 54.180 86.690 ;
        RECT 53.460 85.690 53.720 86.010 ;
        RECT 56.680 85.690 56.940 86.010 ;
        RECT 53.000 84.670 53.260 84.990 ;
        RECT 53.520 83.970 53.660 85.690 ;
        RECT 53.460 83.650 53.720 83.970 ;
        RECT 53.000 82.290 53.260 82.610 ;
        RECT 53.060 75.130 53.200 82.290 ;
        RECT 54.580 81.415 56.460 81.785 ;
        RECT 53.460 76.850 53.720 77.170 ;
        RECT 53.520 75.810 53.660 76.850 ;
        RECT 54.580 75.975 56.460 76.345 ;
        RECT 53.460 75.490 53.720 75.810 ;
        RECT 54.840 75.490 55.100 75.810 ;
        RECT 54.900 75.130 55.040 75.490 ;
        RECT 53.000 74.810 53.260 75.130 ;
        RECT 54.840 74.810 55.100 75.130 ;
        RECT 54.840 74.130 55.100 74.450 ;
        RECT 53.000 73.790 53.260 74.110 ;
        RECT 53.060 72.070 53.200 73.790 ;
        RECT 54.900 72.750 55.040 74.130 ;
        RECT 54.840 72.430 55.100 72.750 ;
        RECT 53.460 72.090 53.720 72.410 ;
        RECT 53.000 71.750 53.260 72.070 ;
        RECT 52.540 67.330 52.800 67.650 ;
        RECT 52.140 66.910 52.740 67.050 ;
        RECT 52.080 65.970 52.340 66.290 ;
        RECT 52.140 63.230 52.280 65.970 ;
        RECT 51.610 62.715 51.890 63.085 ;
        RECT 52.080 62.910 52.340 63.230 ;
        RECT 52.140 61.870 52.280 62.910 ;
        RECT 52.080 61.550 52.340 61.870 ;
        RECT 50.240 60.190 50.500 60.510 ;
        RECT 49.380 59.430 51.360 59.570 ;
        RECT 52.140 59.490 52.280 61.550 ;
        RECT 49.780 58.490 50.040 58.810 ;
        RECT 48.920 56.030 49.520 56.170 ;
        RECT 48.860 55.090 49.120 55.410 ;
        RECT 48.920 53.710 49.060 55.090 ;
        RECT 48.860 53.390 49.120 53.710 ;
        RECT 41.960 53.050 42.220 53.370 ;
        RECT 45.180 53.050 45.440 53.370 ;
        RECT 41.040 52.710 41.300 53.030 ;
        RECT 43.340 52.370 43.600 52.690 ;
        RECT 34.600 52.030 34.860 52.350 ;
        RECT 34.660 50.650 34.800 52.030 ;
        RECT 39.580 51.495 41.460 51.865 ;
        RECT 43.400 51.330 43.540 52.370 ;
        RECT 43.340 51.010 43.600 51.330 ;
        RECT 34.600 50.330 34.860 50.650 ;
        RECT 41.960 49.310 42.220 49.630 ;
        RECT 34.600 48.290 34.860 48.610 ;
        RECT 34.660 47.930 34.800 48.290 ;
        RECT 34.600 47.610 34.860 47.930 ;
        RECT 30.920 45.570 31.180 45.890 ;
        RECT 32.300 45.570 32.560 45.890 ;
        RECT 34.660 44.870 34.800 47.610 ;
        RECT 39.580 46.055 41.460 46.425 ;
        RECT 30.920 44.550 31.180 44.870 ;
        RECT 33.680 44.550 33.940 44.870 ;
        RECT 34.600 44.550 34.860 44.870 ;
        RECT 30.980 42.830 31.120 44.550 ;
        RECT 33.220 43.870 33.480 44.190 ;
        RECT 33.280 42.830 33.420 43.870 ;
        RECT 30.920 42.510 31.180 42.830 ;
        RECT 33.220 42.510 33.480 42.830 ;
        RECT 28.680 39.770 29.740 39.850 ;
        RECT 28.620 39.710 29.740 39.770 ;
        RECT 28.620 39.450 28.880 39.710 ;
        RECT 33.740 39.430 33.880 44.550 ;
        RECT 36.900 42.850 37.160 43.170 ;
        RECT 34.600 39.790 34.860 40.110 ;
        RECT 33.680 39.110 33.940 39.430 ;
        RECT 33.740 36.710 33.880 39.110 ;
        RECT 24.020 36.390 24.280 36.710 ;
        RECT 27.700 36.390 27.960 36.710 ;
        RECT 33.680 36.390 33.940 36.710 ;
        RECT 23.100 33.670 23.360 33.990 ;
        RECT 23.160 31.270 23.300 33.670 ;
        RECT 23.560 31.630 23.820 31.950 ;
        RECT 23.100 30.950 23.360 31.270 ;
        RECT 23.620 29.570 23.760 31.630 ;
        RECT 23.560 29.250 23.820 29.570 ;
        RECT 22.180 28.570 22.440 28.890 ;
        RECT 17.580 27.550 17.840 27.870 ;
        RECT 20.340 27.550 20.600 27.870 ;
        RECT 17.640 26.510 17.780 27.550 ;
        RECT 24.080 26.850 24.220 36.390 ;
        RECT 32.760 35.710 33.020 36.030 ;
        RECT 33.220 35.710 33.480 36.030 ;
        RECT 32.820 33.650 32.960 35.710 ;
        RECT 33.280 35.010 33.420 35.710 ;
        RECT 33.740 35.010 33.880 36.390 ;
        RECT 33.220 34.690 33.480 35.010 ;
        RECT 33.680 34.690 33.940 35.010 ;
        RECT 32.760 33.330 33.020 33.650 ;
        RECT 26.780 32.990 27.040 33.310 ;
        RECT 24.580 32.455 26.460 32.825 ;
        RECT 26.840 31.270 26.980 32.990 ;
        RECT 26.780 30.950 27.040 31.270 ;
        RECT 31.840 30.950 32.100 31.270 ;
        RECT 24.940 30.610 25.200 30.930 ;
        RECT 25.000 28.890 25.140 30.610 ;
        RECT 28.620 30.270 28.880 30.590 ;
        RECT 24.940 28.570 25.200 28.890 ;
        RECT 27.240 27.890 27.500 28.210 ;
        RECT 24.580 27.015 26.460 27.385 ;
        RECT 24.020 26.530 24.280 26.850 ;
        RECT 14.820 26.190 15.080 26.510 ;
        RECT 15.280 26.190 15.540 26.510 ;
        RECT 17.580 26.190 17.840 26.510 ;
        RECT 9.580 24.295 11.460 24.665 ;
        RECT 27.300 23.450 27.440 27.890 ;
        RECT 28.680 23.450 28.820 30.270 ;
        RECT 31.900 26.850 32.040 30.950 ;
        RECT 31.840 26.530 32.100 26.850 ;
        RECT 34.660 26.170 34.800 39.790 ;
        RECT 35.060 39.450 35.320 39.770 ;
        RECT 35.120 31.270 35.260 39.450 ;
        RECT 36.960 39.430 37.100 42.850 ;
        RECT 42.020 42.490 42.160 49.310 ;
        RECT 48.860 47.610 49.120 47.930 ;
        RECT 45.640 47.270 45.900 47.590 ;
        RECT 43.800 44.550 44.060 44.870 ;
        RECT 42.420 43.870 42.680 44.190 ;
        RECT 42.480 42.490 42.620 43.870 ;
        RECT 43.860 43.170 44.000 44.550 ;
        RECT 45.700 43.170 45.840 47.270 ;
        RECT 48.920 44.870 49.060 47.610 ;
        RECT 48.860 44.550 49.120 44.870 ;
        RECT 47.020 44.210 47.280 44.530 ;
        RECT 43.800 42.850 44.060 43.170 ;
        RECT 45.640 42.850 45.900 43.170 ;
        RECT 46.560 42.510 46.820 42.830 ;
        RECT 41.960 42.170 42.220 42.490 ;
        RECT 42.420 42.170 42.680 42.490 ;
        RECT 39.580 40.615 41.460 40.985 ;
        RECT 39.200 39.450 39.460 39.770 ;
        RECT 36.900 39.110 37.160 39.430 ;
        RECT 35.520 38.430 35.780 38.750 ;
        RECT 35.580 37.730 35.720 38.430 ;
        RECT 35.520 37.410 35.780 37.730 ;
        RECT 38.270 34.155 38.550 34.525 ;
        RECT 36.440 31.290 36.700 31.610 ;
        RECT 35.060 30.950 35.320 31.270 ;
        RECT 36.500 28.210 36.640 31.290 ;
        RECT 38.340 28.550 38.480 34.155 ;
        RECT 39.260 31.270 39.400 39.450 ;
        RECT 42.020 39.430 42.160 42.170 ;
        RECT 43.340 41.150 43.600 41.470 ;
        RECT 43.400 40.110 43.540 41.150 ;
        RECT 43.340 39.790 43.600 40.110 ;
        RECT 41.960 39.110 42.220 39.430 ;
        RECT 42.020 36.370 42.160 39.110 ;
        RECT 46.620 37.730 46.760 42.510 ;
        RECT 47.080 37.730 47.220 44.210 ;
        RECT 49.380 43.170 49.520 56.030 ;
        RECT 49.840 54.050 49.980 58.490 ;
        RECT 50.240 57.470 50.500 57.790 ;
        RECT 50.300 56.090 50.440 57.470 ;
        RECT 50.240 55.770 50.500 56.090 ;
        RECT 49.780 53.730 50.040 54.050 ;
        RECT 51.220 48.270 51.360 59.430 ;
        RECT 52.080 59.170 52.340 59.490 ;
        RECT 51.160 47.950 51.420 48.270 ;
        RECT 51.160 46.590 51.420 46.910 ;
        RECT 51.220 44.870 51.360 46.590 ;
        RECT 52.600 45.210 52.740 66.910 ;
        RECT 53.000 63.085 53.260 63.230 ;
        RECT 52.990 62.715 53.270 63.085 ;
        RECT 53.000 61.210 53.260 61.530 ;
        RECT 53.060 56.770 53.200 61.210 ;
        RECT 53.000 56.450 53.260 56.770 ;
        RECT 53.060 53.030 53.200 56.450 ;
        RECT 53.000 52.710 53.260 53.030 ;
        RECT 52.540 44.890 52.800 45.210 ;
        RECT 50.240 44.550 50.500 44.870 ;
        RECT 51.160 44.780 51.420 44.870 ;
        RECT 51.160 44.640 51.820 44.780 ;
        RECT 51.160 44.550 51.420 44.640 ;
        RECT 50.300 43.170 50.440 44.550 ;
        RECT 50.700 43.870 50.960 44.190 ;
        RECT 51.160 43.870 51.420 44.190 ;
        RECT 49.320 42.850 49.580 43.170 ;
        RECT 50.240 42.850 50.500 43.170 ;
        RECT 47.930 42.315 48.210 42.685 ;
        RECT 48.000 42.150 48.140 42.315 ;
        RECT 47.940 41.830 48.200 42.150 ;
        RECT 47.480 41.490 47.740 41.810 ;
        RECT 46.560 37.410 46.820 37.730 ;
        RECT 47.020 37.410 47.280 37.730 ;
        RECT 41.960 36.050 42.220 36.370 ;
        RECT 39.580 35.175 41.460 35.545 ;
        RECT 42.020 34.330 42.160 36.050 ;
        RECT 43.800 35.710 44.060 36.030 ;
        RECT 41.960 34.010 42.220 34.330 ;
        RECT 42.880 34.010 43.140 34.330 ;
        RECT 42.420 32.990 42.680 33.310 ;
        RECT 42.480 31.610 42.620 32.990 ;
        RECT 41.960 31.290 42.220 31.610 ;
        RECT 42.420 31.290 42.680 31.610 ;
        RECT 39.200 30.950 39.460 31.270 ;
        RECT 39.200 30.270 39.460 30.590 ;
        RECT 38.280 28.230 38.540 28.550 ;
        RECT 36.440 27.890 36.700 28.210 ;
        RECT 35.060 27.550 35.320 27.870 ;
        RECT 34.600 25.850 34.860 26.170 ;
        RECT 34.660 24.130 34.800 25.850 ;
        RECT 34.600 23.810 34.860 24.130 ;
        RECT 27.240 23.130 27.500 23.450 ;
        RECT 28.620 23.130 28.880 23.450 ;
        RECT 35.120 22.770 35.260 27.550 ;
        RECT 36.500 26.170 36.640 27.890 ;
        RECT 36.440 25.850 36.700 26.170 ;
        RECT 35.060 22.450 35.320 22.770 ;
        RECT 24.580 21.575 26.460 21.945 ;
        RECT 36.500 20.730 36.640 25.850 ;
        RECT 39.260 25.830 39.400 30.270 ;
        RECT 39.580 29.735 41.460 30.105 ;
        RECT 42.020 29.570 42.160 31.290 ;
        RECT 41.960 29.250 42.220 29.570 ;
        RECT 42.940 28.550 43.080 34.010 ;
        RECT 43.860 33.990 44.000 35.710 ;
        RECT 43.800 33.670 44.060 33.990 ;
        RECT 45.180 32.990 45.440 33.310 ;
        RECT 45.240 31.950 45.380 32.990 ;
        RECT 47.080 32.290 47.220 37.410 ;
        RECT 47.020 31.970 47.280 32.290 ;
        RECT 45.180 31.630 45.440 31.950 ;
        RECT 47.080 28.550 47.220 31.970 ;
        RECT 47.540 30.590 47.680 41.490 ;
        RECT 48.000 40.450 48.140 41.830 ;
        RECT 50.760 41.470 50.900 43.870 ;
        RECT 51.220 42.490 51.360 43.870 ;
        RECT 51.680 42.490 51.820 44.640 ;
        RECT 53.520 44.530 53.660 72.090 ;
        RECT 54.580 70.535 56.460 70.905 ;
        RECT 56.740 67.650 56.880 85.690 ;
        RECT 57.200 73.090 57.340 113.230 ;
        RECT 57.600 104.050 57.860 104.370 ;
        RECT 57.660 103.010 57.800 104.050 ;
        RECT 57.600 102.690 57.860 103.010 ;
        RECT 58.120 94.250 58.260 115.270 ;
        RECT 58.980 111.870 59.240 112.190 ;
        RECT 57.660 94.110 58.260 94.250 ;
        RECT 57.660 78.190 57.800 94.110 ;
        RECT 58.060 93.510 58.320 93.830 ;
        RECT 58.120 92.130 58.260 93.510 ;
        RECT 58.060 91.810 58.320 92.130 ;
        RECT 59.040 91.110 59.180 111.870 ;
        RECT 59.500 106.750 59.640 115.610 ;
        RECT 72.320 115.270 72.580 115.590 ;
        RECT 72.780 115.270 73.040 115.590 ;
        RECT 60.820 114.930 61.080 115.250 ;
        RECT 67.720 114.930 67.980 115.250 ;
        RECT 60.880 113.890 61.020 114.930 ;
        RECT 67.780 113.890 67.920 114.930 ;
        RECT 60.820 113.570 61.080 113.890 ;
        RECT 67.720 113.570 67.980 113.890 ;
        RECT 64.040 112.890 64.300 113.210 ;
        RECT 63.580 107.110 63.840 107.430 ;
        RECT 59.440 106.430 59.700 106.750 ;
        RECT 61.740 106.430 62.000 106.750 ;
        RECT 62.200 106.430 62.460 106.750 ;
        RECT 61.800 105.050 61.940 106.430 ;
        RECT 62.260 105.050 62.400 106.430 ;
        RECT 63.640 105.050 63.780 107.110 ;
        RECT 61.740 104.730 62.000 105.050 ;
        RECT 62.200 104.730 62.460 105.050 ;
        RECT 63.580 104.730 63.840 105.050 ;
        RECT 61.800 103.770 61.940 104.730 ;
        RECT 61.800 103.630 62.400 103.770 ;
        RECT 62.260 102.670 62.400 103.630 ;
        RECT 62.200 102.350 62.460 102.670 ;
        RECT 59.900 102.010 60.160 102.330 ;
        RECT 63.120 102.010 63.380 102.330 ;
        RECT 59.960 99.270 60.100 102.010 ;
        RECT 59.900 98.950 60.160 99.270 ;
        RECT 58.980 90.790 59.240 91.110 ;
        RECT 58.520 87.390 58.780 87.710 ;
        RECT 58.580 85.330 58.720 87.390 ;
        RECT 59.040 85.670 59.180 90.790 ;
        RECT 58.980 85.350 59.240 85.670 ;
        RECT 58.520 85.010 58.780 85.330 ;
        RECT 58.060 84.670 58.320 84.990 ;
        RECT 58.120 83.290 58.260 84.670 ;
        RECT 58.060 82.970 58.320 83.290 ;
        RECT 57.600 77.870 57.860 78.190 ;
        RECT 57.140 72.770 57.400 73.090 ;
        RECT 57.140 71.750 57.400 72.070 ;
        RECT 56.680 67.330 56.940 67.650 ;
        RECT 54.380 66.990 54.640 67.310 ;
        RECT 54.440 66.630 54.580 66.990 ;
        RECT 56.680 66.650 56.940 66.970 ;
        RECT 54.380 66.310 54.640 66.630 ;
        RECT 54.840 66.310 55.100 66.630 ;
        RECT 54.900 65.860 55.040 66.310 ;
        RECT 53.980 65.720 55.040 65.860 ;
        RECT 53.980 64.250 54.120 65.720 ;
        RECT 54.580 65.095 56.460 65.465 ;
        RECT 56.740 64.590 56.880 66.650 ;
        RECT 57.200 64.930 57.340 71.750 ;
        RECT 58.060 71.410 58.320 71.730 ;
        RECT 58.120 70.370 58.260 71.410 ;
        RECT 58.060 70.050 58.320 70.370 ;
        RECT 59.040 69.350 59.180 85.350 ;
        RECT 59.440 75.490 59.700 75.810 ;
        RECT 59.500 74.110 59.640 75.490 ;
        RECT 59.440 73.790 59.700 74.110 ;
        RECT 59.440 69.710 59.700 70.030 ;
        RECT 58.980 69.260 59.240 69.350 ;
        RECT 58.120 69.120 59.240 69.260 ;
        RECT 57.590 65.435 57.870 65.805 ;
        RECT 57.140 64.610 57.400 64.930 ;
        RECT 56.680 64.270 56.940 64.590 ;
        RECT 53.920 63.930 54.180 64.250 ;
        RECT 56.680 63.590 56.940 63.910 ;
        RECT 54.580 59.655 56.460 60.025 ;
        RECT 53.920 58.830 54.180 59.150 ;
        RECT 53.980 54.050 54.120 58.830 ;
        RECT 54.380 58.150 54.640 58.470 ;
        RECT 54.440 56.430 54.580 58.150 ;
        RECT 54.380 56.110 54.640 56.430 ;
        RECT 54.580 54.215 56.460 54.585 ;
        RECT 56.740 54.050 56.880 63.590 ;
        RECT 57.660 59.150 57.800 65.435 ;
        RECT 57.600 58.830 57.860 59.150 ;
        RECT 58.120 56.090 58.260 69.120 ;
        RECT 58.980 69.030 59.240 69.120 ;
        RECT 59.500 68.670 59.640 69.710 ;
        RECT 59.440 68.350 59.700 68.670 ;
        RECT 58.510 66.795 58.790 67.165 ;
        RECT 58.580 66.630 58.720 66.795 ;
        RECT 58.520 66.310 58.780 66.630 ;
        RECT 58.980 65.970 59.240 66.290 ;
        RECT 59.040 64.930 59.180 65.970 ;
        RECT 58.980 64.610 59.240 64.930 ;
        RECT 59.040 64.250 59.180 64.610 ;
        RECT 58.980 63.930 59.240 64.250 ;
        RECT 59.040 62.210 59.180 63.930 ;
        RECT 58.980 61.890 59.240 62.210 ;
        RECT 59.500 61.100 59.640 68.350 ;
        RECT 59.960 65.805 60.100 98.950 ;
        RECT 63.180 97.570 63.320 102.010 ;
        RECT 63.120 97.250 63.380 97.570 ;
        RECT 61.280 96.570 61.540 96.890 ;
        RECT 62.660 96.570 62.920 96.890 ;
        RECT 63.120 96.800 63.380 96.890 ;
        RECT 63.640 96.800 63.780 104.730 ;
        RECT 63.120 96.660 63.780 96.800 ;
        RECT 63.120 96.570 63.380 96.660 ;
        RECT 60.820 95.550 61.080 95.870 ;
        RECT 60.880 93.830 61.020 95.550 ;
        RECT 60.820 93.510 61.080 93.830 ;
        RECT 61.340 92.130 61.480 96.570 ;
        RECT 62.720 92.130 62.860 96.570 ;
        RECT 61.280 91.810 61.540 92.130 ;
        RECT 62.660 91.810 62.920 92.130 ;
        RECT 63.180 91.530 63.320 96.570 ;
        RECT 60.360 91.130 60.620 91.450 ;
        RECT 62.260 91.390 63.320 91.530 ;
        RECT 59.890 65.435 60.170 65.805 ;
        RECT 59.900 63.930 60.160 64.250 ;
        RECT 58.580 60.960 59.640 61.100 ;
        RECT 58.060 55.770 58.320 56.090 ;
        RECT 53.920 53.730 54.180 54.050 ;
        RECT 56.680 53.730 56.940 54.050 ;
        RECT 54.580 48.775 56.460 49.145 ;
        RECT 54.840 47.610 55.100 47.930 ;
        RECT 54.900 45.405 55.040 47.610 ;
        RECT 56.680 46.930 56.940 47.250 ;
        RECT 55.300 46.590 55.560 46.910 ;
        RECT 53.920 44.890 54.180 45.210 ;
        RECT 54.830 45.035 55.110 45.405 ;
        RECT 53.460 44.210 53.720 44.530 ;
        RECT 51.160 42.170 51.420 42.490 ;
        RECT 51.620 42.170 51.880 42.490 ;
        RECT 53.460 41.830 53.720 42.150 ;
        RECT 50.700 41.150 50.960 41.470 ;
        RECT 53.520 40.450 53.660 41.830 ;
        RECT 53.980 41.810 54.120 44.890 ;
        RECT 54.900 44.870 55.040 45.035 ;
        RECT 55.360 44.870 55.500 46.590 ;
        RECT 56.740 44.870 56.880 46.930 ;
        RECT 58.060 45.570 58.320 45.890 ;
        RECT 58.120 44.870 58.260 45.570 ;
        RECT 54.840 44.550 55.100 44.870 ;
        RECT 55.300 44.550 55.560 44.870 ;
        RECT 56.680 44.550 56.940 44.870 ;
        RECT 58.060 44.550 58.320 44.870 ;
        RECT 54.580 43.335 56.460 43.705 ;
        RECT 54.380 42.850 54.640 43.170 ;
        RECT 54.440 42.685 54.580 42.850 ;
        RECT 54.370 42.315 54.650 42.685 ;
        RECT 56.740 42.490 56.880 44.550 ;
        RECT 56.680 42.170 56.940 42.490 ;
        RECT 57.140 41.830 57.400 42.150 ;
        RECT 53.920 41.490 54.180 41.810 ;
        RECT 57.200 40.530 57.340 41.830 ;
        RECT 47.940 40.130 48.200 40.450 ;
        RECT 53.460 40.130 53.720 40.450 ;
        RECT 56.280 40.390 57.340 40.530 ;
        RECT 58.120 40.450 58.260 44.550 ;
        RECT 48.000 36.710 48.140 40.130 ;
        RECT 56.280 39.430 56.420 40.390 ;
        RECT 56.220 39.110 56.480 39.430 ;
        RECT 54.580 37.895 56.460 38.265 ;
        RECT 47.940 36.390 48.200 36.710 ;
        RECT 47.480 30.270 47.740 30.590 ;
        RECT 42.880 28.230 43.140 28.550 ;
        RECT 47.020 28.230 47.280 28.550 ;
        RECT 46.100 27.890 46.360 28.210 ;
        RECT 42.880 27.550 43.140 27.870 ;
        RECT 42.940 26.510 43.080 27.550 ;
        RECT 42.880 26.190 43.140 26.510 ;
        RECT 39.200 25.510 39.460 25.830 ;
        RECT 39.580 24.295 41.460 24.665 ;
        RECT 46.160 23.110 46.300 27.890 ;
        RECT 47.540 27.870 47.680 30.270 ;
        RECT 48.000 28.890 48.140 36.390 ;
        RECT 56.740 36.370 56.880 40.390 ;
        RECT 58.060 40.130 58.320 40.450 ;
        RECT 57.140 39.790 57.400 40.110 ;
        RECT 57.200 39.430 57.340 39.790 ;
        RECT 57.140 39.110 57.400 39.430 ;
        RECT 57.200 37.390 57.340 39.110 ;
        RECT 58.580 37.730 58.720 60.960 ;
        RECT 59.960 58.810 60.100 63.930 ;
        RECT 59.900 58.490 60.160 58.810 ;
        RECT 59.960 56.770 60.100 58.490 ;
        RECT 59.900 56.450 60.160 56.770 ;
        RECT 58.980 55.770 59.240 56.090 ;
        RECT 59.040 44.870 59.180 55.770 ;
        RECT 60.420 50.730 60.560 91.130 ;
        RECT 60.820 82.290 61.080 82.610 ;
        RECT 60.880 81.250 61.020 82.290 ;
        RECT 60.820 80.930 61.080 81.250 ;
        RECT 62.260 80.570 62.400 91.390 ;
        RECT 63.580 90.790 63.840 91.110 ;
        RECT 63.640 86.010 63.780 90.790 ;
        RECT 63.580 85.690 63.840 86.010 ;
        RECT 62.660 82.970 62.920 83.290 ;
        RECT 62.200 80.250 62.460 80.570 ;
        RECT 62.260 78.190 62.400 80.250 ;
        RECT 62.200 77.870 62.460 78.190 ;
        RECT 60.820 74.810 61.080 75.130 ;
        RECT 60.880 70.030 61.020 74.810 ;
        RECT 62.200 74.470 62.460 74.790 ;
        RECT 62.260 72.070 62.400 74.470 ;
        RECT 62.200 71.750 62.460 72.070 ;
        RECT 60.820 69.710 61.080 70.030 ;
        RECT 62.260 69.770 62.400 71.750 ;
        RECT 62.720 70.370 62.860 82.970 ;
        RECT 63.120 80.250 63.380 80.570 ;
        RECT 63.180 78.530 63.320 80.250 ;
        RECT 63.120 78.210 63.380 78.530 ;
        RECT 63.640 77.850 63.780 85.690 ;
        RECT 64.100 79.890 64.240 112.890 ;
        RECT 69.580 111.335 71.460 111.705 ;
        RECT 72.380 110.470 72.520 115.270 ;
        RECT 72.840 113.210 72.980 115.270 ;
        RECT 75.140 113.890 75.280 117.990 ;
        RECT 76.060 117.910 76.660 118.050 ;
        RECT 76.060 116.610 76.200 117.910 ;
        RECT 76.460 117.310 76.720 117.630 ;
        RECT 76.000 116.290 76.260 116.610 ;
        RECT 76.000 115.840 76.260 115.930 ;
        RECT 76.520 115.840 76.660 117.310 ;
        RECT 80.660 115.930 80.800 118.330 ;
        RECT 82.960 118.050 83.100 133.000 ;
        RECT 84.580 119.495 86.460 119.865 ;
        RECT 88.940 119.330 89.080 133.000 ;
        RECT 88.880 119.010 89.140 119.330 ;
        RECT 94.000 118.990 94.140 133.550 ;
        RECT 99.580 122.215 101.460 122.585 ;
        RECT 96.240 120.710 96.500 121.030 ;
        RECT 89.800 118.670 90.060 118.990 ;
        RECT 93.940 118.670 94.200 118.990 ;
        RECT 82.440 117.650 82.700 117.970 ;
        RECT 82.960 117.910 83.560 118.050 ;
        RECT 84.740 117.990 85.000 118.310 ;
        RECT 76.000 115.700 76.660 115.840 ;
        RECT 76.000 115.610 76.260 115.700 ;
        RECT 75.080 113.570 75.340 113.890 ;
        RECT 72.780 112.890 73.040 113.210 ;
        RECT 73.240 112.890 73.500 113.210 ;
        RECT 76.000 112.890 76.260 113.210 ;
        RECT 72.380 110.330 72.980 110.470 ;
        RECT 64.960 107.450 65.220 107.770 ;
        RECT 65.020 100.290 65.160 107.450 ;
        RECT 66.340 106.430 66.600 106.750 ;
        RECT 66.400 104.370 66.540 106.430 ;
        RECT 69.580 105.895 71.460 106.265 ;
        RECT 66.340 104.050 66.600 104.370 ;
        RECT 68.640 103.710 68.900 104.030 ;
        RECT 70.940 103.710 71.200 104.030 ;
        RECT 64.960 99.970 65.220 100.290 ;
        RECT 68.180 99.290 68.440 99.610 ;
        RECT 64.500 96.570 64.760 96.890 ;
        RECT 64.560 93.490 64.700 96.570 ;
        RECT 64.960 93.510 65.220 93.830 ;
        RECT 64.500 93.170 64.760 93.490 ;
        RECT 65.020 91.790 65.160 93.510 ;
        RECT 66.800 92.830 67.060 93.150 ;
        RECT 66.860 92.130 67.000 92.830 ;
        RECT 66.800 91.810 67.060 92.130 ;
        RECT 64.960 91.470 65.220 91.790 ;
        RECT 66.340 86.030 66.600 86.350 ;
        RECT 66.400 83.970 66.540 86.030 ;
        RECT 66.340 83.650 66.600 83.970 ;
        RECT 65.420 83.310 65.680 83.630 ;
        RECT 64.960 82.630 65.220 82.950 ;
        RECT 64.500 80.930 64.760 81.250 ;
        RECT 64.560 80.230 64.700 80.930 ;
        RECT 64.500 79.910 64.760 80.230 ;
        RECT 64.040 79.570 64.300 79.890 ;
        RECT 64.040 77.870 64.300 78.190 ;
        RECT 63.580 77.530 63.840 77.850 ;
        RECT 63.580 71.750 63.840 72.070 ;
        RECT 62.660 70.050 62.920 70.370 ;
        RECT 61.340 69.690 62.400 69.770 ;
        RECT 61.280 69.630 62.460 69.690 ;
        RECT 61.280 69.370 61.540 69.630 ;
        RECT 62.200 69.370 62.460 69.630 ;
        RECT 62.720 68.670 62.860 70.050 ;
        RECT 63.640 69.350 63.780 71.750 ;
        RECT 63.580 69.030 63.840 69.350 ;
        RECT 63.120 68.690 63.380 69.010 ;
        RECT 62.660 68.350 62.920 68.670 ;
        RECT 63.180 67.650 63.320 68.690 ;
        RECT 63.120 67.330 63.380 67.650 ;
        RECT 62.660 63.930 62.920 64.250 ;
        RECT 61.270 63.395 61.550 63.765 ;
        RECT 61.340 63.230 61.480 63.395 ;
        RECT 62.200 63.250 62.460 63.570 ;
        RECT 61.280 62.910 61.540 63.230 ;
        RECT 62.260 61.870 62.400 63.250 ;
        RECT 62.200 61.550 62.460 61.870 ;
        RECT 61.740 60.870 62.000 61.190 ;
        RECT 59.500 50.590 60.560 50.730 ;
        RECT 61.800 55.490 61.940 60.870 ;
        RECT 62.200 55.490 62.460 55.750 ;
        RECT 61.800 55.430 62.460 55.490 ;
        RECT 61.800 55.350 62.400 55.430 ;
        RECT 58.980 44.550 59.240 44.870 ;
        RECT 58.980 42.170 59.240 42.490 ;
        RECT 59.040 38.750 59.180 42.170 ;
        RECT 59.500 39.770 59.640 50.590 ;
        RECT 60.360 47.610 60.620 47.930 ;
        RECT 60.420 44.870 60.560 47.610 ;
        RECT 61.270 45.035 61.550 45.405 ;
        RECT 60.360 44.725 60.620 44.870 ;
        RECT 60.350 44.355 60.630 44.725 ;
        RECT 61.340 44.190 61.480 45.035 ;
        RECT 59.900 43.870 60.160 44.190 ;
        RECT 61.280 43.870 61.540 44.190 ;
        RECT 59.960 42.830 60.100 43.870 ;
        RECT 59.900 42.510 60.160 42.830 ;
        RECT 61.800 42.490 61.940 55.350 ;
        RECT 62.720 55.070 62.860 63.930 ;
        RECT 63.180 62.210 63.320 67.330 ;
        RECT 63.640 64.250 63.780 69.030 ;
        RECT 63.580 63.930 63.840 64.250 ;
        RECT 63.120 61.890 63.380 62.210 ;
        RECT 64.100 56.770 64.240 77.870 ;
        RECT 64.560 69.690 64.700 79.910 ;
        RECT 65.020 69.885 65.160 82.630 ;
        RECT 64.500 69.370 64.760 69.690 ;
        RECT 64.950 69.515 65.230 69.885 ;
        RECT 65.020 63.765 65.160 69.515 ;
        RECT 64.950 63.395 65.230 63.765 ;
        RECT 64.500 58.490 64.760 58.810 ;
        RECT 64.040 56.450 64.300 56.770 ;
        RECT 62.660 54.750 62.920 55.070 ;
        RECT 62.720 53.370 62.860 54.750 ;
        RECT 62.660 53.050 62.920 53.370 ;
        RECT 62.200 52.030 62.460 52.350 ;
        RECT 62.260 48.610 62.400 52.030 ;
        RECT 62.200 48.290 62.460 48.610 ;
        RECT 62.720 44.725 62.860 53.050 ;
        RECT 64.100 50.310 64.240 56.450 ;
        RECT 64.560 55.750 64.700 58.490 ;
        RECT 64.500 55.430 64.760 55.750 ;
        RECT 65.480 52.350 65.620 83.310 ;
        RECT 66.860 82.950 67.000 91.810 ;
        RECT 67.260 91.470 67.520 91.790 ;
        RECT 67.320 88.390 67.460 91.470 ;
        RECT 68.240 91.110 68.380 99.290 ;
        RECT 68.700 99.270 68.840 103.710 ;
        RECT 71.000 102.670 71.140 103.710 ;
        RECT 70.940 102.350 71.200 102.670 ;
        RECT 72.320 100.990 72.580 101.310 ;
        RECT 69.580 100.455 71.460 100.825 ;
        RECT 68.640 98.950 68.900 99.270 ;
        RECT 69.100 98.950 69.360 99.270 ;
        RECT 68.700 91.790 68.840 98.950 ;
        RECT 69.160 94.170 69.300 98.950 ;
        RECT 72.380 98.590 72.520 100.990 ;
        RECT 72.840 99.690 72.980 110.330 ;
        RECT 73.300 104.710 73.440 112.890 ;
        RECT 73.240 104.390 73.500 104.710 ;
        RECT 75.080 104.390 75.340 104.710 ;
        RECT 75.140 102.330 75.280 104.390 ;
        RECT 75.080 102.010 75.340 102.330 ;
        RECT 75.540 100.990 75.800 101.310 ;
        RECT 72.840 99.550 73.440 99.690 ;
        RECT 72.780 98.950 73.040 99.270 ;
        RECT 72.320 98.270 72.580 98.590 ;
        RECT 72.380 96.890 72.520 98.270 ;
        RECT 72.840 97.570 72.980 98.950 ;
        RECT 72.780 97.250 73.040 97.570 ;
        RECT 72.320 96.570 72.580 96.890 ;
        RECT 69.580 95.015 71.460 95.385 ;
        RECT 69.100 93.850 69.360 94.170 ;
        RECT 69.160 93.490 69.300 93.850 ;
        RECT 69.100 93.170 69.360 93.490 ;
        RECT 68.640 91.470 68.900 91.790 ;
        RECT 68.180 90.790 68.440 91.110 ;
        RECT 69.160 88.390 69.300 93.170 ;
        RECT 69.580 89.575 71.460 89.945 ;
        RECT 67.260 88.070 67.520 88.390 ;
        RECT 67.720 88.070 67.980 88.390 ;
        RECT 68.180 88.070 68.440 88.390 ;
        RECT 69.100 88.070 69.360 88.390 ;
        RECT 67.780 86.350 67.920 88.070 ;
        RECT 67.720 86.030 67.980 86.350 ;
        RECT 67.260 85.350 67.520 85.670 ;
        RECT 68.240 85.410 68.380 88.070 ;
        RECT 68.640 87.730 68.900 88.050 ;
        RECT 68.700 86.010 68.840 87.730 ;
        RECT 68.640 85.690 68.900 86.010 ;
        RECT 66.800 82.630 67.060 82.950 ;
        RECT 67.320 82.270 67.460 85.350 ;
        RECT 67.780 85.270 68.380 85.410 ;
        RECT 67.780 84.990 67.920 85.270 ;
        RECT 67.720 84.670 67.980 84.990 ;
        RECT 67.780 82.950 67.920 84.670 ;
        RECT 68.700 83.630 68.840 85.690 ;
        RECT 68.640 83.310 68.900 83.630 ;
        RECT 67.720 82.630 67.980 82.950 ;
        RECT 67.260 81.950 67.520 82.270 ;
        RECT 67.320 77.510 67.460 81.950 ;
        RECT 67.260 77.190 67.520 77.510 ;
        RECT 67.260 74.810 67.520 75.130 ;
        RECT 67.320 72.410 67.460 74.810 ;
        RECT 67.780 73.090 67.920 82.630 ;
        RECT 69.160 81.250 69.300 88.070 ;
        RECT 71.860 86.370 72.120 86.690 ;
        RECT 69.580 84.135 71.460 84.505 ;
        RECT 71.920 82.270 72.060 86.370 ;
        RECT 72.380 86.350 72.520 96.570 ;
        RECT 73.300 88.810 73.440 99.550 ;
        RECT 75.600 98.930 75.740 100.990 ;
        RECT 75.540 98.610 75.800 98.930 ;
        RECT 75.080 96.570 75.340 96.890 ;
        RECT 75.140 94.850 75.280 96.570 ;
        RECT 75.080 94.530 75.340 94.850 ;
        RECT 72.840 88.670 73.440 88.810 ;
        RECT 72.320 86.030 72.580 86.350 ;
        RECT 72.320 84.670 72.580 84.990 ;
        RECT 72.380 82.950 72.520 84.670 ;
        RECT 72.320 82.630 72.580 82.950 ;
        RECT 71.860 81.950 72.120 82.270 ;
        RECT 69.100 80.930 69.360 81.250 ;
        RECT 69.160 78.190 69.300 80.930 ;
        RECT 69.580 78.695 71.460 79.065 ;
        RECT 69.100 77.870 69.360 78.190 ;
        RECT 68.180 77.530 68.440 77.850 ;
        RECT 68.240 74.790 68.380 77.530 ;
        RECT 69.100 75.490 69.360 75.810 ;
        RECT 68.180 74.470 68.440 74.790 ;
        RECT 67.720 72.770 67.980 73.090 ;
        RECT 68.240 72.750 68.380 74.470 ;
        RECT 68.180 72.430 68.440 72.750 ;
        RECT 67.260 72.090 67.520 72.410 ;
        RECT 69.160 72.070 69.300 75.490 ;
        RECT 69.580 73.255 71.460 73.625 ;
        RECT 72.840 72.750 72.980 88.670 ;
        RECT 73.240 88.070 73.500 88.390 ;
        RECT 73.300 86.690 73.440 88.070 ;
        RECT 73.240 86.370 73.500 86.690 ;
        RECT 74.160 80.590 74.420 80.910 ;
        RECT 73.700 79.230 73.960 79.550 ;
        RECT 73.760 77.170 73.900 79.230 ;
        RECT 74.220 78.530 74.360 80.590 ;
        RECT 74.160 78.210 74.420 78.530 ;
        RECT 73.700 76.850 73.960 77.170 ;
        RECT 73.760 75.810 73.900 76.850 ;
        RECT 73.700 75.490 73.960 75.810 ;
        RECT 74.160 75.150 74.420 75.470 ;
        RECT 72.780 72.430 73.040 72.750 ;
        RECT 74.220 72.070 74.360 75.150 ;
        RECT 76.060 74.450 76.200 112.890 ;
        RECT 76.520 105.050 76.660 115.700 ;
        RECT 80.600 115.610 80.860 115.930 ;
        RECT 77.380 114.930 77.640 115.250 ;
        RECT 77.440 113.890 77.580 114.930 ;
        RECT 77.380 113.570 77.640 113.890 ;
        RECT 81.060 112.890 81.320 113.210 ;
        RECT 78.300 106.430 78.560 106.750 ;
        RECT 76.460 104.730 76.720 105.050 ;
        RECT 78.360 104.710 78.500 106.430 ;
        RECT 78.300 104.390 78.560 104.710 ;
        RECT 77.380 98.270 77.640 98.590 ;
        RECT 77.440 96.210 77.580 98.270 ;
        RECT 78.300 96.230 78.560 96.550 ;
        RECT 77.380 95.890 77.640 96.210 ;
        RECT 77.440 93.150 77.580 95.890 ;
        RECT 78.360 94.170 78.500 96.230 ;
        RECT 78.300 93.850 78.560 94.170 ;
        RECT 76.460 92.830 76.720 93.150 ;
        RECT 77.380 92.830 77.640 93.150 ;
        RECT 76.520 87.710 76.660 92.830 ;
        RECT 77.440 89.070 77.580 92.830 ;
        RECT 77.380 88.750 77.640 89.070 ;
        RECT 76.920 87.730 77.180 88.050 ;
        RECT 76.460 87.390 76.720 87.710 ;
        RECT 76.520 86.690 76.660 87.390 ;
        RECT 76.460 86.370 76.720 86.690 ;
        RECT 76.980 82.950 77.120 87.730 ;
        RECT 77.380 86.030 77.640 86.350 ;
        RECT 76.920 82.630 77.180 82.950 ;
        RECT 77.440 82.010 77.580 86.030 ;
        RECT 78.360 85.670 78.500 93.850 ;
        RECT 80.600 88.070 80.860 88.390 ;
        RECT 80.660 86.350 80.800 88.070 ;
        RECT 81.120 86.690 81.260 112.890 ;
        RECT 82.500 110.490 82.640 117.650 ;
        RECT 82.900 117.310 83.160 117.630 ;
        RECT 82.960 115.590 83.100 117.310 ;
        RECT 83.420 115.930 83.560 117.910 ;
        RECT 84.800 116.610 84.940 117.990 ;
        RECT 89.860 116.610 90.000 118.670 ;
        RECT 96.300 117.630 96.440 120.710 ;
        RECT 99.000 120.370 99.260 120.690 ;
        RECT 96.700 117.990 96.960 118.310 ;
        RECT 97.620 117.990 97.880 118.310 ;
        RECT 96.240 117.310 96.500 117.630 ;
        RECT 84.740 116.290 85.000 116.610 ;
        RECT 89.800 116.290 90.060 116.610 ;
        RECT 83.360 115.610 83.620 115.930 ;
        RECT 96.300 115.590 96.440 117.310 ;
        RECT 96.760 116.610 96.900 117.990 ;
        RECT 96.700 116.290 96.960 116.610 ;
        RECT 97.680 115.930 97.820 117.990 ;
        RECT 97.620 115.610 97.880 115.930 ;
        RECT 82.900 115.270 83.160 115.590 ;
        RECT 87.040 115.270 87.300 115.590 ;
        RECT 91.640 115.270 91.900 115.590 ;
        RECT 94.400 115.270 94.660 115.590 ;
        RECT 96.240 115.270 96.500 115.590 ;
        RECT 84.580 114.055 86.460 114.425 ;
        RECT 82.440 110.170 82.700 110.490 ;
        RECT 87.100 110.470 87.240 115.270 ;
        RECT 87.100 110.330 89.080 110.470 ;
        RECT 83.820 109.490 84.080 109.810 ;
        RECT 83.360 107.450 83.620 107.770 ;
        RECT 82.900 107.110 83.160 107.430 ;
        RECT 81.980 104.050 82.240 104.370 ;
        RECT 82.040 103.010 82.180 104.050 ;
        RECT 81.980 102.690 82.240 103.010 ;
        RECT 82.960 102.330 83.100 107.110 ;
        RECT 83.420 103.010 83.560 107.450 ;
        RECT 83.360 102.690 83.620 103.010 ;
        RECT 82.900 102.010 83.160 102.330 ;
        RECT 83.360 92.830 83.620 93.150 ;
        RECT 82.440 89.090 82.700 89.410 ;
        RECT 82.500 88.390 82.640 89.090 ;
        RECT 82.440 88.130 82.700 88.390 ;
        RECT 82.040 88.070 82.700 88.130 ;
        RECT 82.900 88.070 83.160 88.390 ;
        RECT 82.040 87.990 82.640 88.070 ;
        RECT 81.060 86.370 81.320 86.690 ;
        RECT 80.600 86.030 80.860 86.350 ;
        RECT 78.300 85.350 78.560 85.670 ;
        RECT 77.840 82.970 78.100 83.290 ;
        RECT 76.980 81.870 77.580 82.010 ;
        RECT 76.980 80.570 77.120 81.870 ;
        RECT 76.920 80.250 77.180 80.570 ;
        RECT 76.460 75.040 76.720 75.130 ;
        RECT 76.980 75.040 77.120 80.250 ;
        RECT 77.900 77.170 78.040 82.970 ;
        RECT 78.360 77.850 78.500 85.350 ;
        RECT 82.040 84.990 82.180 87.990 ;
        RECT 82.440 87.390 82.700 87.710 ;
        RECT 82.500 86.350 82.640 87.390 ;
        RECT 82.440 86.030 82.700 86.350 ;
        RECT 82.440 85.350 82.700 85.670 ;
        RECT 79.680 84.670 79.940 84.990 ;
        RECT 81.980 84.670 82.240 84.990 ;
        RECT 79.220 83.650 79.480 83.970 ;
        RECT 79.280 80.570 79.420 83.650 ;
        RECT 79.220 80.250 79.480 80.570 ;
        RECT 79.280 79.970 79.420 80.250 ;
        RECT 79.740 80.230 79.880 84.670 ;
        RECT 78.820 79.830 79.420 79.970 ;
        RECT 79.680 79.910 79.940 80.230 ;
        RECT 78.300 77.530 78.560 77.850 ;
        RECT 77.840 76.850 78.100 77.170 ;
        RECT 76.460 74.900 77.120 75.040 ;
        RECT 78.300 75.040 78.560 75.130 ;
        RECT 78.820 75.040 78.960 79.830 ;
        RECT 79.220 76.510 79.480 76.830 ;
        RECT 78.300 74.900 78.960 75.040 ;
        RECT 76.460 74.810 76.720 74.900 ;
        RECT 78.300 74.810 78.560 74.900 ;
        RECT 76.000 74.130 76.260 74.450 ;
        RECT 76.520 72.070 76.660 74.810 ;
        RECT 78.360 74.110 78.500 74.810 ;
        RECT 78.300 73.790 78.560 74.110 ;
        RECT 78.360 72.490 78.500 73.790 ;
        RECT 78.360 72.410 78.960 72.490 ;
        RECT 78.360 72.350 79.020 72.410 ;
        RECT 78.760 72.090 79.020 72.350 ;
        RECT 79.280 72.070 79.420 76.510 ;
        RECT 79.740 74.790 79.880 79.910 ;
        RECT 82.500 77.850 82.640 85.350 ;
        RECT 82.960 83.970 83.100 88.070 ;
        RECT 82.900 83.650 83.160 83.970 ;
        RECT 83.420 77.930 83.560 92.830 ;
        RECT 83.880 91.790 84.020 109.490 ;
        RECT 84.580 108.615 86.460 108.985 ;
        RECT 87.040 107.110 87.300 107.430 ;
        RECT 87.100 105.730 87.240 107.110 ;
        RECT 87.500 106.430 87.760 106.750 ;
        RECT 87.040 105.410 87.300 105.730 ;
        RECT 86.580 104.390 86.840 104.710 ;
        RECT 84.580 103.175 86.460 103.545 ;
        RECT 86.640 102.670 86.780 104.390 ;
        RECT 86.580 102.350 86.840 102.670 ;
        RECT 86.120 101.670 86.380 101.990 ;
        RECT 86.580 101.900 86.840 101.990 ;
        RECT 87.100 101.900 87.240 105.410 ;
        RECT 87.560 102.330 87.700 106.430 ;
        RECT 87.960 104.390 88.220 104.710 ;
        RECT 88.020 103.010 88.160 104.390 ;
        RECT 87.960 102.690 88.220 103.010 ;
        RECT 87.500 102.010 87.760 102.330 ;
        RECT 86.580 101.760 87.240 101.900 ;
        RECT 86.580 101.670 86.840 101.760 ;
        RECT 86.180 99.950 86.320 101.670 ;
        RECT 86.120 99.630 86.380 99.950 ;
        RECT 84.580 97.735 86.460 98.105 ;
        RECT 86.640 96.890 86.780 101.670 ;
        RECT 87.040 99.630 87.300 99.950 ;
        RECT 87.100 97.570 87.240 99.630 ;
        RECT 87.040 97.250 87.300 97.570 ;
        RECT 86.580 96.570 86.840 96.890 ;
        RECT 87.040 96.570 87.300 96.890 ;
        RECT 88.420 96.570 88.680 96.890 ;
        RECT 87.100 93.830 87.240 96.570 ;
        RECT 87.040 93.510 87.300 93.830 ;
        RECT 87.960 92.830 88.220 93.150 ;
        RECT 84.580 92.295 86.460 92.665 ;
        RECT 83.820 91.470 84.080 91.790 ;
        RECT 83.880 90.285 84.020 91.470 ;
        RECT 83.810 89.915 84.090 90.285 ;
        RECT 83.820 88.410 84.080 88.730 ;
        RECT 83.880 86.350 84.020 88.410 ;
        RECT 86.580 88.070 86.840 88.390 ;
        RECT 84.580 86.855 86.460 87.225 ;
        RECT 83.820 86.030 84.080 86.350 ;
        RECT 84.740 85.690 85.000 86.010 ;
        RECT 85.200 85.920 85.460 86.010 ;
        RECT 86.640 85.920 86.780 88.070 ;
        RECT 85.200 85.780 86.780 85.920 ;
        RECT 85.200 85.690 85.460 85.780 ;
        RECT 84.800 84.990 84.940 85.690 ;
        RECT 84.740 84.670 85.000 84.990 ;
        RECT 85.260 83.970 85.400 85.690 ;
        RECT 87.500 85.350 87.760 85.670 ;
        RECT 85.200 83.650 85.460 83.970 ;
        RECT 84.580 81.415 86.460 81.785 ;
        RECT 87.040 80.250 87.300 80.570 ;
        RECT 86.580 79.910 86.840 80.230 ;
        RECT 82.440 77.530 82.700 77.850 ;
        RECT 83.420 77.790 84.020 77.930 ;
        RECT 83.360 77.190 83.620 77.510 ;
        RECT 81.060 76.510 81.320 76.830 ;
        RECT 81.980 76.510 82.240 76.830 ;
        RECT 81.120 75.130 81.260 76.510 ;
        RECT 81.520 75.150 81.780 75.470 ;
        RECT 81.060 74.810 81.320 75.130 ;
        RECT 79.680 74.470 79.940 74.790 ;
        RECT 80.600 74.470 80.860 74.790 ;
        RECT 79.740 72.070 79.880 74.470 ;
        RECT 69.100 71.750 69.360 72.070 ;
        RECT 74.160 71.750 74.420 72.070 ;
        RECT 76.460 71.750 76.720 72.070 ;
        RECT 79.220 71.750 79.480 72.070 ;
        RECT 79.680 71.750 79.940 72.070 ;
        RECT 67.260 71.070 67.520 71.390 ;
        RECT 71.860 71.070 72.120 71.390 ;
        RECT 67.320 69.690 67.460 71.070 ;
        RECT 67.260 69.370 67.520 69.690 ;
        RECT 68.640 69.030 68.900 69.350 ;
        RECT 67.250 66.795 67.530 67.165 ;
        RECT 67.260 66.650 67.520 66.795 ;
        RECT 65.880 65.630 66.140 65.950 ;
        RECT 65.940 62.210 66.080 65.630 ;
        RECT 65.880 61.890 66.140 62.210 ;
        RECT 65.880 61.210 66.140 61.530 ;
        RECT 65.940 59.490 66.080 61.210 ;
        RECT 66.340 60.870 66.600 61.190 ;
        RECT 65.880 59.170 66.140 59.490 ;
        RECT 66.400 56.090 66.540 60.870 ;
        RECT 66.340 55.770 66.600 56.090 ;
        RECT 65.420 52.030 65.680 52.350 ;
        RECT 64.040 49.990 64.300 50.310 ;
        RECT 64.100 47.930 64.240 49.990 ;
        RECT 64.040 47.610 64.300 47.930 ;
        RECT 63.120 47.270 63.380 47.590 ;
        RECT 62.650 44.355 62.930 44.725 ;
        RECT 61.740 42.170 62.000 42.490 ;
        RECT 59.900 41.830 60.160 42.150 ;
        RECT 60.360 41.830 60.620 42.150 ;
        RECT 59.440 39.450 59.700 39.770 ;
        RECT 59.440 39.000 59.700 39.090 ;
        RECT 59.960 39.000 60.100 41.830 ;
        RECT 60.420 40.110 60.560 41.830 ;
        RECT 60.360 39.790 60.620 40.110 ;
        RECT 60.360 39.340 60.620 39.430 ;
        RECT 60.360 39.200 61.020 39.340 ;
        RECT 60.360 39.110 60.620 39.200 ;
        RECT 59.440 38.860 60.100 39.000 ;
        RECT 59.440 38.770 59.700 38.860 ;
        RECT 58.980 38.430 59.240 38.750 ;
        RECT 58.520 37.410 58.780 37.730 ;
        RECT 57.140 37.070 57.400 37.390 ;
        RECT 58.520 36.730 58.780 37.050 ;
        RECT 56.680 36.050 56.940 36.370 ;
        RECT 54.580 32.455 56.460 32.825 ;
        RECT 56.740 32.290 56.880 36.050 ;
        RECT 56.680 31.970 56.940 32.290 ;
        RECT 53.000 30.950 53.260 31.270 ;
        RECT 47.940 28.570 48.200 28.890 ;
        RECT 47.480 27.550 47.740 27.870 ;
        RECT 47.540 26.850 47.680 27.550 ;
        RECT 47.480 26.530 47.740 26.850 ;
        RECT 53.060 25.490 53.200 30.950 ;
        RECT 56.740 28.550 56.880 31.970 ;
        RECT 58.580 31.610 58.720 36.730 ;
        RECT 59.500 36.710 59.640 38.770 ;
        RECT 60.360 38.430 60.620 38.750 ;
        RECT 60.420 37.390 60.560 38.430 ;
        RECT 60.360 37.070 60.620 37.390 ;
        RECT 59.440 36.390 59.700 36.710 ;
        RECT 59.500 31.950 59.640 36.390 ;
        RECT 59.900 32.990 60.160 33.310 ;
        RECT 59.440 31.630 59.700 31.950 ;
        RECT 58.520 31.290 58.780 31.610 ;
        RECT 56.680 28.230 56.940 28.550 ;
        RECT 54.580 27.015 56.460 27.385 ;
        RECT 57.600 26.190 57.860 26.510 ;
        RECT 53.000 25.170 53.260 25.490 ;
        RECT 52.080 23.810 52.340 24.130 ;
        RECT 46.100 22.790 46.360 23.110 ;
        RECT 52.140 22.770 52.280 23.810 ;
        RECT 53.060 23.110 53.200 25.170 ;
        RECT 57.140 23.130 57.400 23.450 ;
        RECT 53.000 22.790 53.260 23.110 ;
        RECT 53.920 22.790 54.180 23.110 ;
        RECT 52.080 22.450 52.340 22.770 ;
        RECT 47.480 22.110 47.740 22.430 ;
        RECT 48.400 22.110 48.660 22.430 ;
        RECT 49.320 22.110 49.580 22.430 ;
        RECT 53.460 22.110 53.720 22.430 ;
        RECT 47.540 21.070 47.680 22.110 ;
        RECT 47.480 20.750 47.740 21.070 ;
        RECT 36.440 20.410 36.700 20.730 ;
        RECT 44.720 20.410 44.980 20.730 ;
        RECT 9.580 18.855 11.460 19.225 ;
        RECT 39.580 18.855 41.460 19.225 ;
        RECT 44.780 18.010 44.920 20.410 ;
        RECT 48.460 20.390 48.600 22.110 ;
        RECT 48.400 20.070 48.660 20.390 ;
        RECT 44.720 17.690 44.980 18.010 ;
        RECT 49.380 17.330 49.520 22.110 ;
        RECT 53.520 21.070 53.660 22.110 ;
        RECT 53.460 20.750 53.720 21.070 ;
        RECT 49.320 17.010 49.580 17.330 ;
        RECT 24.580 16.135 26.460 16.505 ;
        RECT 53.520 14.950 53.660 20.750 ;
        RECT 53.980 20.390 54.120 22.790 ;
        RECT 56.680 22.110 56.940 22.430 ;
        RECT 54.580 21.575 56.460 21.945 ;
        RECT 53.920 20.070 54.180 20.390 ;
        RECT 56.740 20.050 56.880 22.110 ;
        RECT 57.200 21.410 57.340 23.130 ;
        RECT 57.140 21.090 57.400 21.410 ;
        RECT 57.660 21.070 57.800 26.190 ;
        RECT 58.580 26.170 58.720 31.290 ;
        RECT 58.520 25.850 58.780 26.170 ;
        RECT 58.580 22.770 58.720 25.850 ;
        RECT 59.500 25.150 59.640 31.630 ;
        RECT 59.960 31.610 60.100 32.990 ;
        RECT 59.900 31.290 60.160 31.610 ;
        RECT 60.420 31.010 60.560 37.070 ;
        RECT 60.880 34.330 61.020 39.200 ;
        RECT 61.280 39.110 61.540 39.430 ;
        RECT 61.340 38.750 61.480 39.110 ;
        RECT 61.280 38.430 61.540 38.750 ;
        RECT 61.740 38.430 62.000 38.750 ;
        RECT 61.800 36.370 61.940 38.430 ;
        RECT 61.740 36.050 62.000 36.370 ;
        RECT 60.820 34.010 61.080 34.330 ;
        RECT 59.960 30.870 60.560 31.010 ;
        RECT 59.960 28.550 60.100 30.870 ;
        RECT 60.360 29.480 60.620 29.570 ;
        RECT 60.880 29.480 61.020 34.010 ;
        RECT 63.180 32.290 63.320 47.270 ;
        RECT 64.960 46.590 65.220 46.910 ;
        RECT 65.020 45.890 65.160 46.590 ;
        RECT 64.040 45.570 64.300 45.890 ;
        RECT 64.960 45.570 65.220 45.890 ;
        RECT 64.100 44.870 64.240 45.570 ;
        RECT 63.580 44.550 63.840 44.870 ;
        RECT 64.040 44.550 64.300 44.870 ;
        RECT 63.640 40.450 63.780 44.550 ;
        RECT 64.100 42.570 64.240 44.550 ;
        RECT 64.100 42.490 64.700 42.570 ;
        RECT 64.100 42.430 64.760 42.490 ;
        RECT 64.500 42.170 64.760 42.430 ;
        RECT 65.410 42.315 65.690 42.685 ;
        RECT 65.480 41.810 65.620 42.315 ;
        RECT 65.420 41.490 65.680 41.810 ;
        RECT 63.580 40.130 63.840 40.450 ;
        RECT 64.960 39.110 65.220 39.430 ;
        RECT 65.020 36.710 65.160 39.110 ;
        RECT 64.960 36.390 65.220 36.710 ;
        RECT 63.120 31.970 63.380 32.290 ;
        RECT 61.800 31.550 63.320 31.690 ;
        RECT 61.800 31.270 61.940 31.550 ;
        RECT 61.740 30.950 62.000 31.270 ;
        RECT 60.360 29.340 61.020 29.480 ;
        RECT 60.360 29.250 60.620 29.340 ;
        RECT 62.660 29.250 62.920 29.570 ;
        RECT 59.900 28.230 60.160 28.550 ;
        RECT 59.960 25.830 60.100 28.230 ;
        RECT 60.360 27.890 60.620 28.210 ;
        RECT 60.420 25.830 60.560 27.890 ;
        RECT 61.280 27.550 61.540 27.870 ;
        RECT 61.340 26.510 61.480 27.550 ;
        RECT 61.280 26.190 61.540 26.510 ;
        RECT 62.720 25.830 62.860 29.250 ;
        RECT 59.900 25.510 60.160 25.830 ;
        RECT 60.360 25.510 60.620 25.830 ;
        RECT 62.660 25.510 62.920 25.830 ;
        RECT 59.440 24.830 59.700 25.150 ;
        RECT 59.500 23.790 59.640 24.830 ;
        RECT 59.960 23.790 60.100 25.510 ;
        RECT 60.420 24.130 60.560 25.510 ;
        RECT 63.180 25.150 63.320 31.550 ;
        RECT 64.040 28.230 64.300 28.550 ;
        RECT 64.100 26.170 64.240 28.230 ;
        RECT 64.040 25.850 64.300 26.170 ;
        RECT 63.120 24.830 63.380 25.150 ;
        RECT 64.500 24.830 64.760 25.150 ;
        RECT 60.360 23.810 60.620 24.130 ;
        RECT 59.440 23.470 59.700 23.790 ;
        RECT 59.900 23.470 60.160 23.790 ;
        RECT 58.520 22.450 58.780 22.770 ;
        RECT 58.060 22.110 58.320 22.430 ;
        RECT 58.120 21.070 58.260 22.110 ;
        RECT 57.600 20.750 57.860 21.070 ;
        RECT 58.060 20.750 58.320 21.070 ;
        RECT 58.580 20.390 58.720 22.450 ;
        RECT 58.980 22.110 59.240 22.430 ;
        RECT 59.040 20.730 59.180 22.110 ;
        RECT 58.980 20.410 59.240 20.730 ;
        RECT 58.520 20.070 58.780 20.390 ;
        RECT 56.680 19.730 56.940 20.050 ;
        RECT 59.040 18.690 59.180 20.410 ;
        RECT 58.980 18.370 59.240 18.690 ;
        RECT 57.140 17.010 57.400 17.330 ;
        RECT 54.580 16.135 56.460 16.505 ;
        RECT 57.200 15.970 57.340 17.010 ;
        RECT 58.980 16.670 59.240 16.990 ;
        RECT 59.040 15.970 59.180 16.670 ;
        RECT 57.140 15.650 57.400 15.970 ;
        RECT 58.980 15.650 59.240 15.970 ;
        RECT 53.460 14.630 53.720 14.950 ;
        RECT 59.500 14.610 59.640 23.470 ;
        RECT 60.420 21.410 60.560 23.810 ;
        RECT 64.560 23.110 64.700 24.830 ;
        RECT 61.280 22.790 61.540 23.110 ;
        RECT 64.500 22.790 64.760 23.110 ;
        RECT 61.340 21.410 61.480 22.790 ;
        RECT 60.360 21.090 60.620 21.410 ;
        RECT 61.280 21.090 61.540 21.410 ;
        RECT 59.900 20.070 60.160 20.390 ;
        RECT 59.960 18.690 60.100 20.070 ;
        RECT 66.400 19.710 66.540 55.770 ;
        RECT 68.180 49.310 68.440 49.630 ;
        RECT 68.240 48.270 68.380 49.310 ;
        RECT 68.180 47.950 68.440 48.270 ;
        RECT 66.800 47.270 67.060 47.590 ;
        RECT 66.860 46.910 67.000 47.270 ;
        RECT 67.710 47.075 67.990 47.445 ;
        RECT 68.180 47.270 68.440 47.590 ;
        RECT 66.800 46.590 67.060 46.910 ;
        RECT 67.780 45.550 67.920 47.075 ;
        RECT 68.240 45.890 68.380 47.270 ;
        RECT 68.180 45.570 68.440 45.890 ;
        RECT 67.720 45.230 67.980 45.550 ;
        RECT 66.790 44.355 67.070 44.725 ;
        RECT 66.860 43.170 67.000 44.355 ;
        RECT 66.800 42.850 67.060 43.170 ;
        RECT 67.260 42.170 67.520 42.490 ;
        RECT 67.320 34.330 67.460 42.170 ;
        RECT 68.700 35.090 68.840 69.030 ;
        RECT 69.580 67.815 71.460 68.185 ;
        RECT 71.920 66.970 72.060 71.070 ;
        RECT 74.220 70.370 74.360 71.750 ;
        RECT 74.160 70.050 74.420 70.370 ;
        RECT 76.000 69.370 76.260 69.690 ;
        RECT 71.860 66.650 72.120 66.970 ;
        RECT 69.100 66.310 69.360 66.630 ;
        RECT 69.160 58.810 69.300 66.310 ;
        RECT 74.160 65.970 74.420 66.290 ;
        RECT 74.220 64.930 74.360 65.970 ;
        RECT 74.160 64.610 74.420 64.930 ;
        RECT 76.060 64.250 76.200 69.370 ;
        RECT 78.760 68.690 79.020 69.010 ;
        RECT 78.820 67.650 78.960 68.690 ;
        RECT 79.280 67.650 79.420 71.750 ;
        RECT 78.760 67.330 79.020 67.650 ;
        RECT 79.220 67.330 79.480 67.650 ;
        RECT 79.220 66.310 79.480 66.630 ;
        RECT 79.280 64.250 79.420 66.310 ;
        RECT 79.680 65.970 79.940 66.290 ;
        RECT 79.740 64.930 79.880 65.970 ;
        RECT 79.680 64.610 79.940 64.930 ;
        RECT 70.020 64.160 70.280 64.250 ;
        RECT 70.020 64.020 72.060 64.160 ;
        RECT 70.020 63.930 70.280 64.020 ;
        RECT 69.580 62.375 71.460 62.745 ;
        RECT 70.480 60.190 70.740 60.510 ;
        RECT 70.540 59.150 70.680 60.190 ;
        RECT 70.480 58.830 70.740 59.150 ;
        RECT 69.100 58.490 69.360 58.810 ;
        RECT 69.160 56.090 69.300 58.490 ;
        RECT 71.920 58.210 72.060 64.020 ;
        RECT 76.000 63.930 76.260 64.250 ;
        RECT 79.220 63.930 79.480 64.250 ;
        RECT 79.740 61.870 79.880 64.610 ;
        RECT 80.140 63.930 80.400 64.250 ;
        RECT 80.200 63.230 80.340 63.930 ;
        RECT 80.140 62.910 80.400 63.230 ;
        RECT 79.680 61.550 79.940 61.870 ;
        RECT 78.760 60.190 79.020 60.510 ;
        RECT 74.160 58.830 74.420 59.150 ;
        RECT 71.460 58.070 72.060 58.210 ;
        RECT 72.320 58.150 72.580 58.470 ;
        RECT 71.460 57.790 71.600 58.070 ;
        RECT 71.400 57.470 71.660 57.790 ;
        RECT 69.580 56.935 71.460 57.305 ;
        RECT 71.920 56.170 72.060 58.070 ;
        RECT 69.100 55.770 69.360 56.090 ;
        RECT 71.460 56.030 72.060 56.170 ;
        RECT 71.460 55.750 71.600 56.030 ;
        RECT 71.400 55.430 71.660 55.750 ;
        RECT 69.580 51.495 71.460 51.865 ;
        RECT 72.380 50.310 72.520 58.150 ;
        RECT 74.220 56.770 74.360 58.830 ;
        RECT 75.540 57.810 75.800 58.130 ;
        RECT 74.160 56.450 74.420 56.770 ;
        RECT 75.600 56.090 75.740 57.810 ;
        RECT 78.300 57.470 78.560 57.790 ;
        RECT 78.360 56.090 78.500 57.470 ;
        RECT 78.820 56.090 78.960 60.190 ;
        RECT 80.200 59.490 80.340 62.910 ;
        RECT 80.140 59.170 80.400 59.490 ;
        RECT 79.680 58.490 79.940 58.810 ;
        RECT 75.540 55.770 75.800 56.090 ;
        RECT 78.300 55.770 78.560 56.090 ;
        RECT 78.760 55.770 79.020 56.090 ;
        RECT 79.740 55.410 79.880 58.490 ;
        RECT 79.680 55.090 79.940 55.410 ;
        RECT 80.660 51.330 80.800 74.470 ;
        RECT 81.580 73.090 81.720 75.150 ;
        RECT 81.520 72.770 81.780 73.090 ;
        RECT 82.040 69.690 82.180 76.510 ;
        RECT 83.420 75.810 83.560 77.190 ;
        RECT 83.360 75.490 83.620 75.810 ;
        RECT 83.880 74.110 84.020 77.790 ;
        RECT 84.580 75.975 86.460 76.345 ;
        RECT 84.280 74.810 84.540 75.130 ;
        RECT 82.440 73.790 82.700 74.110 ;
        RECT 83.820 73.790 84.080 74.110 ;
        RECT 82.500 72.410 82.640 73.790 ;
        RECT 82.440 72.090 82.700 72.410 ;
        RECT 82.900 71.750 83.160 72.070 ;
        RECT 83.360 71.750 83.620 72.070 ;
        RECT 84.340 71.810 84.480 74.810 ;
        RECT 82.440 70.050 82.700 70.370 ;
        RECT 81.980 69.370 82.240 69.690 ;
        RECT 82.500 65.950 82.640 70.050 ;
        RECT 82.440 65.630 82.700 65.950 ;
        RECT 82.960 64.930 83.100 71.750 ;
        RECT 82.900 64.610 83.160 64.930 ;
        RECT 83.420 64.330 83.560 71.750 ;
        RECT 83.880 71.670 84.480 71.810 ;
        RECT 83.880 67.650 84.020 71.670 ;
        RECT 84.580 70.535 86.460 70.905 ;
        RECT 83.820 67.330 84.080 67.650 ;
        RECT 86.120 66.990 86.380 67.310 ;
        RECT 86.180 66.630 86.320 66.990 ;
        RECT 86.120 66.310 86.380 66.630 ;
        RECT 83.820 65.630 84.080 65.950 ;
        RECT 82.960 64.190 83.560 64.330 ;
        RECT 82.440 63.590 82.700 63.910 ;
        RECT 82.500 63.230 82.640 63.590 ;
        RECT 82.440 62.910 82.700 63.230 ;
        RECT 81.980 57.470 82.240 57.790 ;
        RECT 82.040 55.410 82.180 57.470 ;
        RECT 81.980 55.090 82.240 55.410 ;
        RECT 80.600 51.010 80.860 51.330 ;
        RECT 72.320 49.990 72.580 50.310 ;
        RECT 78.300 49.990 78.560 50.310 ;
        RECT 79.220 49.990 79.480 50.310 ;
        RECT 79.680 49.990 79.940 50.310 ;
        RECT 81.980 49.990 82.240 50.310 ;
        RECT 71.860 49.310 72.120 49.630 ;
        RECT 70.020 48.290 70.280 48.610 ;
        RECT 70.080 48.125 70.220 48.290 ;
        RECT 71.920 48.270 72.060 49.310 ;
        RECT 70.010 47.755 70.290 48.125 ;
        RECT 71.860 47.950 72.120 48.270 ;
        RECT 69.100 46.590 69.360 46.910 ;
        RECT 69.160 45.210 69.300 46.590 ;
        RECT 69.580 46.055 71.460 46.425 ;
        RECT 69.100 44.890 69.360 45.210 ;
        RECT 71.860 44.210 72.120 44.530 ;
        RECT 70.940 43.930 71.200 44.190 ;
        RECT 71.920 43.930 72.060 44.210 ;
        RECT 70.940 43.870 72.060 43.930 ;
        RECT 71.000 43.790 72.060 43.870 ;
        RECT 69.580 40.615 71.460 40.985 ;
        RECT 72.380 39.430 72.520 49.990 ;
        RECT 76.000 49.650 76.260 49.970 ;
        RECT 76.060 48.610 76.200 49.650 ;
        RECT 78.360 49.630 78.500 49.990 ;
        RECT 78.300 49.310 78.560 49.630 ;
        RECT 76.000 48.290 76.260 48.610 ;
        RECT 78.360 48.125 78.500 49.310 ;
        RECT 76.460 47.610 76.720 47.930 ;
        RECT 78.290 47.755 78.570 48.125 ;
        RECT 75.080 47.270 75.340 47.590 ;
        RECT 73.700 44.890 73.960 45.210 ;
        RECT 73.760 39.430 73.900 44.890 ;
        RECT 75.140 43.170 75.280 47.270 ;
        RECT 75.080 42.850 75.340 43.170 ;
        RECT 76.520 41.810 76.660 47.610 ;
        RECT 79.280 47.590 79.420 49.990 ;
        RECT 79.740 48.270 79.880 49.990 ;
        RECT 82.040 49.630 82.180 49.990 ;
        RECT 81.980 49.310 82.240 49.630 ;
        RECT 79.680 47.950 79.940 48.270 ;
        RECT 78.760 47.270 79.020 47.590 ;
        RECT 79.220 47.270 79.480 47.590 ;
        RECT 78.820 46.910 78.960 47.270 ;
        RECT 78.760 46.590 79.020 46.910 ;
        RECT 76.920 44.210 77.180 44.530 ;
        RECT 76.460 41.490 76.720 41.810 ;
        RECT 72.320 39.110 72.580 39.430 ;
        RECT 73.700 39.110 73.960 39.430 ;
        RECT 72.380 36.370 72.520 39.110 ;
        RECT 73.760 36.710 73.900 39.110 ;
        RECT 75.080 38.430 75.340 38.750 ;
        RECT 75.140 37.390 75.280 38.430 ;
        RECT 75.080 37.070 75.340 37.390 ;
        RECT 73.700 36.390 73.960 36.710 ;
        RECT 72.320 36.050 72.580 36.370 ;
        RECT 69.580 35.175 71.460 35.545 ;
        RECT 68.240 34.950 68.840 35.090 ;
        RECT 67.260 34.010 67.520 34.330 ;
        RECT 66.800 31.970 67.060 32.290 ;
        RECT 66.860 28.550 67.000 31.970 ;
        RECT 67.260 31.630 67.520 31.950 ;
        RECT 67.320 29.570 67.460 31.630 ;
        RECT 67.260 29.250 67.520 29.570 ;
        RECT 66.800 28.230 67.060 28.550 ;
        RECT 66.340 19.390 66.600 19.710 ;
        RECT 59.900 18.370 60.160 18.690 ;
        RECT 59.960 15.290 60.100 18.370 ;
        RECT 66.860 17.670 67.000 28.230 ;
        RECT 68.240 24.130 68.380 34.950 ;
        RECT 73.760 34.670 73.900 36.390 ;
        RECT 73.700 34.350 73.960 34.670 ;
        RECT 70.940 34.010 71.200 34.330 ;
        RECT 71.000 32.290 71.140 34.010 ;
        RECT 72.780 32.990 73.040 33.310 ;
        RECT 70.940 31.970 71.200 32.290 ;
        RECT 72.840 31.950 72.980 32.990 ;
        RECT 72.780 31.630 73.040 31.950 ;
        RECT 73.760 31.270 73.900 34.350 ;
        RECT 76.520 33.990 76.660 41.490 ;
        RECT 76.980 40.450 77.120 44.210 ;
        RECT 78.820 42.150 78.960 46.590 ;
        RECT 82.040 45.550 82.180 49.310 ;
        RECT 82.960 45.890 83.100 64.190 ;
        RECT 83.360 62.910 83.620 63.230 ;
        RECT 83.420 61.190 83.560 62.910 ;
        RECT 83.880 61.530 84.020 65.630 ;
        RECT 84.580 65.095 86.460 65.465 ;
        RECT 86.640 62.170 86.780 79.910 ;
        RECT 87.100 64.930 87.240 80.250 ;
        RECT 87.040 64.610 87.300 64.930 ;
        RECT 86.640 62.030 87.240 62.170 ;
        RECT 83.820 61.210 84.080 61.530 ;
        RECT 83.360 60.870 83.620 61.190 ;
        RECT 83.360 60.190 83.620 60.510 ;
        RECT 83.820 60.190 84.080 60.510 ;
        RECT 86.580 60.190 86.840 60.510 ;
        RECT 83.420 56.770 83.560 60.190 ;
        RECT 83.880 58.810 84.020 60.190 ;
        RECT 84.580 59.655 86.460 60.025 ;
        RECT 86.640 59.150 86.780 60.190 ;
        RECT 86.580 58.830 86.840 59.150 ;
        RECT 83.820 58.490 84.080 58.810 ;
        RECT 83.360 56.450 83.620 56.770 ;
        RECT 84.580 54.215 86.460 54.585 ;
        RECT 85.660 52.030 85.920 52.350 ;
        RECT 83.360 50.670 83.620 50.990 ;
        RECT 83.420 50.310 83.560 50.670 ;
        RECT 85.720 50.310 85.860 52.030 ;
        RECT 87.100 51.330 87.240 62.030 ;
        RECT 87.040 51.010 87.300 51.330 ;
        RECT 83.360 49.990 83.620 50.310 ;
        RECT 83.820 49.990 84.080 50.310 ;
        RECT 85.660 49.990 85.920 50.310 ;
        RECT 83.880 49.630 84.020 49.990 ;
        RECT 83.360 49.310 83.620 49.630 ;
        RECT 83.820 49.310 84.080 49.630 ;
        RECT 82.900 45.570 83.160 45.890 ;
        RECT 81.980 45.230 82.240 45.550 ;
        RECT 82.440 44.550 82.700 44.870 ;
        RECT 80.600 44.210 80.860 44.530 ;
        RECT 79.220 43.870 79.480 44.190 ;
        RECT 79.280 42.830 79.420 43.870 ;
        RECT 79.220 42.510 79.480 42.830 ;
        RECT 80.660 42.150 80.800 44.210 ;
        RECT 82.500 43.170 82.640 44.550 ;
        RECT 82.440 42.850 82.700 43.170 ;
        RECT 78.760 41.830 79.020 42.150 ;
        RECT 80.600 41.830 80.860 42.150 ;
        RECT 76.920 40.130 77.180 40.450 ;
        RECT 77.370 34.155 77.650 34.525 ;
        RECT 77.440 33.990 77.580 34.155 ;
        RECT 76.460 33.670 76.720 33.990 ;
        RECT 77.380 33.670 77.640 33.990 ;
        RECT 75.080 32.990 75.340 33.310 ;
        RECT 75.140 32.290 75.280 32.990 ;
        RECT 75.080 31.970 75.340 32.290 ;
        RECT 73.700 30.950 73.960 31.270 ;
        RECT 69.100 30.610 69.360 30.930 ;
        RECT 68.180 23.810 68.440 24.130 ;
        RECT 68.180 20.750 68.440 21.070 ;
        RECT 68.240 18.690 68.380 20.750 ;
        RECT 69.160 19.710 69.300 30.610 ;
        RECT 69.580 29.735 71.460 30.105 ;
        RECT 75.140 26.850 75.280 31.970 ;
        RECT 78.760 31.290 79.020 31.610 ;
        RECT 78.820 29.570 78.960 31.290 ;
        RECT 80.660 31.270 80.800 41.830 ;
        RECT 82.900 41.150 83.160 41.470 ;
        RECT 82.960 39.770 83.100 41.150 ;
        RECT 82.900 39.450 83.160 39.770 ;
        RECT 82.900 38.430 83.160 38.750 ;
        RECT 82.960 35.010 83.100 38.430 ;
        RECT 82.900 34.690 83.160 35.010 ;
        RECT 80.600 30.950 80.860 31.270 ;
        RECT 82.440 30.270 82.700 30.590 ;
        RECT 78.760 29.250 79.020 29.570 ;
        RECT 82.500 28.890 82.640 30.270 ;
        RECT 82.440 28.570 82.700 28.890 ;
        RECT 79.680 27.890 79.940 28.210 ;
        RECT 79.740 26.850 79.880 27.890 ;
        RECT 82.440 27.780 82.700 27.870 ;
        RECT 83.420 27.780 83.560 49.310 ;
        RECT 83.880 44.870 84.020 49.310 ;
        RECT 84.580 48.775 86.460 49.145 ;
        RECT 87.560 48.270 87.700 85.350 ;
        RECT 88.020 79.890 88.160 92.830 ;
        RECT 88.480 84.990 88.620 96.570 ;
        RECT 88.940 89.410 89.080 110.330 ;
        RECT 90.720 107.790 90.980 108.110 ;
        RECT 89.340 106.770 89.600 107.090 ;
        RECT 89.400 101.990 89.540 106.770 ;
        RECT 89.800 106.430 90.060 106.750 ;
        RECT 89.860 104.370 90.000 106.430 ;
        RECT 89.800 104.050 90.060 104.370 ;
        RECT 90.780 104.030 90.920 107.790 ;
        RECT 90.720 103.710 90.980 104.030 ;
        RECT 90.780 103.010 90.920 103.710 ;
        RECT 90.720 102.690 90.980 103.010 ;
        RECT 89.340 101.670 89.600 101.990 ;
        RECT 89.400 99.950 89.540 101.670 ;
        RECT 89.340 99.630 89.600 99.950 ;
        RECT 90.260 98.270 90.520 98.590 ;
        RECT 89.800 96.910 90.060 97.230 ;
        RECT 89.340 92.830 89.600 93.150 ;
        RECT 88.880 89.090 89.140 89.410 ;
        RECT 89.400 88.810 89.540 92.830 ;
        RECT 89.860 89.410 90.000 96.910 ;
        RECT 90.320 94.170 90.460 98.270 ;
        RECT 90.780 96.890 90.920 102.690 ;
        RECT 91.180 102.010 91.440 102.330 ;
        RECT 91.240 99.610 91.380 102.010 ;
        RECT 91.180 99.290 91.440 99.610 ;
        RECT 90.720 96.570 90.980 96.890 ;
        RECT 90.260 93.850 90.520 94.170 ;
        RECT 90.260 93.170 90.520 93.490 ;
        RECT 90.320 92.130 90.460 93.170 ;
        RECT 90.260 91.810 90.520 92.130 ;
        RECT 91.700 89.410 91.840 115.270 ;
        RECT 92.100 114.930 92.360 115.250 ;
        RECT 92.160 113.550 92.300 114.930 ;
        RECT 92.100 113.230 92.360 113.550 ;
        RECT 93.020 107.450 93.280 107.770 ;
        RECT 93.080 103.010 93.220 107.450 ;
        RECT 93.940 106.430 94.200 106.750 ;
        RECT 94.000 105.050 94.140 106.430 ;
        RECT 93.940 104.730 94.200 105.050 ;
        RECT 93.020 102.690 93.280 103.010 ;
        RECT 93.020 96.910 93.280 97.230 ;
        RECT 92.560 96.570 92.820 96.890 ;
        RECT 92.620 89.410 92.760 96.570 ;
        RECT 93.080 90.770 93.220 96.910 ;
        RECT 93.480 93.510 93.740 93.830 ;
        RECT 93.020 90.450 93.280 90.770 ;
        RECT 93.540 89.410 93.680 93.510 ;
        RECT 89.800 89.090 90.060 89.410 ;
        RECT 91.640 89.090 91.900 89.410 ;
        RECT 92.560 89.090 92.820 89.410 ;
        RECT 93.480 89.090 93.740 89.410 ;
        RECT 88.940 88.670 89.540 88.810 ;
        RECT 88.420 84.670 88.680 84.990 ;
        RECT 87.960 79.570 88.220 79.890 ;
        RECT 88.420 74.810 88.680 75.130 ;
        RECT 87.960 71.750 88.220 72.070 ;
        RECT 88.020 67.650 88.160 71.750 ;
        RECT 88.480 69.885 88.620 74.810 ;
        RECT 88.940 73.090 89.080 88.670 ;
        RECT 89.340 88.070 89.600 88.390 ;
        RECT 90.260 88.070 90.520 88.390 ;
        RECT 92.100 88.070 92.360 88.390 ;
        RECT 92.560 88.070 92.820 88.390 ;
        RECT 88.880 72.770 89.140 73.090 ;
        RECT 88.410 69.515 88.690 69.885 ;
        RECT 88.420 69.370 88.680 69.515 ;
        RECT 89.400 67.650 89.540 88.070 ;
        RECT 89.800 75.150 90.060 75.470 ;
        RECT 89.860 72.070 90.000 75.150 ;
        RECT 89.800 71.750 90.060 72.070 ;
        RECT 89.860 70.030 90.000 71.750 ;
        RECT 89.800 69.710 90.060 70.030 ;
        RECT 87.960 67.330 88.220 67.650 ;
        RECT 89.340 67.330 89.600 67.650 ;
        RECT 89.340 66.880 89.600 66.970 ;
        RECT 89.340 66.740 90.000 66.880 ;
        RECT 89.340 66.650 89.600 66.740 ;
        RECT 89.860 66.485 90.000 66.740 ;
        RECT 89.790 66.115 90.070 66.485 ;
        RECT 87.960 65.630 88.220 65.950 ;
        RECT 88.020 64.250 88.160 65.630 ;
        RECT 89.860 64.930 90.000 66.115 ;
        RECT 89.800 64.610 90.060 64.930 ;
        RECT 87.960 63.930 88.220 64.250 ;
        RECT 89.800 63.930 90.060 64.250 ;
        RECT 89.860 56.090 90.000 63.930 ;
        RECT 90.320 62.170 90.460 88.070 ;
        RECT 90.720 85.690 90.980 86.010 ;
        RECT 90.780 64.930 90.920 85.690 ;
        RECT 91.640 82.290 91.900 82.610 ;
        RECT 91.180 75.490 91.440 75.810 ;
        RECT 91.240 72.070 91.380 75.490 ;
        RECT 91.180 71.750 91.440 72.070 ;
        RECT 91.240 70.370 91.380 71.750 ;
        RECT 91.180 70.050 91.440 70.370 ;
        RECT 91.180 66.485 91.440 66.630 ;
        RECT 91.170 66.115 91.450 66.485 ;
        RECT 91.180 65.630 91.440 65.950 ;
        RECT 90.720 64.610 90.980 64.930 ;
        RECT 91.240 64.250 91.380 65.630 ;
        RECT 91.180 63.930 91.440 64.250 ;
        RECT 90.320 62.030 90.920 62.170 ;
        RECT 90.260 60.190 90.520 60.510 ;
        RECT 90.320 56.770 90.460 60.190 ;
        RECT 90.260 56.450 90.520 56.770 ;
        RECT 89.800 55.770 90.060 56.090 ;
        RECT 88.880 53.050 89.140 53.370 ;
        RECT 88.940 52.885 89.080 53.050 ;
        RECT 88.870 52.515 89.150 52.885 ;
        RECT 90.260 49.990 90.520 50.310 ;
        RECT 88.420 49.310 88.680 49.630 ;
        RECT 85.200 47.950 85.460 48.270 ;
        RECT 87.500 47.950 87.760 48.270 ;
        RECT 85.260 44.870 85.400 47.950 ;
        RECT 88.480 47.930 88.620 49.310 ;
        RECT 88.420 47.610 88.680 47.930 ;
        RECT 88.880 47.610 89.140 47.930 ;
        RECT 89.340 47.610 89.600 47.930 ;
        RECT 87.500 47.270 87.760 47.590 ;
        RECT 86.580 46.590 86.840 46.910 ;
        RECT 83.820 44.550 84.080 44.870 ;
        RECT 85.200 44.550 85.460 44.870 ;
        RECT 84.580 43.335 86.460 43.705 ;
        RECT 86.640 42.740 86.780 46.590 ;
        RECT 87.560 44.870 87.700 47.270 ;
        RECT 87.500 44.550 87.760 44.870 ;
        RECT 87.040 43.870 87.300 44.190 ;
        RECT 87.100 43.170 87.240 43.870 ;
        RECT 87.040 42.850 87.300 43.170 ;
        RECT 86.180 42.600 86.780 42.740 ;
        RECT 86.180 42.150 86.320 42.600 ;
        RECT 87.560 42.490 87.700 44.550 ;
        RECT 88.480 43.170 88.620 47.610 ;
        RECT 88.420 42.850 88.680 43.170 ;
        RECT 88.940 42.490 89.080 47.610 ;
        RECT 89.400 44.870 89.540 47.610 ;
        RECT 90.320 45.890 90.460 49.990 ;
        RECT 90.260 45.570 90.520 45.890 ;
        RECT 89.340 44.550 89.600 44.870 ;
        RECT 90.780 43.170 90.920 62.030 ;
        RECT 91.700 51.330 91.840 82.290 ;
        RECT 92.160 73.090 92.300 88.070 ;
        RECT 92.100 72.770 92.360 73.090 ;
        RECT 92.100 65.970 92.360 66.290 ;
        RECT 92.160 52.690 92.300 65.970 ;
        RECT 92.100 52.370 92.360 52.690 ;
        RECT 91.640 51.010 91.900 51.330 ;
        RECT 92.160 50.310 92.300 52.370 ;
        RECT 92.100 49.990 92.360 50.310 ;
        RECT 91.180 47.950 91.440 48.270 ;
        RECT 90.720 42.850 90.980 43.170 ;
        RECT 91.240 42.685 91.380 47.950 ;
        RECT 92.160 46.910 92.300 49.990 ;
        RECT 92.620 47.250 92.760 88.070 ;
        RECT 94.460 86.690 94.600 115.270 ;
        RECT 96.300 110.830 96.440 115.270 ;
        RECT 99.060 113.890 99.200 120.370 ;
        RECT 99.580 116.775 101.460 117.145 ;
        RECT 102.740 115.930 102.880 133.550 ;
        RECT 106.880 121.370 107.020 133.000 ;
        RECT 106.820 121.050 107.080 121.370 ;
        RECT 104.980 120.710 105.240 121.030 ;
        RECT 105.040 119.330 105.180 120.710 ;
        RECT 104.980 119.010 105.240 119.330 ;
        RECT 105.440 118.330 105.700 118.650 ;
        RECT 104.060 117.310 104.320 117.630 ;
        RECT 104.120 115.930 104.260 117.310 ;
        RECT 102.680 115.610 102.940 115.930 ;
        RECT 104.060 115.610 104.320 115.930 ;
        RECT 101.300 114.930 101.560 115.250 ;
        RECT 100.840 114.590 101.100 114.910 ;
        RECT 100.900 113.890 101.040 114.590 ;
        RECT 101.360 113.890 101.500 114.930 ;
        RECT 99.000 113.570 99.260 113.890 ;
        RECT 100.840 113.570 101.100 113.890 ;
        RECT 101.300 113.570 101.560 113.890 ;
        RECT 105.500 113.550 105.640 118.330 ;
        RECT 114.240 115.930 114.380 133.550 ;
        RECT 114.580 119.495 116.460 119.865 ;
        RECT 114.180 115.610 114.440 115.930 ;
        RECT 109.580 114.930 109.840 115.250 ;
        RECT 109.640 113.890 109.780 114.930 ;
        RECT 114.580 114.055 116.460 114.425 ;
        RECT 109.580 113.570 109.840 113.890 ;
        RECT 105.440 113.230 105.700 113.550 ;
        RECT 98.540 112.890 98.800 113.210 ;
        RECT 103.600 112.890 103.860 113.210 ;
        RECT 96.240 110.510 96.500 110.830 ;
        RECT 97.160 109.830 97.420 110.150 ;
        RECT 97.220 108.450 97.360 109.830 ;
        RECT 98.080 109.150 98.340 109.470 ;
        RECT 97.160 108.130 97.420 108.450 ;
        RECT 97.220 107.770 97.360 108.130 ;
        RECT 96.240 107.450 96.500 107.770 ;
        RECT 97.160 107.450 97.420 107.770 ;
        RECT 95.320 106.430 95.580 106.750 ;
        RECT 95.380 102.330 95.520 106.430 ;
        RECT 95.320 102.010 95.580 102.330 ;
        RECT 96.300 100.290 96.440 107.450 ;
        RECT 97.620 106.430 97.880 106.750 ;
        RECT 97.680 104.370 97.820 106.430 ;
        RECT 97.620 104.050 97.880 104.370 ;
        RECT 96.700 103.710 96.960 104.030 ;
        RECT 96.240 99.970 96.500 100.290 ;
        RECT 96.240 99.520 96.500 99.610 ;
        RECT 96.760 99.520 96.900 103.710 ;
        RECT 98.140 102.670 98.280 109.150 ;
        RECT 98.080 102.350 98.340 102.670 ;
        RECT 97.160 101.670 97.420 101.990 ;
        RECT 96.240 99.380 96.900 99.520 ;
        RECT 96.240 99.290 96.500 99.380 ;
        RECT 96.300 96.890 96.440 99.290 ;
        RECT 94.860 96.570 95.120 96.890 ;
        RECT 96.240 96.570 96.500 96.890 ;
        RECT 94.400 86.370 94.660 86.690 ;
        RECT 94.400 85.690 94.660 86.010 ;
        RECT 93.940 85.350 94.200 85.670 ;
        RECT 93.020 82.970 93.280 83.290 ;
        RECT 93.080 67.650 93.220 82.970 ;
        RECT 93.480 81.950 93.740 82.270 ;
        RECT 93.540 80.910 93.680 81.950 ;
        RECT 93.480 80.590 93.740 80.910 ;
        RECT 93.020 67.330 93.280 67.650 ;
        RECT 93.480 49.990 93.740 50.310 ;
        RECT 93.540 48.270 93.680 49.990 ;
        RECT 94.000 48.270 94.140 85.350 ;
        RECT 94.460 75.810 94.600 85.690 ;
        RECT 94.920 84.990 95.060 96.570 ;
        RECT 97.220 96.550 97.360 101.670 ;
        RECT 98.080 100.990 98.340 101.310 ;
        RECT 98.140 99.270 98.280 100.990 ;
        RECT 98.080 98.950 98.340 99.270 ;
        RECT 97.160 96.230 97.420 96.550 ;
        RECT 95.320 92.830 95.580 93.150 ;
        RECT 95.380 91.110 95.520 92.830 ;
        RECT 95.320 90.790 95.580 91.110 ;
        RECT 96.700 90.790 96.960 91.110 ;
        RECT 96.760 88.050 96.900 90.790 ;
        RECT 97.160 89.090 97.420 89.410 ;
        RECT 96.700 87.730 96.960 88.050 ;
        RECT 96.240 85.690 96.500 86.010 ;
        RECT 94.860 84.670 95.120 84.990 ;
        RECT 96.300 75.810 96.440 85.690 ;
        RECT 96.760 77.850 96.900 87.730 ;
        RECT 97.220 82.950 97.360 89.090 ;
        RECT 98.140 89.070 98.280 98.950 ;
        RECT 98.080 88.750 98.340 89.070 ;
        RECT 98.600 86.690 98.740 112.890 ;
        RECT 101.760 112.550 102.020 112.870 ;
        RECT 99.580 111.335 101.460 111.705 ;
        RECT 99.580 105.895 101.460 106.265 ;
        RECT 99.580 100.455 101.460 100.825 ;
        RECT 99.580 95.015 101.460 95.385 ;
        RECT 99.000 92.830 99.260 93.150 ;
        RECT 99.060 91.790 99.200 92.830 ;
        RECT 99.000 91.470 99.260 91.790 ;
        RECT 99.000 90.110 99.260 90.430 ;
        RECT 99.060 88.810 99.200 90.110 ;
        RECT 99.580 89.575 101.460 89.945 ;
        RECT 101.820 89.410 101.960 112.550 ;
        RECT 102.220 106.430 102.480 106.750 ;
        RECT 102.280 102.670 102.420 106.430 ;
        RECT 102.220 102.350 102.480 102.670 ;
        RECT 102.680 96.230 102.940 96.550 ;
        RECT 102.740 93.830 102.880 96.230 ;
        RECT 102.680 93.510 102.940 93.830 ;
        RECT 103.140 93.510 103.400 93.830 ;
        RECT 102.220 90.110 102.480 90.430 ;
        RECT 101.760 89.090 102.020 89.410 ;
        RECT 99.060 88.670 101.040 88.810 ;
        RECT 99.000 87.390 99.260 87.710 ;
        RECT 98.540 86.370 98.800 86.690 ;
        RECT 98.080 85.690 98.340 86.010 ;
        RECT 97.620 85.350 97.880 85.670 ;
        RECT 97.160 82.630 97.420 82.950 ;
        RECT 97.160 81.950 97.420 82.270 ;
        RECT 97.220 79.550 97.360 81.950 ;
        RECT 97.160 79.230 97.420 79.550 ;
        RECT 96.700 77.530 96.960 77.850 ;
        RECT 94.400 75.490 94.660 75.810 ;
        RECT 96.240 75.490 96.500 75.810 ;
        RECT 96.760 72.410 96.900 77.530 ;
        RECT 97.160 74.810 97.420 75.130 ;
        RECT 97.220 74.110 97.360 74.810 ;
        RECT 97.160 73.790 97.420 74.110 ;
        RECT 96.700 72.090 96.960 72.410 ;
        RECT 95.780 71.070 96.040 71.390 ;
        RECT 95.840 69.350 95.980 71.070 ;
        RECT 96.240 69.600 96.500 69.690 ;
        RECT 96.760 69.600 96.900 72.090 ;
        RECT 97.160 71.750 97.420 72.070 ;
        RECT 96.240 69.460 96.900 69.600 ;
        RECT 96.240 69.370 96.500 69.460 ;
        RECT 95.320 69.030 95.580 69.350 ;
        RECT 95.780 69.030 96.040 69.350 ;
        RECT 95.380 61.870 95.520 69.030 ;
        RECT 97.220 67.650 97.360 71.750 ;
        RECT 97.160 67.330 97.420 67.650 ;
        RECT 96.700 64.270 96.960 64.590 ;
        RECT 95.320 61.550 95.580 61.870 ;
        RECT 96.760 60.850 96.900 64.270 ;
        RECT 97.160 63.930 97.420 64.250 ;
        RECT 96.700 60.530 96.960 60.850 ;
        RECT 96.760 59.490 96.900 60.530 ;
        RECT 97.220 59.490 97.360 63.930 ;
        RECT 96.700 59.170 96.960 59.490 ;
        RECT 97.160 59.170 97.420 59.490 ;
        RECT 94.860 58.490 95.120 58.810 ;
        RECT 94.920 56.770 95.060 58.490 ;
        RECT 96.240 58.150 96.500 58.470 ;
        RECT 94.860 56.450 95.120 56.770 ;
        RECT 96.300 55.750 96.440 58.150 ;
        RECT 96.240 55.430 96.500 55.750 ;
        RECT 96.300 54.050 96.440 55.430 ;
        RECT 97.160 55.090 97.420 55.410 ;
        RECT 96.240 53.730 96.500 54.050 ;
        RECT 94.860 49.990 95.120 50.310 ;
        RECT 93.480 47.950 93.740 48.270 ;
        RECT 93.940 47.950 94.200 48.270 ;
        RECT 94.920 47.930 95.060 49.990 ;
        RECT 95.780 49.650 96.040 49.970 ;
        RECT 93.020 47.610 93.280 47.930 ;
        RECT 94.860 47.610 95.120 47.930 ;
        RECT 93.080 47.445 93.220 47.610 ;
        RECT 92.560 46.930 92.820 47.250 ;
        RECT 93.010 47.075 93.290 47.445 ;
        RECT 95.320 47.270 95.580 47.590 ;
        RECT 92.100 46.590 92.360 46.910 ;
        RECT 92.160 43.170 92.300 46.590 ;
        RECT 93.080 43.170 93.220 47.075 ;
        RECT 94.860 46.590 95.120 46.910 ;
        RECT 94.920 45.210 95.060 46.590 ;
        RECT 94.860 44.890 95.120 45.210 ;
        RECT 93.480 43.870 93.740 44.190 ;
        RECT 92.100 42.850 92.360 43.170 ;
        RECT 92.560 42.850 92.820 43.170 ;
        RECT 93.020 42.850 93.280 43.170 ;
        RECT 92.620 42.685 92.760 42.850 ;
        RECT 87.500 42.170 87.760 42.490 ;
        RECT 88.880 42.170 89.140 42.490 ;
        RECT 91.170 42.315 91.450 42.685 ;
        RECT 92.100 42.400 92.360 42.490 ;
        RECT 91.700 42.260 92.360 42.400 ;
        RECT 92.550 42.315 92.830 42.685 ;
        RECT 85.660 41.830 85.920 42.150 ;
        RECT 86.120 41.830 86.380 42.150 ;
        RECT 86.580 41.830 86.840 42.150 ;
        RECT 85.720 40.450 85.860 41.830 ;
        RECT 86.180 41.470 86.320 41.830 ;
        RECT 86.120 41.150 86.380 41.470 ;
        RECT 85.660 40.130 85.920 40.450 ;
        RECT 86.640 39.430 86.780 41.830 ;
        RECT 87.500 41.150 87.760 41.470 ;
        RECT 87.040 40.130 87.300 40.450 ;
        RECT 86.580 39.110 86.840 39.430 ;
        RECT 84.580 37.895 86.460 38.265 ;
        RECT 86.640 37.730 86.780 39.110 ;
        RECT 87.100 37.730 87.240 40.130 ;
        RECT 86.580 37.410 86.840 37.730 ;
        RECT 87.040 37.410 87.300 37.730 ;
        RECT 87.560 37.050 87.700 41.150 ;
        RECT 89.340 39.450 89.600 39.770 ;
        RECT 88.880 39.110 89.140 39.430 ;
        RECT 87.960 38.430 88.220 38.750 ;
        RECT 87.500 36.730 87.760 37.050 ;
        RECT 86.580 36.050 86.840 36.370 ;
        RECT 83.820 34.350 84.080 34.670 ;
        RECT 86.640 34.410 86.780 36.050 ;
        RECT 87.040 35.710 87.300 36.030 ;
        RECT 83.880 31.950 84.020 34.350 ;
        RECT 86.180 34.330 86.780 34.410 ;
        RECT 86.120 34.270 86.780 34.330 ;
        RECT 86.120 34.010 86.380 34.270 ;
        RECT 84.580 32.455 86.460 32.825 ;
        RECT 83.820 31.630 84.080 31.950 ;
        RECT 83.880 28.890 84.020 31.630 ;
        RECT 86.640 31.270 86.780 34.270 ;
        RECT 86.580 30.950 86.840 31.270 ;
        RECT 83.820 28.570 84.080 28.890 ;
        RECT 87.100 28.550 87.240 35.710 ;
        RECT 88.020 31.610 88.160 38.430 ;
        RECT 88.940 37.730 89.080 39.110 ;
        RECT 89.400 37.730 89.540 39.450 ;
        RECT 88.880 37.410 89.140 37.730 ;
        RECT 89.340 37.410 89.600 37.730 ;
        RECT 91.700 36.710 91.840 42.260 ;
        RECT 92.100 42.170 92.360 42.260 ;
        RECT 93.540 40.450 93.680 43.870 ;
        RECT 93.480 40.130 93.740 40.450 ;
        RECT 94.920 39.770 95.060 44.890 ;
        RECT 94.860 39.450 95.120 39.770 ;
        RECT 94.920 36.710 95.060 39.450 ;
        RECT 95.380 39.430 95.520 47.270 ;
        RECT 95.840 42.490 95.980 49.650 ;
        RECT 96.300 45.210 96.440 53.730 ;
        RECT 97.220 53.370 97.360 55.090 ;
        RECT 97.160 53.050 97.420 53.370 ;
        RECT 97.220 51.410 97.360 53.050 ;
        RECT 96.760 51.270 97.360 51.410 ;
        RECT 97.680 51.330 97.820 85.350 ;
        RECT 98.140 82.950 98.280 85.690 ;
        RECT 99.060 85.330 99.200 87.390 ;
        RECT 99.520 86.010 99.660 88.670 ;
        RECT 100.900 88.390 101.040 88.670 ;
        RECT 100.380 88.070 100.640 88.390 ;
        RECT 100.840 88.070 101.100 88.390 ;
        RECT 101.760 88.070 102.020 88.390 ;
        RECT 100.440 86.690 100.580 88.070 ;
        RECT 100.380 86.370 100.640 86.690 ;
        RECT 99.460 85.690 99.720 86.010 ;
        RECT 101.820 85.670 101.960 88.070 ;
        RECT 102.280 86.690 102.420 90.110 ;
        RECT 103.200 88.390 103.340 93.510 ;
        RECT 103.140 88.070 103.400 88.390 ;
        RECT 102.220 86.370 102.480 86.690 ;
        RECT 102.680 86.030 102.940 86.350 ;
        RECT 101.760 85.350 102.020 85.670 ;
        RECT 99.000 85.010 99.260 85.330 ;
        RECT 98.540 84.670 98.800 84.990 ;
        RECT 98.600 83.970 98.740 84.670 ;
        RECT 99.580 84.135 101.460 84.505 ;
        RECT 98.540 83.650 98.800 83.970 ;
        RECT 102.740 83.290 102.880 86.030 ;
        RECT 103.200 83.290 103.340 88.070 ;
        RECT 102.680 82.970 102.940 83.290 ;
        RECT 103.140 82.970 103.400 83.290 ;
        RECT 98.080 82.630 98.340 82.950 ;
        RECT 103.660 81.250 103.800 112.890 ;
        RECT 105.440 111.870 105.700 112.190 ;
        RECT 111.880 111.870 112.140 112.190 ;
        RECT 105.500 111.170 105.640 111.870 ;
        RECT 105.440 110.850 105.700 111.170 ;
        RECT 106.820 109.830 107.080 110.150 ;
        RECT 104.520 107.790 104.780 108.110 ;
        RECT 104.580 105.730 104.720 107.790 ;
        RECT 106.880 107.170 107.020 109.830 ;
        RECT 111.940 109.810 112.080 111.870 ;
        RECT 118.840 110.490 118.980 133.000 ;
        RECT 118.780 110.170 119.040 110.490 ;
        RECT 111.880 109.490 112.140 109.810 ;
        RECT 114.580 108.615 116.460 108.985 ;
        RECT 111.880 107.450 112.140 107.770 ;
        RECT 107.280 107.170 107.540 107.430 ;
        RECT 106.880 107.110 107.540 107.170 ;
        RECT 106.880 107.030 107.480 107.110 ;
        RECT 104.520 105.410 104.780 105.730 ;
        RECT 107.340 105.050 107.480 107.030 ;
        RECT 109.580 106.430 109.840 106.750 ;
        RECT 107.280 104.730 107.540 105.050 ;
        RECT 107.740 104.390 108.000 104.710 ;
        RECT 107.800 103.010 107.940 104.390 ;
        RECT 109.640 104.370 109.780 106.430 ;
        RECT 109.580 104.050 109.840 104.370 ;
        RECT 110.500 103.710 110.760 104.030 ;
        RECT 107.740 102.690 108.000 103.010 ;
        RECT 106.360 102.010 106.620 102.330 ;
        RECT 106.420 100.290 106.560 102.010 ;
        RECT 110.560 101.990 110.700 103.710 ;
        RECT 111.940 103.010 112.080 107.450 ;
        RECT 113.260 107.110 113.520 107.430 ;
        RECT 113.320 104.450 113.460 107.110 ;
        RECT 113.720 104.450 113.980 104.710 ;
        RECT 113.320 104.390 113.980 104.450 ;
        RECT 113.320 104.310 113.920 104.390 ;
        RECT 111.880 102.690 112.140 103.010 ;
        RECT 110.500 101.670 110.760 101.990 ;
        RECT 106.360 99.970 106.620 100.290 ;
        RECT 110.560 98.590 110.700 101.670 ;
        RECT 110.960 101.330 111.220 101.650 ;
        RECT 111.020 99.610 111.160 101.330 ;
        RECT 110.960 99.290 111.220 99.610 ;
        RECT 109.580 98.270 109.840 98.590 ;
        RECT 110.500 98.270 110.760 98.590 ;
        RECT 109.120 95.550 109.380 95.870 ;
        RECT 109.180 94.170 109.320 95.550 ;
        RECT 109.120 93.850 109.380 94.170 ;
        RECT 109.640 93.150 109.780 98.270 ;
        RECT 110.040 96.570 110.300 96.890 ;
        RECT 109.580 92.830 109.840 93.150 ;
        RECT 109.640 91.790 109.780 92.830 ;
        RECT 110.100 92.130 110.240 96.570 ;
        RECT 110.500 94.530 110.760 94.850 ;
        RECT 110.560 92.130 110.700 94.530 ;
        RECT 110.040 91.810 110.300 92.130 ;
        RECT 110.500 91.810 110.760 92.130 ;
        RECT 109.580 91.470 109.840 91.790 ;
        RECT 104.520 91.130 104.780 91.450 ;
        RECT 104.060 90.110 104.320 90.430 ;
        RECT 104.120 88.730 104.260 90.110 ;
        RECT 104.060 88.410 104.320 88.730 ;
        RECT 104.580 86.690 104.720 91.130 ;
        RECT 109.580 88.750 109.840 89.070 ;
        RECT 104.520 86.370 104.780 86.690 ;
        RECT 109.640 83.290 109.780 88.750 ;
        RECT 110.560 86.010 110.700 91.810 ;
        RECT 111.020 91.110 111.160 99.290 ;
        RECT 111.880 96.570 112.140 96.890 ;
        RECT 111.940 93.490 112.080 96.570 ;
        RECT 113.320 96.550 113.460 104.310 ;
        RECT 114.580 103.175 116.460 103.545 ;
        RECT 114.580 97.735 116.460 98.105 ;
        RECT 113.260 96.230 113.520 96.550 ;
        RECT 111.880 93.170 112.140 93.490 ;
        RECT 110.960 90.790 111.220 91.110 ;
        RECT 111.020 88.730 111.160 90.790 ;
        RECT 113.320 88.730 113.460 96.230 ;
        RECT 114.580 92.295 116.460 92.665 ;
        RECT 110.960 88.410 111.220 88.730 ;
        RECT 113.260 88.410 113.520 88.730 ;
        RECT 111.020 88.130 111.160 88.410 ;
        RECT 111.020 87.990 111.620 88.130 ;
        RECT 114.180 88.070 114.440 88.390 ;
        RECT 110.960 87.390 111.220 87.710 ;
        RECT 111.020 86.690 111.160 87.390 ;
        RECT 110.960 86.370 111.220 86.690 ;
        RECT 110.500 85.690 110.760 86.010 ;
        RECT 110.560 83.970 110.700 85.690 ;
        RECT 111.480 85.670 111.620 87.990 ;
        RECT 113.720 87.390 113.980 87.710 ;
        RECT 111.420 85.350 111.680 85.670 ;
        RECT 110.500 83.650 110.760 83.970 ;
        RECT 109.580 82.970 109.840 83.290 ;
        RECT 113.780 82.610 113.920 87.390 ;
        RECT 114.240 86.690 114.380 88.070 ;
        RECT 114.580 86.855 116.460 87.225 ;
        RECT 114.180 86.370 114.440 86.690 ;
        RECT 113.720 82.290 113.980 82.610 ;
        RECT 114.580 81.415 116.460 81.785 ;
        RECT 103.600 80.930 103.860 81.250 ;
        RECT 98.080 80.250 98.340 80.570 ;
        RECT 98.140 70.370 98.280 80.250 ;
        RECT 98.540 79.910 98.800 80.230 ;
        RECT 98.080 70.050 98.340 70.370 ;
        RECT 98.080 65.630 98.340 65.950 ;
        RECT 98.140 64.930 98.280 65.630 ;
        RECT 98.080 64.610 98.340 64.930 ;
        RECT 98.140 62.210 98.280 64.610 ;
        RECT 98.080 61.890 98.340 62.210 ;
        RECT 98.600 60.930 98.740 79.910 ;
        RECT 99.580 78.695 101.460 79.065 ;
        RECT 103.140 78.210 103.400 78.530 ;
        RECT 102.680 77.250 102.940 77.510 ;
        RECT 103.200 77.250 103.340 78.210 ;
        RECT 104.060 77.530 104.320 77.850 ;
        RECT 102.680 77.190 103.340 77.250 ;
        RECT 102.740 77.110 103.340 77.190 ;
        RECT 101.760 74.810 102.020 75.130 ;
        RECT 99.000 74.470 99.260 74.790 ;
        RECT 99.060 66.970 99.200 74.470 ;
        RECT 99.580 73.255 101.460 73.625 ;
        RECT 101.820 71.730 101.960 74.810 ;
        RECT 103.200 72.070 103.340 77.110 ;
        RECT 104.120 75.810 104.260 77.530 ;
        RECT 110.040 76.510 110.300 76.830 ;
        RECT 112.800 76.510 113.060 76.830 ;
        RECT 104.060 75.490 104.320 75.810 ;
        RECT 104.520 75.490 104.780 75.810 ;
        RECT 104.580 74.450 104.720 75.490 ;
        RECT 110.100 75.470 110.240 76.510 ;
        RECT 110.500 75.490 110.760 75.810 ;
        RECT 110.040 75.150 110.300 75.470 ;
        RECT 104.520 74.130 104.780 74.450 ;
        RECT 108.200 73.790 108.460 74.110 ;
        RECT 108.260 72.410 108.400 73.790 ;
        RECT 110.560 72.410 110.700 75.490 ;
        RECT 111.880 74.470 112.140 74.790 ;
        RECT 108.200 72.090 108.460 72.410 ;
        RECT 110.500 72.090 110.760 72.410 ;
        RECT 103.140 71.750 103.400 72.070 ;
        RECT 101.760 71.410 102.020 71.730 ;
        RECT 99.460 71.070 99.720 71.390 ;
        RECT 99.520 70.030 99.660 71.070 ;
        RECT 101.820 70.370 101.960 71.410 ;
        RECT 101.760 70.050 102.020 70.370 ;
        RECT 99.460 69.710 99.720 70.030 ;
        RECT 99.580 67.815 101.460 68.185 ;
        RECT 100.840 66.990 101.100 67.310 ;
        RECT 99.000 66.650 99.260 66.970 ;
        RECT 99.460 66.310 99.720 66.630 ;
        RECT 99.520 65.950 99.660 66.310 ;
        RECT 99.460 65.630 99.720 65.950 ;
        RECT 100.900 64.250 101.040 66.990 ;
        RECT 101.820 66.630 101.960 70.050 ;
        RECT 102.220 66.650 102.480 66.970 ;
        RECT 101.760 66.310 102.020 66.630 ;
        RECT 100.840 63.930 101.100 64.250 ;
        RECT 102.280 63.570 102.420 66.650 ;
        RECT 103.200 63.910 103.340 71.750 ;
        RECT 110.560 70.370 110.700 72.090 ;
        RECT 110.500 70.050 110.760 70.370 ;
        RECT 111.940 69.350 112.080 74.470 ;
        RECT 112.860 71.730 113.000 76.510 ;
        RECT 114.580 75.975 116.460 76.345 ;
        RECT 112.800 71.410 113.060 71.730 ;
        RECT 114.580 70.535 116.460 70.905 ;
        RECT 110.960 69.030 111.220 69.350 ;
        RECT 111.880 69.030 112.140 69.350 ;
        RECT 105.440 68.350 105.700 68.670 ;
        RECT 105.500 66.630 105.640 68.350 ;
        RECT 105.440 66.310 105.700 66.630 ;
        RECT 105.900 66.310 106.160 66.630 ;
        RECT 103.140 63.590 103.400 63.910 ;
        RECT 102.220 63.250 102.480 63.570 ;
        RECT 101.760 62.910 102.020 63.230 ;
        RECT 99.580 62.375 101.460 62.745 ;
        RECT 99.000 61.890 99.260 62.210 ;
        RECT 99.060 61.190 99.200 61.890 ;
        RECT 98.140 60.790 98.740 60.930 ;
        RECT 99.000 60.870 99.260 61.190 ;
        RECT 101.820 60.850 101.960 62.910 ;
        RECT 102.280 61.530 102.420 63.250 ;
        RECT 102.220 61.210 102.480 61.530 ;
        RECT 105.960 61.190 106.100 66.310 ;
        RECT 111.020 65.950 111.160 69.030 ;
        RECT 110.960 65.630 111.220 65.950 ;
        RECT 111.020 64.930 111.160 65.630 ;
        RECT 110.960 64.610 111.220 64.930 ;
        RECT 111.940 63.910 112.080 69.030 ;
        RECT 113.720 65.970 113.980 66.290 ;
        RECT 113.780 64.930 113.920 65.970 ;
        RECT 114.580 65.095 116.460 65.465 ;
        RECT 113.720 64.610 113.980 64.930 ;
        RECT 111.420 63.590 111.680 63.910 ;
        RECT 111.880 63.590 112.140 63.910 ;
        RECT 107.280 62.910 107.540 63.230 ;
        RECT 107.340 61.530 107.480 62.910 ;
        RECT 111.480 62.210 111.620 63.590 ;
        RECT 114.180 62.910 114.440 63.230 ;
        RECT 111.420 61.890 111.680 62.210 ;
        RECT 107.280 61.210 107.540 61.530 ;
        RECT 104.060 60.870 104.320 61.190 ;
        RECT 105.900 60.870 106.160 61.190 ;
        RECT 96.240 44.890 96.500 45.210 ;
        RECT 96.300 43.170 96.440 44.890 ;
        RECT 96.240 42.850 96.500 43.170 ;
        RECT 95.780 42.170 96.040 42.490 ;
        RECT 95.320 39.110 95.580 39.430 ;
        RECT 95.380 37.390 95.520 39.110 ;
        RECT 95.320 37.070 95.580 37.390 ;
        RECT 91.640 36.390 91.900 36.710 ;
        RECT 94.860 36.390 95.120 36.710 ;
        RECT 88.420 36.050 88.680 36.370 ;
        RECT 88.480 34.330 88.620 36.050 ;
        RECT 88.420 34.010 88.680 34.330 ;
        RECT 87.960 31.290 88.220 31.610 ;
        RECT 91.700 31.270 91.840 36.390 ;
        RECT 93.940 35.710 94.200 36.030 ;
        RECT 94.000 31.950 94.140 35.710 ;
        RECT 95.380 35.010 95.520 37.070 ;
        RECT 96.760 37.050 96.900 51.270 ;
        RECT 97.620 51.010 97.880 51.330 ;
        RECT 97.160 50.330 97.420 50.650 ;
        RECT 97.220 39.430 97.360 50.330 ;
        RECT 97.620 49.310 97.880 49.630 ;
        RECT 97.680 45.210 97.820 49.310 ;
        RECT 97.620 44.890 97.880 45.210 ;
        RECT 98.140 42.830 98.280 60.790 ;
        RECT 101.760 60.530 102.020 60.850 ;
        RECT 98.540 60.190 98.800 60.510 ;
        RECT 103.140 60.190 103.400 60.510 ;
        RECT 98.600 55.750 98.740 60.190 ;
        RECT 99.000 58.490 99.260 58.810 ;
        RECT 98.540 55.430 98.800 55.750 ;
        RECT 99.060 54.050 99.200 58.490 ;
        RECT 99.580 56.935 101.460 57.305 ;
        RECT 103.200 56.430 103.340 60.190 ;
        RECT 104.120 59.150 104.260 60.870 ;
        RECT 114.240 60.850 114.380 62.910 ;
        RECT 114.180 60.530 114.440 60.850 ;
        RECT 106.360 60.190 106.620 60.510 ;
        RECT 104.060 58.830 104.320 59.150 ;
        RECT 104.120 58.470 104.260 58.830 ;
        RECT 106.420 58.810 106.560 60.190 ;
        RECT 114.580 59.655 116.460 60.025 ;
        RECT 105.900 58.490 106.160 58.810 ;
        RECT 106.360 58.490 106.620 58.810 ;
        RECT 104.060 58.150 104.320 58.470 ;
        RECT 104.520 58.150 104.780 58.470 ;
        RECT 104.580 56.770 104.720 58.150 ;
        RECT 104.520 56.450 104.780 56.770 ;
        RECT 103.140 56.110 103.400 56.430 ;
        RECT 105.960 56.090 106.100 58.490 ;
        RECT 108.200 57.470 108.460 57.790 ;
        RECT 105.900 55.770 106.160 56.090 ;
        RECT 108.260 55.410 108.400 57.470 ;
        RECT 103.140 55.090 103.400 55.410 ;
        RECT 108.200 55.090 108.460 55.410 ;
        RECT 103.200 54.050 103.340 55.090 ;
        RECT 114.580 54.215 116.460 54.585 ;
        RECT 99.000 53.730 99.260 54.050 ;
        RECT 103.140 53.730 103.400 54.050 ;
        RECT 102.680 53.050 102.940 53.370 ;
        RECT 99.580 51.495 101.460 51.865 ;
        RECT 99.000 47.950 99.260 48.270 ;
        RECT 98.540 47.610 98.800 47.930 ;
        RECT 98.600 45.890 98.740 47.610 ;
        RECT 98.540 45.570 98.800 45.890 ;
        RECT 99.060 42.830 99.200 47.950 ;
        RECT 99.580 46.055 101.460 46.425 ;
        RECT 102.740 45.210 102.880 53.050 ;
        RECT 114.580 48.775 116.460 49.145 ;
        RECT 104.980 47.950 105.240 48.270 ;
        RECT 105.040 45.890 105.180 47.950 ;
        RECT 106.820 46.590 107.080 46.910 ;
        RECT 104.980 45.570 105.240 45.890 ;
        RECT 102.680 44.890 102.940 45.210 ;
        RECT 105.440 43.870 105.700 44.190 ;
        RECT 105.500 42.830 105.640 43.870 ;
        RECT 106.880 42.830 107.020 46.590 ;
        RECT 114.580 43.335 116.460 43.705 ;
        RECT 98.080 42.510 98.340 42.830 ;
        RECT 99.000 42.510 99.260 42.830 ;
        RECT 105.440 42.510 105.700 42.830 ;
        RECT 106.820 42.510 107.080 42.830 ;
        RECT 97.160 39.110 97.420 39.430 ;
        RECT 99.060 39.090 99.200 42.510 ;
        RECT 99.580 40.615 101.460 40.985 ;
        RECT 103.140 39.110 103.400 39.430 ;
        RECT 99.000 38.770 99.260 39.090 ;
        RECT 102.680 38.430 102.940 38.750 ;
        RECT 102.740 37.730 102.880 38.430 ;
        RECT 103.200 37.730 103.340 39.110 ;
        RECT 110.040 38.430 110.300 38.750 ;
        RECT 102.680 37.410 102.940 37.730 ;
        RECT 103.140 37.410 103.400 37.730 ;
        RECT 104.520 37.070 104.780 37.390 ;
        RECT 96.700 36.730 96.960 37.050 ;
        RECT 95.320 34.690 95.580 35.010 ;
        RECT 96.760 34.330 96.900 36.730 ;
        RECT 99.580 35.175 101.460 35.545 ;
        RECT 104.580 34.330 104.720 37.070 ;
        RECT 110.100 36.710 110.240 38.430 ;
        RECT 114.580 37.895 116.460 38.265 ;
        RECT 110.040 36.390 110.300 36.710 ;
        RECT 96.700 34.010 96.960 34.330 ;
        RECT 104.520 34.010 104.780 34.330 ;
        RECT 114.580 32.455 116.460 32.825 ;
        RECT 93.940 31.630 94.200 31.950 ;
        RECT 91.640 30.950 91.900 31.270 ;
        RECT 99.580 29.735 101.460 30.105 ;
        RECT 87.040 28.230 87.300 28.550 ;
        RECT 83.820 27.890 84.080 28.210 ;
        RECT 82.440 27.640 83.560 27.780 ;
        RECT 82.440 27.550 82.700 27.640 ;
        RECT 75.080 26.530 75.340 26.850 ;
        RECT 79.680 26.530 79.940 26.850 ;
        RECT 82.500 25.830 82.640 27.550 ;
        RECT 83.880 26.170 84.020 27.890 ;
        RECT 84.580 27.015 86.460 27.385 ;
        RECT 114.580 27.015 116.460 27.385 ;
        RECT 83.820 25.850 84.080 26.170 ;
        RECT 82.440 25.510 82.700 25.830 ;
        RECT 69.580 24.295 71.460 24.665 ;
        RECT 99.580 24.295 101.460 24.665 ;
        RECT 71.860 22.110 72.120 22.430 ;
        RECT 71.920 20.390 72.060 22.110 ;
        RECT 84.580 21.575 86.460 21.945 ;
        RECT 114.580 21.575 116.460 21.945 ;
        RECT 71.860 20.070 72.120 20.390 ;
        RECT 69.100 19.390 69.360 19.710 ;
        RECT 68.180 18.370 68.440 18.690 ;
        RECT 69.160 18.010 69.300 19.390 ;
        RECT 69.580 18.855 71.460 19.225 ;
        RECT 99.580 18.855 101.460 19.225 ;
        RECT 69.100 17.690 69.360 18.010 ;
        RECT 66.800 17.350 67.060 17.670 ;
        RECT 66.860 15.290 67.000 17.350 ;
        RECT 84.580 16.135 86.460 16.505 ;
        RECT 114.580 16.135 116.460 16.505 ;
        RECT 59.900 14.970 60.160 15.290 ;
        RECT 66.800 14.970 67.060 15.290 ;
        RECT 59.440 14.290 59.700 14.610 ;
        RECT 9.580 13.415 11.460 13.785 ;
        RECT 39.580 13.415 41.460 13.785 ;
        RECT 69.580 13.415 71.460 13.785 ;
        RECT 99.580 13.415 101.460 13.785 ;
        RECT 24.580 10.695 26.460 11.065 ;
        RECT 54.580 10.695 56.460 11.065 ;
        RECT 84.580 10.695 86.460 11.065 ;
        RECT 114.580 10.695 116.460 11.065 ;
      LAYER met3 ;
        RECT 9.530 122.235 11.510 122.565 ;
        RECT 39.530 122.235 41.510 122.565 ;
        RECT 69.530 122.235 71.510 122.565 ;
        RECT 99.530 122.235 101.510 122.565 ;
        RECT 24.530 119.515 26.510 119.845 ;
        RECT 54.530 119.515 56.510 119.845 ;
        RECT 84.530 119.515 86.510 119.845 ;
        RECT 114.530 119.515 116.510 119.845 ;
        RECT 9.530 116.795 11.510 117.125 ;
        RECT 39.530 116.795 41.510 117.125 ;
        RECT 69.530 116.795 71.510 117.125 ;
        RECT 99.530 116.795 101.510 117.125 ;
        RECT 6.965 116.090 7.295 116.105 ;
        RECT 2.000 115.790 7.295 116.090 ;
        RECT 6.965 115.775 7.295 115.790 ;
        RECT 24.530 114.075 26.510 114.405 ;
        RECT 54.530 114.075 56.510 114.405 ;
        RECT 84.530 114.075 86.510 114.405 ;
        RECT 114.530 114.075 116.510 114.405 ;
        RECT 9.530 111.355 11.510 111.685 ;
        RECT 39.530 111.355 41.510 111.685 ;
        RECT 69.530 111.355 71.510 111.685 ;
        RECT 99.530 111.355 101.510 111.685 ;
        RECT 37.990 109.290 38.370 109.300 ;
        RECT 40.085 109.290 40.415 109.305 ;
        RECT 37.990 108.990 40.415 109.290 ;
        RECT 37.990 108.980 38.370 108.990 ;
        RECT 40.085 108.975 40.415 108.990 ;
        RECT 24.530 108.635 26.510 108.965 ;
        RECT 54.530 108.635 56.510 108.965 ;
        RECT 84.530 108.635 86.510 108.965 ;
        RECT 114.530 108.635 116.510 108.965 ;
        RECT 9.530 105.915 11.510 106.245 ;
        RECT 39.530 105.915 41.510 106.245 ;
        RECT 69.530 105.915 71.510 106.245 ;
        RECT 99.530 105.915 101.510 106.245 ;
        RECT 24.530 103.195 26.510 103.525 ;
        RECT 54.530 103.195 56.510 103.525 ;
        RECT 84.530 103.195 86.510 103.525 ;
        RECT 114.530 103.195 116.510 103.525 ;
        RECT 9.530 100.475 11.510 100.805 ;
        RECT 39.530 100.475 41.510 100.805 ;
        RECT 69.530 100.475 71.510 100.805 ;
        RECT 99.530 100.475 101.510 100.805 ;
        RECT 24.530 97.755 26.510 98.085 ;
        RECT 54.530 97.755 56.510 98.085 ;
        RECT 84.530 97.755 86.510 98.085 ;
        RECT 114.530 97.755 116.510 98.085 ;
        RECT 9.530 95.035 11.510 95.365 ;
        RECT 39.530 95.035 41.510 95.365 ;
        RECT 69.530 95.035 71.510 95.365 ;
        RECT 99.530 95.035 101.510 95.365 ;
        RECT 37.325 92.970 37.655 92.985 ;
        RECT 37.990 92.970 38.370 92.980 ;
        RECT 37.325 92.670 38.370 92.970 ;
        RECT 37.325 92.655 37.655 92.670 ;
        RECT 37.990 92.660 38.370 92.670 ;
        RECT 24.530 92.315 26.510 92.645 ;
        RECT 54.530 92.315 56.510 92.645 ;
        RECT 84.530 92.315 86.510 92.645 ;
        RECT 114.530 92.315 116.510 92.645 ;
        RECT 83.785 90.250 84.115 90.265 ;
        RECT 88.590 90.250 88.970 90.260 ;
        RECT 83.785 89.950 88.970 90.250 ;
        RECT 83.785 89.935 84.115 89.950 ;
        RECT 88.590 89.940 88.970 89.950 ;
        RECT 9.530 89.595 11.510 89.925 ;
        RECT 39.530 89.595 41.510 89.925 ;
        RECT 69.530 89.595 71.510 89.925 ;
        RECT 99.530 89.595 101.510 89.925 ;
        RECT 24.905 88.210 25.235 88.225 ;
        RECT 33.645 88.210 33.975 88.225 ;
        RECT 24.905 87.910 33.975 88.210 ;
        RECT 24.905 87.895 25.235 87.910 ;
        RECT 33.645 87.895 33.975 87.910 ;
        RECT 24.530 86.875 26.510 87.205 ;
        RECT 54.530 86.875 56.510 87.205 ;
        RECT 84.530 86.875 86.510 87.205 ;
        RECT 114.530 86.875 116.510 87.205 ;
        RECT 9.530 84.155 11.510 84.485 ;
        RECT 39.530 84.155 41.510 84.485 ;
        RECT 69.530 84.155 71.510 84.485 ;
        RECT 99.530 84.155 101.510 84.485 ;
        RECT 20.510 83.450 20.890 83.460 ;
        RECT 2.000 83.150 20.890 83.450 ;
        RECT 20.510 83.140 20.890 83.150 ;
        RECT 24.530 81.435 26.510 81.765 ;
        RECT 54.530 81.435 56.510 81.765 ;
        RECT 84.530 81.435 86.510 81.765 ;
        RECT 114.530 81.435 116.510 81.765 ;
        RECT 9.530 78.715 11.510 79.045 ;
        RECT 39.530 78.715 41.510 79.045 ;
        RECT 69.530 78.715 71.510 79.045 ;
        RECT 99.530 78.715 101.510 79.045 ;
        RECT 24.530 75.995 26.510 76.325 ;
        RECT 54.530 75.995 56.510 76.325 ;
        RECT 84.530 75.995 86.510 76.325 ;
        RECT 114.530 75.995 116.510 76.325 ;
        RECT 9.530 73.275 11.510 73.605 ;
        RECT 39.530 73.275 41.510 73.605 ;
        RECT 69.530 73.275 71.510 73.605 ;
        RECT 99.530 73.275 101.510 73.605 ;
        RECT 25.365 71.890 25.695 71.905 ;
        RECT 33.645 71.890 33.975 71.905 ;
        RECT 45.145 71.890 45.475 71.905 ;
        RECT 25.365 71.590 45.475 71.890 ;
        RECT 25.365 71.575 25.695 71.590 ;
        RECT 33.645 71.575 33.975 71.590 ;
        RECT 45.145 71.575 45.475 71.590 ;
        RECT 24.530 70.555 26.510 70.885 ;
        RECT 54.530 70.555 56.510 70.885 ;
        RECT 84.530 70.555 86.510 70.885 ;
        RECT 114.530 70.555 116.510 70.885 ;
        RECT 64.925 69.850 65.255 69.865 ;
        RECT 88.385 69.850 88.715 69.865 ;
        RECT 64.925 69.550 88.715 69.850 ;
        RECT 64.925 69.535 65.255 69.550 ;
        RECT 88.385 69.535 88.715 69.550 ;
        RECT 9.530 67.835 11.510 68.165 ;
        RECT 39.530 67.835 41.510 68.165 ;
        RECT 69.530 67.835 71.510 68.165 ;
        RECT 99.530 67.835 101.510 68.165 ;
        RECT 20.510 67.130 20.890 67.140 ;
        RECT 58.485 67.130 58.815 67.145 ;
        RECT 67.225 67.130 67.555 67.145 ;
        RECT 88.590 67.130 88.970 67.140 ;
        RECT 20.510 66.830 58.815 67.130 ;
        RECT 20.510 66.820 20.890 66.830 ;
        RECT 58.485 66.815 58.815 66.830 ;
        RECT 61.950 66.830 88.970 67.130 ;
        RECT 37.990 66.450 38.370 66.460 ;
        RECT 61.950 66.450 62.250 66.830 ;
        RECT 67.225 66.815 67.555 66.830 ;
        RECT 88.590 66.820 88.970 66.830 ;
        RECT 37.990 66.150 62.250 66.450 ;
        RECT 89.765 66.450 90.095 66.465 ;
        RECT 91.145 66.450 91.475 66.465 ;
        RECT 89.765 66.150 91.475 66.450 ;
        RECT 37.990 66.140 38.370 66.150 ;
        RECT 89.765 66.135 90.095 66.150 ;
        RECT 91.145 66.135 91.475 66.150 ;
        RECT 57.565 65.770 57.895 65.785 ;
        RECT 59.865 65.770 60.195 65.785 ;
        RECT 57.565 65.470 60.195 65.770 ;
        RECT 57.565 65.455 57.895 65.470 ;
        RECT 59.865 65.455 60.195 65.470 ;
        RECT 24.530 65.115 26.510 65.445 ;
        RECT 54.530 65.115 56.510 65.445 ;
        RECT 84.530 65.115 86.510 65.445 ;
        RECT 114.530 65.115 116.510 65.445 ;
        RECT 48.365 63.730 48.695 63.745 ;
        RECT 61.245 63.730 61.575 63.745 ;
        RECT 64.925 63.730 65.255 63.745 ;
        RECT 48.365 63.430 65.255 63.730 ;
        RECT 48.365 63.415 48.695 63.430 ;
        RECT 61.245 63.415 61.575 63.430 ;
        RECT 64.925 63.415 65.255 63.430 ;
        RECT 51.585 63.050 51.915 63.065 ;
        RECT 52.965 63.050 53.295 63.065 ;
        RECT 51.585 62.750 53.295 63.050 ;
        RECT 51.585 62.735 51.915 62.750 ;
        RECT 52.965 62.735 53.295 62.750 ;
        RECT 9.530 62.395 11.510 62.725 ;
        RECT 39.530 62.395 41.510 62.725 ;
        RECT 69.530 62.395 71.510 62.725 ;
        RECT 99.530 62.395 101.510 62.725 ;
        RECT 24.530 59.675 26.510 60.005 ;
        RECT 54.530 59.675 56.510 60.005 ;
        RECT 84.530 59.675 86.510 60.005 ;
        RECT 114.530 59.675 116.510 60.005 ;
        RECT 31.805 58.290 32.135 58.305 ;
        RECT 34.310 58.290 34.690 58.300 ;
        RECT 37.990 58.290 38.370 58.300 ;
        RECT 31.805 57.990 38.370 58.290 ;
        RECT 31.805 57.975 32.135 57.990 ;
        RECT 34.310 57.980 34.690 57.990 ;
        RECT 37.990 57.980 38.370 57.990 ;
        RECT 9.530 56.955 11.510 57.285 ;
        RECT 39.530 56.955 41.510 57.285 ;
        RECT 69.530 56.955 71.510 57.285 ;
        RECT 99.530 56.955 101.510 57.285 ;
        RECT 24.530 54.235 26.510 54.565 ;
        RECT 54.530 54.235 56.510 54.565 ;
        RECT 84.530 54.235 86.510 54.565 ;
        RECT 114.530 54.235 116.510 54.565 ;
        RECT 88.845 52.860 89.175 52.865 ;
        RECT 88.590 52.850 89.175 52.860 ;
        RECT 88.590 52.550 89.400 52.850 ;
        RECT 88.590 52.540 89.175 52.550 ;
        RECT 88.845 52.535 89.175 52.540 ;
        RECT 9.530 51.515 11.510 51.845 ;
        RECT 39.530 51.515 41.510 51.845 ;
        RECT 69.530 51.515 71.510 51.845 ;
        RECT 99.530 51.515 101.510 51.845 ;
        RECT 5.125 50.810 5.455 50.825 ;
        RECT 2.000 50.510 5.455 50.810 ;
        RECT 5.125 50.495 5.455 50.510 ;
        RECT 24.530 48.795 26.510 49.125 ;
        RECT 54.530 48.795 56.510 49.125 ;
        RECT 84.530 48.795 86.510 49.125 ;
        RECT 114.530 48.795 116.510 49.125 ;
        RECT 69.985 48.090 70.315 48.105 ;
        RECT 78.265 48.090 78.595 48.105 ;
        RECT 69.985 47.790 78.595 48.090 ;
        RECT 69.985 47.775 70.315 47.790 ;
        RECT 78.265 47.775 78.595 47.790 ;
        RECT 67.685 47.410 68.015 47.425 ;
        RECT 92.985 47.410 93.315 47.425 ;
        RECT 67.685 47.110 93.315 47.410 ;
        RECT 67.685 47.095 68.015 47.110 ;
        RECT 92.985 47.095 93.315 47.110 ;
        RECT 9.530 46.075 11.510 46.405 ;
        RECT 39.530 46.075 41.510 46.405 ;
        RECT 69.530 46.075 71.510 46.405 ;
        RECT 99.530 46.075 101.510 46.405 ;
        RECT 54.805 45.370 55.135 45.385 ;
        RECT 61.245 45.370 61.575 45.385 ;
        RECT 54.805 45.070 61.575 45.370 ;
        RECT 54.805 45.055 55.135 45.070 ;
        RECT 61.245 45.055 61.575 45.070 ;
        RECT 60.325 44.690 60.655 44.705 ;
        RECT 62.625 44.690 62.955 44.705 ;
        RECT 66.765 44.690 67.095 44.705 ;
        RECT 60.325 44.390 67.095 44.690 ;
        RECT 60.325 44.375 60.655 44.390 ;
        RECT 62.625 44.375 62.955 44.390 ;
        RECT 66.765 44.375 67.095 44.390 ;
        RECT 24.530 43.355 26.510 43.685 ;
        RECT 54.530 43.355 56.510 43.685 ;
        RECT 84.530 43.355 86.510 43.685 ;
        RECT 114.530 43.355 116.510 43.685 ;
        RECT 47.905 42.650 48.235 42.665 ;
        RECT 54.345 42.650 54.675 42.665 ;
        RECT 47.905 42.350 54.675 42.650 ;
        RECT 47.905 42.335 48.235 42.350 ;
        RECT 54.345 42.335 54.675 42.350 ;
        RECT 65.385 42.650 65.715 42.665 ;
        RECT 91.145 42.650 91.475 42.665 ;
        RECT 92.525 42.650 92.855 42.665 ;
        RECT 65.385 42.350 92.855 42.650 ;
        RECT 65.385 42.335 65.715 42.350 ;
        RECT 91.145 42.335 91.475 42.350 ;
        RECT 92.525 42.335 92.855 42.350 ;
        RECT 9.530 40.635 11.510 40.965 ;
        RECT 39.530 40.635 41.510 40.965 ;
        RECT 69.530 40.635 71.510 40.965 ;
        RECT 99.530 40.635 101.510 40.965 ;
        RECT 24.530 37.915 26.510 38.245 ;
        RECT 54.530 37.915 56.510 38.245 ;
        RECT 84.530 37.915 86.510 38.245 ;
        RECT 114.530 37.915 116.510 38.245 ;
        RECT 9.530 35.195 11.510 35.525 ;
        RECT 39.530 35.195 41.510 35.525 ;
        RECT 69.530 35.195 71.510 35.525 ;
        RECT 99.530 35.195 101.510 35.525 ;
        RECT 34.310 34.490 34.690 34.500 ;
        RECT 38.245 34.490 38.575 34.505 ;
        RECT 34.310 34.190 38.575 34.490 ;
        RECT 34.310 34.180 34.690 34.190 ;
        RECT 38.245 34.175 38.575 34.190 ;
        RECT 77.345 34.490 77.675 34.505 ;
        RECT 88.590 34.490 88.970 34.500 ;
        RECT 77.345 34.190 88.970 34.490 ;
        RECT 77.345 34.175 77.675 34.190 ;
        RECT 88.590 34.180 88.970 34.190 ;
        RECT 24.530 32.475 26.510 32.805 ;
        RECT 54.530 32.475 56.510 32.805 ;
        RECT 84.530 32.475 86.510 32.805 ;
        RECT 114.530 32.475 116.510 32.805 ;
        RECT 9.530 29.755 11.510 30.085 ;
        RECT 39.530 29.755 41.510 30.085 ;
        RECT 69.530 29.755 71.510 30.085 ;
        RECT 99.530 29.755 101.510 30.085 ;
        RECT 24.530 27.035 26.510 27.365 ;
        RECT 54.530 27.035 56.510 27.365 ;
        RECT 84.530 27.035 86.510 27.365 ;
        RECT 114.530 27.035 116.510 27.365 ;
        RECT 9.530 24.315 11.510 24.645 ;
        RECT 39.530 24.315 41.510 24.645 ;
        RECT 69.530 24.315 71.510 24.645 ;
        RECT 99.530 24.315 101.510 24.645 ;
        RECT 24.530 21.595 26.510 21.925 ;
        RECT 54.530 21.595 56.510 21.925 ;
        RECT 84.530 21.595 86.510 21.925 ;
        RECT 114.530 21.595 116.510 21.925 ;
        RECT 9.530 18.875 11.510 19.205 ;
        RECT 39.530 18.875 41.510 19.205 ;
        RECT 69.530 18.875 71.510 19.205 ;
        RECT 99.530 18.875 101.510 19.205 ;
        RECT 24.530 16.155 26.510 16.485 ;
        RECT 54.530 16.155 56.510 16.485 ;
        RECT 84.530 16.155 86.510 16.485 ;
        RECT 114.530 16.155 116.510 16.485 ;
        RECT 9.530 13.435 11.510 13.765 ;
        RECT 39.530 13.435 41.510 13.765 ;
        RECT 69.530 13.435 71.510 13.765 ;
        RECT 99.530 13.435 101.510 13.765 ;
        RECT 24.530 10.715 26.510 11.045 ;
        RECT 54.530 10.715 56.510 11.045 ;
        RECT 84.530 10.715 86.510 11.045 ;
        RECT 114.530 10.715 116.510 11.045 ;
      LAYER met4 ;
        RECT 38.015 108.975 38.345 109.305 ;
        RECT 38.030 92.985 38.330 108.975 ;
        RECT 38.015 92.655 38.345 92.985 ;
        RECT 20.535 83.135 20.865 83.465 ;
        RECT 20.550 67.145 20.850 83.135 ;
        RECT 20.535 66.815 20.865 67.145 ;
        RECT 38.030 66.465 38.330 92.655 ;
        RECT 88.615 89.935 88.945 90.265 ;
        RECT 88.630 67.145 88.930 89.935 ;
        RECT 88.615 66.815 88.945 67.145 ;
        RECT 38.015 66.135 38.345 66.465 ;
        RECT 38.030 58.305 38.330 66.135 ;
        RECT 34.335 57.975 34.665 58.305 ;
        RECT 38.015 57.975 38.345 58.305 ;
        RECT 34.350 34.505 34.650 57.975 ;
        RECT 88.630 52.865 88.930 66.815 ;
        RECT 88.615 52.535 88.945 52.865 ;
        RECT 88.630 34.505 88.930 52.535 ;
        RECT 34.335 34.175 34.665 34.505 ;
        RECT 88.615 34.175 88.945 34.505 ;
  END
END digital_top
END LIBRARY

