MACRO digital_top
  CLASS BLOCK ;
  FOREIGN digital_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 119.560 BY 130.280 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.520 10.640 26.520 117.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.520 10.640 56.520 117.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 84.520 10.640 86.520 117.200 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.520 10.640 11.520 117.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 39.520 10.640 41.520 117.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 69.520 10.640 71.520 117.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.520 10.640 101.520 117.200 ;
    END
  END VPWR
  PIN i_dem_dis
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 2.000 113.520 ;
    END
  END i_dem_dis
  PIN i_reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 2.000 48.240 ;
    END
  END i_reset
  PIN i_sys_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 2.000 80.880 ;
    END
  END i_sys_clk
  PIN o_cs_cell_hi[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 2.850 128.280 3.130 130.280 ;
    END
  END o_cs_cell_hi[0]
  PIN o_cs_cell_hi[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 8.830 128.280 9.110 130.280 ;
    END
  END o_cs_cell_hi[1]
  PIN o_cs_cell_hi[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 14.810 128.280 15.090 130.280 ;
    END
  END o_cs_cell_hi[2]
  PIN o_cs_cell_hi[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 20.790 128.280 21.070 130.280 ;
    END
  END o_cs_cell_hi[3]
  PIN o_cs_cell_hi[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 26.770 128.280 27.050 130.280 ;
    END
  END o_cs_cell_hi[4]
  PIN o_cs_cell_hi[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 32.750 128.280 33.030 130.280 ;
    END
  END o_cs_cell_hi[5]
  PIN o_cs_cell_hi[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 38.730 128.280 39.010 130.280 ;
    END
  END o_cs_cell_hi[6]
  PIN o_cs_cell_hi[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 44.710 128.280 44.990 130.280 ;
    END
  END o_cs_cell_hi[7]
  PIN o_cs_cell_hi[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 50.690 128.280 50.970 130.280 ;
    END
  END o_cs_cell_hi[8]
  PIN o_cs_cell_hi[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 56.670 128.280 56.950 130.280 ;
    END
  END o_cs_cell_hi[9]
  PIN o_cs_cell_lo[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 62.650 128.280 62.930 130.280 ;
    END
  END o_cs_cell_lo[0]
  PIN o_cs_cell_lo[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 68.630 128.280 68.910 130.280 ;
    END
  END o_cs_cell_lo[1]
  PIN o_cs_cell_lo[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 74.610 128.280 74.890 130.280 ;
    END
  END o_cs_cell_lo[2]
  PIN o_cs_cell_lo[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 80.590 128.280 80.870 130.280 ;
    END
  END o_cs_cell_lo[3]
  PIN o_cs_cell_lo[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 86.570 128.280 86.850 130.280 ;
    END
  END o_cs_cell_lo[4]
  PIN o_cs_cell_lo[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 92.550 128.280 92.830 130.280 ;
    END
  END o_cs_cell_lo[5]
  PIN o_cs_cell_lo[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 98.530 128.280 98.810 130.280 ;
    END
  END o_cs_cell_lo[6]
  PIN o_cs_cell_lo[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 104.510 128.280 104.790 130.280 ;
    END
  END o_cs_cell_lo[7]
  PIN o_cs_cell_lo[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 110.490 128.280 110.770 130.280 ;
    END
  END o_cs_cell_lo[8]
  PIN o_cs_cell_lo[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 116.470 128.280 116.750 130.280 ;
    END
  END o_cs_cell_lo[9]
  OBS
      LAYER nwell ;
        RECT 5.330 115.545 113.810 117.150 ;
      LAYER pwell ;
        RECT 5.525 114.345 6.895 115.155 ;
        RECT 6.905 114.345 8.275 115.125 ;
        RECT 8.285 114.345 13.795 115.155 ;
        RECT 13.805 114.345 17.475 115.155 ;
        RECT 18.415 114.430 18.845 115.215 ;
        RECT 18.865 114.345 24.375 115.155 ;
        RECT 24.385 114.345 29.895 115.155 ;
        RECT 29.905 114.345 31.275 115.155 ;
        RECT 31.295 114.430 31.725 115.215 ;
        RECT 31.745 115.025 32.665 115.255 ;
        RECT 35.495 115.025 36.425 115.245 ;
        RECT 31.745 114.345 40.935 115.025 ;
        RECT 40.945 114.345 43.695 115.155 ;
        RECT 44.175 114.430 44.605 115.215 ;
        RECT 44.625 114.345 50.135 115.155 ;
        RECT 51.075 114.345 52.425 115.255 ;
        RECT 52.915 114.345 54.265 115.255 ;
        RECT 54.285 114.345 57.035 115.155 ;
        RECT 57.055 114.430 57.485 115.215 ;
        RECT 57.505 114.345 63.015 115.155 ;
        RECT 63.025 114.345 68.535 115.155 ;
        RECT 68.545 114.345 69.915 115.155 ;
        RECT 69.935 114.430 70.365 115.215 ;
        RECT 70.385 114.345 75.895 115.155 ;
        RECT 75.905 114.345 81.415 115.155 ;
        RECT 81.425 114.345 82.795 115.155 ;
        RECT 82.815 114.430 83.245 115.215 ;
        RECT 83.265 114.345 84.635 115.155 ;
        RECT 84.655 114.345 86.005 115.255 ;
        RECT 86.025 114.345 89.695 115.155 ;
        RECT 90.635 114.345 91.985 115.255 ;
        RECT 92.005 114.345 95.675 115.155 ;
        RECT 95.695 114.430 96.125 115.215 ;
        RECT 97.075 114.345 98.425 115.255 ;
        RECT 103.875 115.025 104.805 115.245 ;
        RECT 107.635 115.025 108.555 115.255 ;
        RECT 99.365 114.345 108.555 115.025 ;
        RECT 108.575 114.430 109.005 115.215 ;
        RECT 109.025 114.345 111.775 115.155 ;
        RECT 112.245 114.345 113.615 115.155 ;
        RECT 5.665 114.135 5.835 114.345 ;
        RECT 7.055 114.325 7.225 114.345 ;
        RECT 7.045 114.155 7.225 114.325 ;
        RECT 8.425 114.155 8.595 114.345 ;
        RECT 9.800 114.185 9.920 114.295 ;
        RECT 13.945 114.155 14.115 114.345 ;
        RECT 17.635 114.190 17.795 114.300 ;
        RECT 7.045 114.135 7.215 114.155 ;
        RECT 19.005 114.135 19.175 114.345 ;
        RECT 19.465 114.135 19.635 114.325 ;
        RECT 21.305 114.135 21.475 114.325 ;
        RECT 24.525 114.155 24.695 114.345 ;
        RECT 30.045 114.155 30.215 114.345 ;
        RECT 30.515 114.180 30.675 114.290 ;
        RECT 31.885 114.135 32.055 114.325 ;
        RECT 37.415 114.180 37.575 114.290 ;
        RECT 38.325 114.135 38.495 114.325 ;
        RECT 40.625 114.155 40.795 114.345 ;
        RECT 41.085 114.155 41.255 114.345 ;
        RECT 43.840 114.185 43.960 114.295 ;
        RECT 44.765 114.155 44.935 114.345 ;
        RECT 47.520 114.185 47.640 114.295 ;
        RECT 47.985 114.135 48.155 114.325 ;
        RECT 50.295 114.190 50.455 114.300 ;
        RECT 51.205 114.155 51.375 114.345 ;
        RECT 52.580 114.185 52.700 114.295 ;
        RECT 53.045 114.155 53.215 114.345 ;
        RECT 54.425 114.155 54.595 114.345 ;
        RECT 57.645 114.135 57.815 114.345 ;
        RECT 61.335 114.180 61.495 114.290 ;
        RECT 62.245 114.135 62.415 114.325 ;
        RECT 63.165 114.155 63.335 114.345 ;
        RECT 68.685 114.155 68.855 114.345 ;
        RECT 70.525 114.155 70.695 114.345 ;
        RECT 71.445 114.135 71.615 114.325 ;
        RECT 76.045 114.155 76.215 114.345 ;
        RECT 81.565 114.135 81.735 114.345 ;
        RECT 82.035 114.180 82.195 114.290 ;
        RECT 83.405 114.135 83.575 114.345 ;
        RECT 84.785 114.155 84.955 114.345 ;
        RECT 86.165 114.155 86.335 114.345 ;
        RECT 89.855 114.190 90.015 114.300 ;
        RECT 90.765 114.155 90.935 114.345 ;
        RECT 92.145 114.155 92.315 114.345 ;
        RECT 92.605 114.135 92.775 114.325 ;
        RECT 96.295 114.190 96.455 114.300 ;
        RECT 97.205 114.155 97.375 114.345 ;
        RECT 98.595 114.190 98.755 114.300 ;
        RECT 99.505 114.155 99.675 114.345 ;
        RECT 102.725 114.135 102.895 114.325 ;
        RECT 104.105 114.135 104.275 114.325 ;
        RECT 104.565 114.135 104.735 114.325 ;
        RECT 106.400 114.185 106.520 114.295 ;
        RECT 106.865 114.135 107.035 114.325 ;
        RECT 108.240 114.185 108.360 114.295 ;
        RECT 109.165 114.135 109.335 114.345 ;
        RECT 111.920 114.185 112.040 114.295 ;
        RECT 113.305 114.135 113.475 114.345 ;
        RECT 5.525 113.325 6.895 114.135 ;
        RECT 6.905 113.325 9.655 114.135 ;
        RECT 10.125 113.455 19.315 114.135 ;
        RECT 10.125 113.225 11.045 113.455 ;
        RECT 13.875 113.235 14.805 113.455 ;
        RECT 19.325 113.325 21.155 114.135 ;
        RECT 21.165 113.455 30.355 114.135 ;
        RECT 25.675 113.235 26.605 113.455 ;
        RECT 29.435 113.225 30.355 113.455 ;
        RECT 31.295 113.265 31.725 114.050 ;
        RECT 31.745 113.325 37.255 114.135 ;
        RECT 38.185 113.455 47.375 114.135 ;
        RECT 47.845 113.455 57.035 114.135 ;
        RECT 42.695 113.235 43.625 113.455 ;
        RECT 46.455 113.225 47.375 113.455 ;
        RECT 52.355 113.235 53.285 113.455 ;
        RECT 56.115 113.225 57.035 113.455 ;
        RECT 57.055 113.265 57.485 114.050 ;
        RECT 57.505 113.325 61.175 114.135 ;
        RECT 62.105 113.455 71.295 114.135 ;
        RECT 71.305 113.455 80.495 114.135 ;
        RECT 66.615 113.235 67.545 113.455 ;
        RECT 70.375 113.225 71.295 113.455 ;
        RECT 75.815 113.235 76.745 113.455 ;
        RECT 79.575 113.225 80.495 113.455 ;
        RECT 80.515 113.225 81.865 114.135 ;
        RECT 82.815 113.265 83.245 114.050 ;
        RECT 83.265 113.455 92.455 114.135 ;
        RECT 92.465 113.455 101.655 114.135 ;
        RECT 87.775 113.235 88.705 113.455 ;
        RECT 91.535 113.225 92.455 113.455 ;
        RECT 96.975 113.235 97.905 113.455 ;
        RECT 100.735 113.225 101.655 113.455 ;
        RECT 101.665 113.355 103.035 114.135 ;
        RECT 103.055 113.225 104.405 114.135 ;
        RECT 104.425 113.325 106.255 114.135 ;
        RECT 106.735 113.225 108.085 114.135 ;
        RECT 108.575 113.265 109.005 114.050 ;
        RECT 109.025 113.325 111.775 114.135 ;
        RECT 112.245 113.325 113.615 114.135 ;
      LAYER nwell ;
        RECT 5.330 110.105 113.810 112.935 ;
      LAYER pwell ;
        RECT 5.525 108.905 6.895 109.715 ;
        RECT 6.905 108.905 8.275 109.715 ;
        RECT 8.285 109.585 9.205 109.815 ;
        RECT 12.035 109.585 12.965 109.805 ;
        RECT 8.285 108.905 17.475 109.585 ;
        RECT 18.415 108.990 18.845 109.775 ;
        RECT 19.785 109.585 20.705 109.815 ;
        RECT 23.535 109.585 24.465 109.805 ;
        RECT 19.785 108.905 28.975 109.585 ;
        RECT 28.995 108.905 30.345 109.815 ;
        RECT 30.365 108.905 31.735 109.715 ;
        RECT 31.745 108.905 33.115 109.685 ;
        RECT 33.135 108.905 34.485 109.815 ;
        RECT 39.015 109.585 39.945 109.805 ;
        RECT 42.775 109.585 43.695 109.815 ;
        RECT 34.505 108.905 43.695 109.585 ;
        RECT 44.175 108.990 44.605 109.775 ;
        RECT 45.545 108.905 46.915 109.685 ;
        RECT 51.435 109.585 52.365 109.805 ;
        RECT 55.195 109.585 56.115 109.815 ;
        RECT 46.925 108.905 56.115 109.585 ;
        RECT 56.135 108.905 57.485 109.815 ;
        RECT 57.505 108.905 58.875 109.715 ;
        RECT 63.395 109.585 64.325 109.805 ;
        RECT 67.155 109.585 68.075 109.815 ;
        RECT 58.885 108.905 68.075 109.585 ;
        RECT 68.085 108.905 69.455 109.685 ;
        RECT 69.935 108.990 70.365 109.775 ;
        RECT 70.395 108.905 71.745 109.815 ;
        RECT 72.685 108.905 74.055 109.685 ;
        RECT 78.575 109.585 79.505 109.805 ;
        RECT 82.335 109.585 83.255 109.815 ;
        RECT 74.065 108.905 83.255 109.585 ;
        RECT 83.265 108.905 84.635 109.685 ;
        RECT 90.075 109.585 91.005 109.805 ;
        RECT 93.835 109.585 94.755 109.815 ;
        RECT 85.565 108.905 94.755 109.585 ;
        RECT 95.695 108.990 96.125 109.775 ;
        RECT 96.145 108.905 97.515 109.685 ;
        RECT 102.035 109.585 102.965 109.805 ;
        RECT 105.795 109.585 106.715 109.815 ;
        RECT 97.525 108.905 106.715 109.585 ;
        RECT 106.725 108.905 112.235 109.715 ;
        RECT 112.245 108.905 113.615 109.715 ;
        RECT 5.665 108.695 5.835 108.905 ;
        RECT 7.045 108.695 7.215 108.905 ;
        RECT 17.165 108.695 17.335 108.905 ;
        RECT 17.635 108.750 17.795 108.860 ;
        RECT 18.545 108.695 18.715 108.885 ;
        RECT 19.015 108.740 19.175 108.860 ;
        RECT 20.845 108.695 21.015 108.885 ;
        RECT 21.305 108.695 21.475 108.885 ;
        RECT 23.605 108.695 23.775 108.885 ;
        RECT 24.060 108.745 24.180 108.855 ;
        RECT 25.445 108.695 25.615 108.885 ;
        RECT 26.825 108.695 26.995 108.885 ;
        RECT 27.285 108.695 27.455 108.885 ;
        RECT 28.665 108.715 28.835 108.905 ;
        RECT 30.045 108.715 30.215 108.905 ;
        RECT 30.505 108.715 30.675 108.905 ;
        RECT 30.960 108.745 31.080 108.855 ;
        RECT 31.885 108.695 32.055 108.905 ;
        RECT 33.265 108.715 33.435 108.905 ;
        RECT 34.645 108.715 34.815 108.905 ;
        RECT 37.405 108.695 37.575 108.885 ;
        RECT 40.165 108.695 40.335 108.885 ;
        RECT 41.545 108.695 41.715 108.885 ;
        RECT 42.000 108.745 42.120 108.855 ;
        RECT 43.385 108.695 43.555 108.885 ;
        RECT 43.840 108.745 43.960 108.855 ;
        RECT 44.765 108.695 44.935 108.885 ;
        RECT 45.225 108.695 45.395 108.885 ;
        RECT 45.685 108.715 45.855 108.905 ;
        RECT 47.065 108.715 47.235 108.905 ;
        RECT 48.915 108.740 49.075 108.850 ;
        RECT 52.120 108.695 52.290 108.885 ;
        RECT 53.505 108.695 53.675 108.885 ;
        RECT 53.965 108.695 54.135 108.885 ;
        RECT 56.265 108.715 56.435 108.905 ;
        RECT 56.720 108.745 56.840 108.855 ;
        RECT 57.645 108.695 57.815 108.905 ;
        RECT 59.025 108.715 59.195 108.905 ;
        RECT 61.325 108.695 61.495 108.885 ;
        RECT 63.625 108.695 63.795 108.885 ;
        RECT 64.085 108.695 64.255 108.885 ;
        RECT 66.845 108.695 67.015 108.885 ;
        RECT 67.305 108.695 67.475 108.885 ;
        RECT 69.145 108.715 69.315 108.905 ;
        RECT 69.600 108.745 69.720 108.855 ;
        RECT 70.980 108.695 71.150 108.885 ;
        RECT 71.445 108.695 71.615 108.905 ;
        RECT 71.915 108.750 72.075 108.860 ;
        RECT 73.285 108.695 73.455 108.885 ;
        RECT 73.745 108.715 73.915 108.905 ;
        RECT 74.205 108.715 74.375 108.905 ;
        RECT 74.665 108.695 74.835 108.885 ;
        RECT 79.265 108.695 79.435 108.885 ;
        RECT 79.725 108.695 79.895 108.885 ;
        RECT 82.480 108.745 82.600 108.855 ;
        RECT 83.405 108.695 83.575 108.905 ;
        RECT 84.795 108.750 84.955 108.860 ;
        RECT 85.705 108.715 85.875 108.905 ;
        RECT 88.005 108.695 88.175 108.885 ;
        RECT 88.465 108.695 88.635 108.885 ;
        RECT 93.985 108.695 94.155 108.885 ;
        RECT 94.915 108.750 95.075 108.860 ;
        RECT 95.820 108.745 95.940 108.855 ;
        RECT 96.285 108.695 96.455 108.885 ;
        RECT 97.205 108.715 97.375 108.905 ;
        RECT 97.665 108.715 97.835 108.905 ;
        RECT 98.585 108.695 98.755 108.885 ;
        RECT 106.865 108.715 107.035 108.905 ;
        RECT 107.795 108.740 107.955 108.850 ;
        RECT 109.165 108.695 109.335 108.885 ;
        RECT 111.920 108.745 112.040 108.855 ;
        RECT 113.305 108.695 113.475 108.905 ;
        RECT 5.525 107.885 6.895 108.695 ;
        RECT 6.905 108.015 16.095 108.695 ;
        RECT 11.415 107.795 12.345 108.015 ;
        RECT 15.175 107.785 16.095 108.015 ;
        RECT 16.115 107.785 17.465 108.695 ;
        RECT 17.495 107.785 18.845 108.695 ;
        RECT 19.785 107.915 21.155 108.695 ;
        RECT 21.165 107.885 22.535 108.695 ;
        RECT 22.545 107.915 23.915 108.695 ;
        RECT 24.385 107.915 25.755 108.695 ;
        RECT 25.775 107.785 27.125 108.695 ;
        RECT 27.145 107.885 30.815 108.695 ;
        RECT 31.295 107.825 31.725 108.610 ;
        RECT 31.745 107.885 37.255 108.695 ;
        RECT 37.265 107.885 39.095 108.695 ;
        RECT 39.105 107.915 40.475 108.695 ;
        RECT 40.495 107.785 41.845 108.695 ;
        RECT 42.325 107.915 43.695 108.695 ;
        RECT 43.715 107.785 45.065 108.695 ;
        RECT 45.085 107.885 48.755 108.695 ;
        RECT 49.825 107.785 52.435 108.695 ;
        RECT 52.445 107.915 53.815 108.695 ;
        RECT 53.825 107.885 56.575 108.695 ;
        RECT 57.055 107.825 57.485 108.610 ;
        RECT 57.505 107.885 61.175 108.695 ;
        RECT 61.185 107.885 62.555 108.695 ;
        RECT 62.565 107.915 63.935 108.695 ;
        RECT 63.945 107.885 65.775 108.695 ;
        RECT 65.795 107.785 67.145 108.695 ;
        RECT 67.165 107.885 68.535 108.695 ;
        RECT 68.685 107.785 71.295 108.695 ;
        RECT 71.305 107.885 73.135 108.695 ;
        RECT 73.155 107.785 74.505 108.695 ;
        RECT 74.525 107.885 78.195 108.695 ;
        RECT 78.205 107.915 79.575 108.695 ;
        RECT 79.585 107.885 82.335 108.695 ;
        RECT 82.815 107.825 83.245 108.610 ;
        RECT 83.265 107.885 86.935 108.695 ;
        RECT 86.945 107.915 88.315 108.695 ;
        RECT 88.325 107.885 93.835 108.695 ;
        RECT 93.845 107.885 95.675 108.695 ;
        RECT 96.145 107.915 97.515 108.695 ;
        RECT 98.445 108.015 107.635 108.695 ;
        RECT 102.955 107.795 103.885 108.015 ;
        RECT 106.715 107.785 107.635 108.015 ;
        RECT 108.575 107.825 109.005 108.610 ;
        RECT 109.025 107.885 111.775 108.695 ;
        RECT 112.245 107.885 113.615 108.695 ;
      LAYER nwell ;
        RECT 5.330 104.665 113.810 107.495 ;
      LAYER pwell ;
        RECT 5.525 103.465 6.895 104.275 ;
        RECT 6.905 103.465 9.655 104.275 ;
        RECT 9.665 103.465 11.035 104.245 ;
        RECT 11.965 103.465 13.335 104.245 ;
        RECT 14.275 103.465 15.625 104.375 ;
        RECT 15.645 103.465 18.395 104.275 ;
        RECT 18.415 103.550 18.845 104.335 ;
        RECT 18.865 103.465 24.375 104.275 ;
        RECT 24.385 103.465 29.895 104.275 ;
        RECT 29.905 103.465 35.415 104.275 ;
        RECT 35.435 103.465 36.785 104.375 ;
        RECT 36.805 103.465 42.315 104.275 ;
        RECT 42.325 103.465 44.155 104.275 ;
        RECT 44.175 103.550 44.605 104.335 ;
        RECT 44.625 103.465 45.995 104.275 ;
        RECT 46.005 104.145 46.935 104.375 ;
        RECT 46.005 103.465 49.905 104.145 ;
        RECT 50.145 103.465 55.655 104.275 ;
        RECT 55.665 103.465 61.175 104.275 ;
        RECT 61.185 103.465 66.695 104.275 ;
        RECT 66.705 103.465 69.455 104.275 ;
        RECT 69.935 103.550 70.365 104.335 ;
        RECT 70.385 104.145 71.315 104.375 ;
        RECT 70.385 103.465 74.285 104.145 ;
        RECT 74.535 103.465 75.885 104.375 ;
        RECT 75.905 103.465 81.415 104.275 ;
        RECT 81.425 103.465 86.935 104.275 ;
        RECT 86.945 103.465 92.455 104.275 ;
        RECT 92.465 103.465 95.215 104.275 ;
        RECT 95.695 103.550 96.125 104.335 ;
        RECT 96.155 103.465 97.505 104.375 ;
        RECT 97.525 103.465 98.895 104.245 ;
        RECT 98.905 103.465 102.575 104.275 ;
        RECT 102.585 103.465 103.955 104.275 ;
        RECT 103.975 103.465 105.325 104.375 ;
        RECT 105.345 103.465 110.855 104.275 ;
        RECT 110.865 103.465 112.235 104.275 ;
        RECT 112.245 103.465 113.615 104.275 ;
        RECT 5.665 103.255 5.835 103.465 ;
        RECT 7.045 103.255 7.215 103.465 ;
        RECT 10.725 103.275 10.895 103.465 ;
        RECT 11.195 103.310 11.355 103.420 ;
        RECT 12.565 103.255 12.735 103.445 ;
        RECT 13.025 103.275 13.195 103.465 ;
        RECT 13.495 103.310 13.655 103.420 ;
        RECT 15.325 103.275 15.495 103.465 ;
        RECT 15.785 103.275 15.955 103.465 ;
        RECT 16.245 103.255 16.415 103.445 ;
        RECT 19.005 103.275 19.175 103.465 ;
        RECT 24.525 103.275 24.695 103.465 ;
        RECT 25.905 103.255 26.075 103.445 ;
        RECT 27.745 103.255 27.915 103.445 ;
        RECT 29.125 103.255 29.295 103.445 ;
        RECT 30.045 103.275 30.215 103.465 ;
        RECT 30.960 103.305 31.080 103.415 ;
        RECT 36.485 103.275 36.655 103.465 ;
        RECT 36.945 103.275 37.115 103.465 ;
        RECT 41.085 103.255 41.255 103.445 ;
        RECT 42.465 103.255 42.635 103.465 ;
        RECT 42.935 103.300 43.095 103.410 ;
        RECT 43.845 103.255 44.015 103.445 ;
        RECT 44.765 103.275 44.935 103.465 ;
        RECT 46.420 103.275 46.590 103.465 ;
        RECT 50.285 103.275 50.455 103.465 ;
        RECT 53.505 103.255 53.675 103.445 ;
        RECT 54.885 103.255 55.055 103.445 ;
        RECT 55.805 103.275 55.975 103.465 ;
        RECT 56.720 103.305 56.840 103.415 ;
        RECT 57.645 103.255 57.815 103.445 ;
        RECT 60.405 103.255 60.575 103.445 ;
        RECT 61.325 103.275 61.495 103.465 ;
        RECT 62.060 103.255 62.230 103.445 ;
        RECT 65.925 103.255 66.095 103.445 ;
        RECT 66.845 103.275 67.015 103.465 ;
        RECT 69.600 103.305 69.720 103.415 ;
        RECT 70.800 103.275 70.970 103.465 ;
        RECT 75.585 103.445 75.755 103.465 ;
        RECT 75.585 103.275 75.760 103.445 ;
        RECT 76.045 103.275 76.215 103.465 ;
        RECT 75.590 103.255 75.760 103.275 ;
        RECT 78.345 103.255 78.515 103.445 ;
        RECT 79.725 103.255 79.895 103.445 ;
        RECT 81.100 103.305 81.220 103.415 ;
        RECT 81.565 103.255 81.735 103.465 ;
        RECT 83.405 103.255 83.575 103.445 ;
        RECT 84.785 103.255 84.955 103.445 ;
        RECT 86.165 103.255 86.335 103.445 ;
        RECT 87.085 103.275 87.255 103.465 ;
        RECT 92.605 103.275 92.775 103.465 ;
        RECT 95.360 103.305 95.480 103.415 ;
        RECT 95.820 103.305 95.940 103.415 ;
        RECT 96.285 103.255 96.455 103.445 ;
        RECT 97.205 103.275 97.375 103.465 ;
        RECT 97.665 103.275 97.835 103.465 ;
        RECT 99.045 103.275 99.215 103.465 ;
        RECT 102.725 103.275 102.895 103.465 ;
        RECT 105.025 103.275 105.195 103.465 ;
        RECT 105.485 103.275 105.655 103.465 ;
        RECT 106.405 103.255 106.575 103.445 ;
        RECT 106.865 103.255 107.035 103.445 ;
        RECT 108.240 103.305 108.360 103.415 ;
        RECT 109.165 103.255 109.335 103.445 ;
        RECT 111.005 103.275 111.175 103.465 ;
        RECT 111.920 103.305 112.040 103.415 ;
        RECT 113.305 103.255 113.475 103.465 ;
        RECT 5.525 102.445 6.895 103.255 ;
        RECT 6.905 102.445 12.415 103.255 ;
        RECT 12.425 102.445 16.095 103.255 ;
        RECT 16.105 102.575 25.385 103.255 ;
        RECT 17.465 102.355 18.385 102.575 ;
        RECT 23.050 102.455 25.385 102.575 ;
        RECT 24.465 102.345 25.385 102.455 ;
        RECT 25.765 102.445 27.595 103.255 ;
        RECT 27.605 102.475 28.975 103.255 ;
        RECT 28.985 102.445 30.815 103.255 ;
        RECT 31.295 102.385 31.725 103.170 ;
        RECT 32.115 102.575 41.395 103.255 ;
        RECT 32.115 102.455 34.450 102.575 ;
        RECT 32.115 102.345 33.035 102.455 ;
        RECT 39.115 102.355 40.035 102.575 ;
        RECT 41.415 102.345 42.765 103.255 ;
        RECT 43.705 102.575 52.985 103.255 ;
        RECT 45.065 102.355 45.985 102.575 ;
        RECT 50.650 102.455 52.985 102.575 ;
        RECT 53.365 102.475 54.735 103.255 ;
        RECT 52.065 102.345 52.985 102.455 ;
        RECT 54.745 102.445 56.575 103.255 ;
        RECT 57.055 102.385 57.485 103.170 ;
        RECT 57.505 102.445 60.255 103.255 ;
        RECT 60.275 102.345 61.625 103.255 ;
        RECT 61.645 102.575 65.545 103.255 ;
        RECT 65.785 102.575 75.065 103.255 ;
        RECT 61.645 102.345 62.575 102.575 ;
        RECT 67.145 102.355 68.065 102.575 ;
        RECT 72.730 102.455 75.065 102.575 ;
        RECT 74.145 102.345 75.065 102.455 ;
        RECT 75.445 102.345 78.055 103.255 ;
        RECT 78.205 102.445 79.575 103.255 ;
        RECT 79.585 102.475 80.955 103.255 ;
        RECT 81.435 102.345 82.785 103.255 ;
        RECT 82.815 102.385 83.245 103.170 ;
        RECT 83.265 102.445 84.635 103.255 ;
        RECT 84.645 102.475 86.015 103.255 ;
        RECT 86.025 102.575 95.305 103.255 ;
        RECT 96.145 102.575 105.250 103.255 ;
        RECT 87.385 102.355 88.305 102.575 ;
        RECT 92.970 102.455 95.305 102.575 ;
        RECT 105.345 102.475 106.715 103.255 ;
        RECT 94.385 102.345 95.305 102.455 ;
        RECT 106.735 102.345 108.085 103.255 ;
        RECT 108.575 102.385 109.005 103.170 ;
        RECT 109.025 102.445 111.775 103.255 ;
        RECT 112.245 102.445 113.615 103.255 ;
      LAYER nwell ;
        RECT 5.330 99.225 113.810 102.055 ;
      LAYER pwell ;
        RECT 5.525 98.025 6.895 98.835 ;
        RECT 9.185 98.705 10.105 98.925 ;
        RECT 16.185 98.825 17.105 98.935 ;
        RECT 14.770 98.705 17.105 98.825 ;
        RECT 7.825 98.025 17.105 98.705 ;
        RECT 18.415 98.110 18.845 98.895 ;
        RECT 18.865 98.705 19.795 98.935 ;
        RECT 18.865 98.025 22.765 98.705 ;
        RECT 23.015 98.025 24.365 98.935 ;
        RECT 25.305 98.025 26.675 98.805 ;
        RECT 26.685 98.705 27.615 98.935 ;
        RECT 26.685 98.025 30.585 98.705 ;
        RECT 31.285 98.025 32.655 98.805 ;
        RECT 34.025 98.705 34.945 98.925 ;
        RECT 41.025 98.825 41.945 98.935 ;
        RECT 39.610 98.705 41.945 98.825 ;
        RECT 32.665 98.025 41.945 98.705 ;
        RECT 42.325 98.025 43.695 98.805 ;
        RECT 44.175 98.110 44.605 98.895 ;
        RECT 47.295 98.825 48.215 98.935 ;
        RECT 45.545 98.025 46.915 98.805 ;
        RECT 47.295 98.705 49.630 98.825 ;
        RECT 54.295 98.705 55.215 98.925 ;
        RECT 57.945 98.705 58.865 98.925 ;
        RECT 64.945 98.825 65.865 98.935 ;
        RECT 63.530 98.705 65.865 98.825 ;
        RECT 47.295 98.025 56.575 98.705 ;
        RECT 56.585 98.025 65.865 98.705 ;
        RECT 66.245 98.025 68.075 98.835 ;
        RECT 68.085 98.025 69.455 98.805 ;
        RECT 69.935 98.110 70.365 98.895 ;
        RECT 70.385 98.025 72.215 98.835 ;
        RECT 72.685 98.025 83.695 98.935 ;
        RECT 85.085 98.705 86.005 98.925 ;
        RECT 92.085 98.825 93.005 98.935 ;
        RECT 90.670 98.705 93.005 98.825 ;
        RECT 83.725 98.025 93.005 98.705 ;
        RECT 93.845 98.025 95.215 98.805 ;
        RECT 95.695 98.110 96.125 98.895 ;
        RECT 96.145 98.705 97.075 98.935 ;
        RECT 103.945 98.705 104.865 98.925 ;
        RECT 110.945 98.825 111.865 98.935 ;
        RECT 109.530 98.705 111.865 98.825 ;
        RECT 96.145 98.025 100.045 98.705 ;
        RECT 100.700 98.025 101.655 98.705 ;
        RECT 102.585 98.025 111.865 98.705 ;
        RECT 112.245 98.025 113.615 98.835 ;
        RECT 5.665 97.815 5.835 98.025 ;
        RECT 7.045 97.815 7.215 98.005 ;
        RECT 7.965 97.835 8.135 98.025 ;
        RECT 10.720 97.865 10.840 97.975 ;
        RECT 12.105 97.815 12.275 98.005 ;
        RECT 12.560 97.865 12.680 97.975 ;
        RECT 13.945 97.815 14.115 98.005 ;
        RECT 14.405 97.815 14.575 98.005 ;
        RECT 17.160 97.865 17.280 97.975 ;
        RECT 17.635 97.870 17.795 97.980 ;
        RECT 18.545 97.815 18.715 98.005 ;
        RECT 19.005 97.835 19.175 98.005 ;
        RECT 19.280 97.835 19.450 98.025 ;
        RECT 20.385 97.815 20.555 98.005 ;
        RECT 24.065 97.835 24.235 98.025 ;
        RECT 24.535 97.870 24.695 97.980 ;
        RECT 26.365 97.835 26.535 98.025 ;
        RECT 27.100 97.835 27.270 98.025 ;
        RECT 30.505 97.815 30.675 98.005 ;
        RECT 30.960 97.865 31.080 97.975 ;
        RECT 31.425 97.835 31.595 98.025 ;
        RECT 31.885 97.815 32.055 98.005 ;
        RECT 32.805 97.835 32.975 98.025 ;
        RECT 33.540 97.815 33.710 98.005 ;
        RECT 42.465 97.835 42.635 98.025 ;
        RECT 43.840 97.865 43.960 97.975 ;
        RECT 44.775 97.870 44.935 97.980 ;
        RECT 46.605 97.815 46.775 98.025 ;
        RECT 47.065 97.815 47.235 98.005 ;
        RECT 56.265 97.835 56.435 98.025 ;
        RECT 56.725 97.835 56.895 98.025 ;
        RECT 58.565 97.815 58.735 98.005 ;
        RECT 59.035 97.860 59.195 97.970 ;
        RECT 60.865 97.815 61.035 98.005 ;
        RECT 61.325 97.815 61.495 98.005 ;
        RECT 65.000 97.865 65.120 97.975 ;
        RECT 65.465 97.815 65.635 98.005 ;
        RECT 66.385 97.835 66.555 98.025 ;
        RECT 69.145 97.835 69.315 98.025 ;
        RECT 69.600 97.865 69.720 97.975 ;
        RECT 70.525 97.835 70.695 98.025 ;
        RECT 72.360 97.865 72.480 97.975 ;
        RECT 72.830 97.835 73.000 98.025 ;
        RECT 78.340 97.815 78.510 98.005 ;
        RECT 78.805 97.835 78.975 98.005 ;
        RECT 78.825 97.815 78.975 97.835 ;
        RECT 81.105 97.815 81.275 98.005 ;
        RECT 83.680 97.815 83.850 98.005 ;
        RECT 83.865 97.835 84.035 98.025 ;
        RECT 87.820 97.815 87.990 98.005 ;
        RECT 91.685 97.815 91.855 98.005 ;
        RECT 93.520 97.865 93.640 97.975 ;
        RECT 94.905 97.835 95.075 98.025 ;
        RECT 95.360 97.865 95.480 97.975 ;
        RECT 96.560 97.835 96.730 98.025 ;
        RECT 100.425 97.835 100.595 98.005 ;
        RECT 101.815 97.870 101.975 97.980 ;
        RECT 102.265 97.815 102.435 98.005 ;
        RECT 102.725 97.835 102.895 98.025 ;
        RECT 107.050 97.815 107.220 98.005 ;
        RECT 107.795 97.860 107.955 97.970 ;
        RECT 109.165 97.815 109.335 98.005 ;
        RECT 111.920 97.865 112.040 97.975 ;
        RECT 113.305 97.815 113.475 98.025 ;
        RECT 5.525 97.005 6.895 97.815 ;
        RECT 6.905 97.005 10.575 97.815 ;
        RECT 11.045 97.035 12.415 97.815 ;
        RECT 12.895 96.905 14.245 97.815 ;
        RECT 14.265 97.005 17.015 97.815 ;
        RECT 17.485 97.035 18.855 97.815 ;
        RECT 19.280 97.135 20.235 97.815 ;
        RECT 20.245 97.135 29.350 97.815 ;
        RECT 29.455 96.905 30.805 97.815 ;
        RECT 31.295 96.945 31.725 97.730 ;
        RECT 31.745 97.005 33.115 97.815 ;
        RECT 33.125 97.135 37.025 97.815 ;
        RECT 37.635 97.135 46.915 97.815 ;
        RECT 46.925 97.135 56.030 97.815 ;
        RECT 33.125 96.905 34.055 97.135 ;
        RECT 37.635 97.015 39.970 97.135 ;
        RECT 37.635 96.905 38.555 97.015 ;
        RECT 44.635 96.915 45.555 97.135 ;
        RECT 57.055 96.945 57.485 97.730 ;
        RECT 57.515 96.905 58.865 97.815 ;
        RECT 59.805 97.035 61.175 97.815 ;
        RECT 61.185 97.005 64.855 97.815 ;
        RECT 65.325 97.135 74.605 97.815 ;
        RECT 66.685 96.915 67.605 97.135 ;
        RECT 72.270 97.015 74.605 97.135 ;
        RECT 73.685 96.905 74.605 97.015 ;
        RECT 75.180 96.905 78.655 97.815 ;
        RECT 78.825 96.995 80.755 97.815 ;
        RECT 80.965 97.005 82.795 97.815 ;
        RECT 79.805 96.905 80.755 96.995 ;
        RECT 82.815 96.945 83.245 97.730 ;
        RECT 83.265 97.135 87.165 97.815 ;
        RECT 87.405 97.135 91.305 97.815 ;
        RECT 91.545 97.135 100.825 97.815 ;
        RECT 83.265 96.905 84.195 97.135 ;
        RECT 87.405 96.905 88.335 97.135 ;
        RECT 92.905 96.915 93.825 97.135 ;
        RECT 98.490 97.015 100.825 97.135 ;
        RECT 99.905 96.905 100.825 97.015 ;
        RECT 101.215 96.905 102.565 97.815 ;
        RECT 103.735 97.135 107.635 97.815 ;
        RECT 106.705 96.905 107.635 97.135 ;
        RECT 108.575 96.945 109.005 97.730 ;
        RECT 109.025 97.005 111.775 97.815 ;
        RECT 112.245 97.005 113.615 97.815 ;
      LAYER nwell ;
        RECT 5.330 93.785 113.810 96.615 ;
      LAYER pwell ;
        RECT 5.525 92.585 6.895 93.395 ;
        RECT 6.905 92.585 10.575 93.395 ;
        RECT 11.045 92.585 12.415 93.365 ;
        RECT 12.895 92.585 14.245 93.495 ;
        RECT 14.265 93.265 15.195 93.495 ;
        RECT 14.265 92.585 18.165 93.265 ;
        RECT 18.415 92.670 18.845 93.455 ;
        RECT 18.865 92.585 21.615 93.395 ;
        RECT 23.445 93.265 24.365 93.485 ;
        RECT 30.445 93.385 31.365 93.495 ;
        RECT 29.030 93.265 31.365 93.385 ;
        RECT 22.085 92.585 31.365 93.265 ;
        RECT 31.745 92.585 37.255 93.395 ;
        RECT 37.265 92.585 40.935 93.395 ;
        RECT 41.415 92.585 42.765 93.495 ;
        RECT 42.785 92.585 44.155 93.395 ;
        RECT 44.175 92.670 44.605 93.455 ;
        RECT 44.625 93.265 45.555 93.495 ;
        RECT 44.625 92.585 48.525 93.265 ;
        RECT 48.775 92.585 50.125 93.495 ;
        RECT 53.345 93.265 54.275 93.495 ;
        RECT 50.375 92.585 54.275 93.265 ;
        RECT 54.485 93.405 55.435 93.495 ;
        RECT 54.485 92.585 56.415 93.405 ;
        RECT 56.585 92.585 62.095 93.395 ;
        RECT 62.105 92.585 67.615 93.395 ;
        RECT 67.625 92.585 68.995 93.365 ;
        RECT 69.935 92.670 70.365 93.455 ;
        RECT 82.085 93.405 83.035 93.495 ;
        RECT 84.385 93.405 85.335 93.495 ;
        RECT 86.685 93.405 87.635 93.495 ;
        RECT 70.385 92.585 72.215 93.395 ;
        RECT 72.685 92.585 81.790 93.265 ;
        RECT 82.085 92.585 84.015 93.405 ;
        RECT 84.385 92.585 86.315 93.405 ;
        RECT 86.685 92.585 88.615 93.405 ;
        RECT 88.785 92.585 90.155 93.395 ;
        RECT 90.165 92.585 91.535 93.365 ;
        RECT 91.545 92.585 95.215 93.395 ;
        RECT 95.695 92.670 96.125 93.455 ;
        RECT 96.145 92.585 98.895 93.395 ;
        RECT 99.365 92.585 100.735 93.365 ;
        RECT 102.105 93.265 103.025 93.485 ;
        RECT 109.105 93.385 110.025 93.495 ;
        RECT 107.690 93.265 110.025 93.385 ;
        RECT 100.745 92.585 110.025 93.265 ;
        RECT 110.415 92.585 111.765 93.495 ;
        RECT 112.245 92.585 113.615 93.395 ;
        RECT 5.665 92.375 5.835 92.585 ;
        RECT 7.045 92.395 7.215 92.585 ;
        RECT 7.965 92.375 8.135 92.565 ;
        RECT 10.720 92.425 10.840 92.535 ;
        RECT 12.105 92.395 12.275 92.585 ;
        RECT 12.560 92.425 12.680 92.535 ;
        RECT 13.945 92.395 14.115 92.585 ;
        RECT 14.680 92.395 14.850 92.585 ;
        RECT 17.900 92.375 18.070 92.565 ;
        RECT 19.005 92.395 19.175 92.585 ;
        RECT 21.765 92.535 21.935 92.565 ;
        RECT 21.760 92.425 21.935 92.535 ;
        RECT 21.765 92.375 21.935 92.425 ;
        RECT 22.225 92.395 22.395 92.585 ;
        RECT 24.525 92.395 24.695 92.565 ;
        RECT 26.820 92.425 26.940 92.535 ;
        RECT 24.545 92.375 24.695 92.395 ;
        RECT 27.560 92.375 27.730 92.565 ;
        RECT 31.885 92.395 32.055 92.585 ;
        RECT 33.725 92.395 33.895 92.565 ;
        RECT 33.725 92.375 33.875 92.395 ;
        RECT 34.185 92.375 34.355 92.565 ;
        RECT 37.405 92.395 37.575 92.585 ;
        RECT 39.705 92.375 39.875 92.565 ;
        RECT 41.080 92.425 41.200 92.535 ;
        RECT 42.465 92.395 42.635 92.585 ;
        RECT 42.925 92.395 43.095 92.585 ;
        RECT 45.040 92.395 45.210 92.585 ;
        RECT 45.225 92.375 45.395 92.565 ;
        RECT 47.980 92.425 48.100 92.535 ;
        RECT 48.445 92.395 48.615 92.565 ;
        RECT 49.825 92.395 49.995 92.585 ;
        RECT 50.745 92.395 50.915 92.565 ;
        RECT 53.045 92.395 53.215 92.565 ;
        RECT 53.690 92.395 53.860 92.585 ;
        RECT 56.265 92.565 56.415 92.585 ;
        RECT 48.465 92.375 48.615 92.395 ;
        RECT 50.765 92.375 50.915 92.395 ;
        RECT 53.065 92.375 53.215 92.395 ;
        RECT 55.345 92.375 55.515 92.565 ;
        RECT 56.265 92.395 56.435 92.565 ;
        RECT 56.725 92.395 56.895 92.585 ;
        RECT 59.945 92.375 60.115 92.565 ;
        RECT 62.245 92.395 62.415 92.585 ;
        RECT 62.245 92.375 62.395 92.395 ;
        RECT 63.625 92.375 63.795 92.565 ;
        RECT 64.085 92.375 64.255 92.565 ;
        RECT 67.765 92.375 67.935 92.565 ;
        RECT 68.685 92.395 68.855 92.585 ;
        RECT 69.145 92.375 69.315 92.565 ;
        RECT 70.525 92.395 70.695 92.585 ;
        RECT 70.800 92.375 70.970 92.565 ;
        RECT 72.360 92.425 72.480 92.535 ;
        RECT 72.825 92.395 72.995 92.585 ;
        RECT 83.865 92.565 84.015 92.585 ;
        RECT 86.165 92.565 86.315 92.585 ;
        RECT 88.465 92.565 88.615 92.585 ;
        RECT 74.675 92.420 74.835 92.530 ;
        RECT 78.800 92.375 78.970 92.565 ;
        RECT 5.525 91.565 6.895 92.375 ;
        RECT 7.825 91.695 17.105 92.375 ;
        RECT 9.185 91.475 10.105 91.695 ;
        RECT 14.770 91.575 17.105 91.695 ;
        RECT 16.185 91.465 17.105 91.575 ;
        RECT 17.485 91.695 21.385 92.375 ;
        RECT 17.485 91.465 18.415 91.695 ;
        RECT 21.625 91.565 24.375 92.375 ;
        RECT 24.545 91.555 26.475 92.375 ;
        RECT 25.525 91.465 26.475 91.555 ;
        RECT 27.145 91.695 31.045 92.375 ;
        RECT 27.145 91.465 28.075 91.695 ;
        RECT 31.295 91.505 31.725 92.290 ;
        RECT 31.945 91.555 33.875 92.375 ;
        RECT 34.045 91.565 39.555 92.375 ;
        RECT 39.565 91.565 45.075 92.375 ;
        RECT 45.085 91.565 47.835 92.375 ;
        RECT 48.465 91.555 50.395 92.375 ;
        RECT 50.765 91.555 52.695 92.375 ;
        RECT 53.065 91.555 54.995 92.375 ;
        RECT 55.205 91.565 57.035 92.375 ;
        RECT 31.945 91.465 32.895 91.555 ;
        RECT 49.445 91.465 50.395 91.555 ;
        RECT 51.745 91.465 52.695 91.555 ;
        RECT 54.045 91.465 54.995 91.555 ;
        RECT 57.055 91.505 57.485 92.290 ;
        RECT 57.515 91.695 60.255 92.375 ;
        RECT 60.465 91.555 62.395 92.375 ;
        RECT 60.465 91.465 61.415 91.555 ;
        RECT 62.575 91.465 63.925 92.375 ;
        RECT 63.945 91.565 67.615 92.375 ;
        RECT 67.625 91.565 68.995 92.375 ;
        RECT 69.015 91.465 70.365 92.375 ;
        RECT 70.385 91.695 74.285 92.375 ;
        RECT 70.385 91.465 71.315 91.695 ;
        RECT 75.640 91.465 79.115 92.375 ;
        RECT 79.270 92.345 79.440 92.565 ;
        RECT 82.035 92.420 82.195 92.530 ;
        RECT 83.405 92.375 83.575 92.565 ;
        RECT 83.865 92.395 84.035 92.565 ;
        RECT 86.165 92.395 86.335 92.565 ;
        RECT 88.005 92.395 88.175 92.565 ;
        RECT 88.005 92.375 88.155 92.395 ;
        RECT 88.465 92.375 88.635 92.565 ;
        RECT 88.925 92.395 89.095 92.585 ;
        RECT 91.225 92.395 91.395 92.585 ;
        RECT 91.685 92.395 91.855 92.585 ;
        RECT 95.360 92.425 95.480 92.535 ;
        RECT 96.285 92.395 96.455 92.585 ;
        RECT 99.045 92.535 99.215 92.565 ;
        RECT 98.135 92.420 98.295 92.530 ;
        RECT 99.040 92.425 99.215 92.535 ;
        RECT 99.045 92.375 99.215 92.425 ;
        RECT 99.505 92.395 99.675 92.585 ;
        RECT 100.885 92.395 101.055 92.585 ;
        RECT 110.085 92.375 110.255 92.565 ;
        RECT 110.545 92.375 110.715 92.585 ;
        RECT 111.920 92.425 112.040 92.535 ;
        RECT 113.305 92.375 113.475 92.585 ;
        RECT 80.930 92.345 81.875 92.375 ;
        RECT 79.125 91.665 81.875 92.345 ;
        RECT 80.930 91.465 81.875 91.665 ;
        RECT 82.815 91.505 83.245 92.290 ;
        RECT 83.265 91.695 86.005 92.375 ;
        RECT 86.225 91.555 88.155 92.375 ;
        RECT 88.325 91.695 97.605 92.375 ;
        RECT 98.905 91.695 108.185 92.375 ;
        RECT 86.225 91.465 87.175 91.555 ;
        RECT 89.685 91.475 90.605 91.695 ;
        RECT 95.270 91.575 97.605 91.695 ;
        RECT 96.685 91.465 97.605 91.575 ;
        RECT 100.265 91.475 101.185 91.695 ;
        RECT 105.850 91.575 108.185 91.695 ;
        RECT 107.265 91.465 108.185 91.575 ;
        RECT 108.575 91.505 109.005 92.290 ;
        RECT 109.025 91.595 110.395 92.375 ;
        RECT 110.415 91.465 111.765 92.375 ;
        RECT 112.245 91.565 113.615 92.375 ;
      LAYER nwell ;
        RECT 5.330 88.345 113.810 91.175 ;
      LAYER pwell ;
        RECT 5.525 87.145 6.895 87.955 ;
        RECT 6.905 87.145 8.735 87.955 ;
        RECT 10.105 87.825 11.025 88.045 ;
        RECT 17.105 87.945 18.025 88.055 ;
        RECT 15.690 87.825 18.025 87.945 ;
        RECT 8.745 87.145 18.025 87.825 ;
        RECT 18.415 87.230 18.845 88.015 ;
        RECT 18.865 87.825 19.795 88.055 ;
        RECT 23.205 87.965 24.155 88.055 ;
        RECT 27.825 87.965 28.775 88.055 ;
        RECT 18.865 87.145 22.765 87.825 ;
        RECT 23.205 87.145 25.135 87.965 ;
        RECT 25.305 87.145 26.675 87.955 ;
        RECT 26.845 87.145 28.775 87.965 ;
        RECT 28.985 87.145 34.495 87.955 ;
        RECT 34.505 87.145 38.175 87.955 ;
        RECT 38.185 87.145 39.555 87.955 ;
        RECT 39.565 87.145 40.935 87.925 ;
        RECT 40.945 87.145 43.695 87.955 ;
        RECT 44.175 87.230 44.605 88.015 ;
        RECT 44.625 87.145 48.295 87.955 ;
        RECT 49.225 87.855 50.170 88.055 ;
        RECT 49.225 87.175 51.975 87.855 ;
        RECT 49.225 87.145 50.170 87.175 ;
        RECT 5.665 86.935 5.835 87.145 ;
        RECT 7.045 86.935 7.215 87.145 ;
        RECT 8.885 86.955 9.055 87.145 ;
        RECT 12.565 86.935 12.735 87.125 ;
        RECT 14.865 86.935 15.035 87.125 ;
        RECT 16.245 86.935 16.415 87.125 ;
        RECT 16.705 86.935 16.875 87.125 ;
        RECT 19.280 86.955 19.450 87.145 ;
        RECT 24.985 87.125 25.135 87.145 ;
        RECT 20.380 86.985 20.500 87.095 ;
        RECT 22.685 86.955 22.855 87.125 ;
        RECT 23.145 86.955 23.315 87.125 ;
        RECT 24.985 86.955 25.155 87.125 ;
        RECT 22.685 86.935 22.835 86.955 ;
        RECT 5.525 86.125 6.895 86.935 ;
        RECT 6.905 86.125 12.415 86.935 ;
        RECT 12.425 86.125 13.795 86.935 ;
        RECT 13.815 86.025 15.165 86.935 ;
        RECT 15.185 86.155 16.555 86.935 ;
        RECT 16.565 86.125 20.235 86.935 ;
        RECT 20.905 86.115 22.835 86.935 ;
        RECT 23.165 86.935 23.315 86.955 ;
        RECT 25.445 86.935 25.615 87.145 ;
        RECT 26.845 87.125 26.995 87.145 ;
        RECT 26.825 86.955 26.995 87.125 ;
        RECT 29.125 86.955 29.295 87.145 ;
        RECT 30.960 86.985 31.080 87.095 ;
        RECT 31.880 86.985 32.000 87.095 ;
        RECT 32.345 86.935 32.515 87.125 ;
        RECT 33.725 86.935 33.895 87.125 ;
        RECT 34.645 86.955 34.815 87.145 ;
        RECT 35.565 86.935 35.735 87.125 ;
        RECT 36.945 86.935 37.115 87.125 ;
        RECT 38.325 86.955 38.495 87.145 ;
        RECT 40.625 86.955 40.795 87.145 ;
        RECT 41.085 86.955 41.255 87.145 ;
        RECT 43.840 86.985 43.960 87.095 ;
        RECT 44.765 86.955 44.935 87.145 ;
        RECT 46.880 86.935 47.050 87.125 ;
        RECT 48.455 86.990 48.615 87.100 ;
        RECT 51.660 86.955 51.830 87.175 ;
        RECT 51.985 87.145 54.735 87.955 ;
        RECT 56.105 87.825 57.025 88.045 ;
        RECT 63.105 87.945 64.025 88.055 ;
        RECT 61.690 87.825 64.025 87.945 ;
        RECT 54.745 87.145 64.025 87.825 ;
        RECT 64.405 87.145 66.235 87.825 ;
        RECT 67.165 87.145 68.535 87.925 ;
        RECT 68.545 87.145 69.915 87.955 ;
        RECT 69.935 87.230 70.365 88.015 ;
        RECT 70.385 87.145 74.055 87.955 ;
        RECT 74.260 87.145 77.735 88.055 ;
        RECT 80.010 87.855 80.955 88.055 ;
        RECT 82.770 87.855 83.715 88.055 ;
        RECT 78.205 87.175 80.955 87.855 ;
        RECT 80.965 87.175 83.715 87.855 ;
        RECT 52.125 86.955 52.295 87.145 ;
        RECT 53.960 86.935 54.130 87.125 ;
        RECT 23.165 86.115 25.095 86.935 ;
        RECT 25.305 86.125 30.815 86.935 ;
        RECT 20.905 86.025 21.855 86.115 ;
        RECT 24.145 86.025 25.095 86.115 ;
        RECT 31.295 86.065 31.725 86.850 ;
        RECT 32.205 86.155 33.575 86.935 ;
        RECT 33.585 86.125 35.415 86.935 ;
        RECT 35.435 86.025 36.785 86.935 ;
        RECT 36.805 86.255 46.085 86.935 ;
        RECT 38.165 86.035 39.085 86.255 ;
        RECT 43.750 86.135 46.085 86.255 ;
        RECT 45.165 86.025 46.085 86.135 ;
        RECT 46.465 86.255 50.365 86.935 ;
        RECT 46.465 86.025 47.395 86.255 ;
        RECT 50.800 86.025 54.275 86.935 ;
        RECT 54.430 86.905 54.600 87.125 ;
        RECT 54.885 86.955 55.055 87.145 ;
        RECT 58.565 86.935 58.735 87.125 ;
        RECT 59.300 86.935 59.470 87.125 ;
        RECT 63.175 86.980 63.335 87.090 ;
        RECT 64.085 86.935 64.255 87.125 ;
        RECT 64.545 86.955 64.715 87.145 ;
        RECT 66.395 86.990 66.555 87.100 ;
        RECT 68.225 86.955 68.395 87.145 ;
        RECT 68.685 86.955 68.855 87.145 ;
        RECT 70.525 86.955 70.695 87.145 ;
        RECT 74.020 86.935 74.190 87.125 ;
        RECT 77.420 86.955 77.590 87.145 ;
        RECT 77.890 87.095 78.060 87.125 ;
        RECT 77.880 86.985 78.060 87.095 ;
        RECT 77.890 86.935 78.060 86.985 ;
        RECT 78.350 86.955 78.520 87.175 ;
        RECT 80.010 87.145 80.955 87.175 ;
        RECT 81.110 86.955 81.280 87.175 ;
        RECT 82.770 87.145 83.715 87.175 ;
        RECT 83.725 87.145 85.095 87.955 ;
        RECT 86.910 87.855 87.855 88.055 ;
        RECT 85.105 87.175 87.855 87.855 ;
        RECT 81.565 86.935 81.735 87.125 ;
        RECT 83.405 86.935 83.575 87.125 ;
        RECT 83.865 86.955 84.035 87.145 ;
        RECT 85.250 86.955 85.420 87.175 ;
        RECT 86.910 87.145 87.855 87.175 ;
        RECT 88.065 87.965 89.015 88.055 ;
        RECT 88.065 87.145 89.995 87.965 ;
        RECT 90.625 87.825 91.555 88.055 ;
        RECT 90.625 87.145 94.525 87.825 ;
        RECT 95.695 87.230 96.125 88.015 ;
        RECT 96.155 87.145 97.505 88.055 ;
        RECT 97.525 87.145 101.195 87.955 ;
        RECT 105.325 87.825 106.255 88.055 ;
        RECT 102.355 87.145 106.255 87.825 ;
        RECT 106.265 87.825 107.195 88.055 ;
        RECT 106.265 87.145 110.165 87.825 ;
        RECT 110.405 87.145 112.235 87.955 ;
        RECT 112.245 87.145 113.615 87.955 ;
        RECT 89.845 87.125 89.995 87.145 ;
        RECT 88.925 86.935 89.095 87.125 ;
        RECT 89.845 86.955 90.015 87.125 ;
        RECT 90.300 86.985 90.420 87.095 ;
        RECT 91.040 86.955 91.210 87.145 ;
        RECT 94.445 86.935 94.615 87.125 ;
        RECT 94.915 86.990 95.075 87.100 ;
        RECT 97.205 86.955 97.375 87.145 ;
        RECT 97.665 86.955 97.835 87.145 ;
        RECT 99.965 86.935 100.135 87.125 ;
        RECT 101.355 86.990 101.515 87.100 ;
        RECT 105.485 86.935 105.655 87.125 ;
        RECT 105.670 86.955 105.840 87.145 ;
        RECT 106.680 86.955 106.850 87.145 ;
        RECT 108.240 86.985 108.360 87.095 ;
        RECT 109.165 86.935 109.335 87.125 ;
        RECT 110.545 86.955 110.715 87.145 ;
        RECT 111.920 86.985 112.040 87.095 ;
        RECT 113.305 86.935 113.475 87.145 ;
        RECT 56.090 86.905 57.035 86.935 ;
        RECT 54.285 86.225 57.035 86.905 ;
        RECT 56.090 86.025 57.035 86.225 ;
        RECT 57.055 86.065 57.485 86.850 ;
        RECT 57.505 86.155 58.875 86.935 ;
        RECT 58.885 86.255 62.785 86.935 ;
        RECT 63.945 86.255 73.225 86.935 ;
        RECT 58.885 86.025 59.815 86.255 ;
        RECT 65.305 86.035 66.225 86.255 ;
        RECT 70.890 86.135 73.225 86.255 ;
        RECT 72.305 86.025 73.225 86.135 ;
        RECT 73.605 86.255 77.505 86.935 ;
        RECT 73.605 86.025 74.535 86.255 ;
        RECT 77.745 86.025 81.220 86.935 ;
        RECT 81.425 86.125 82.795 86.935 ;
        RECT 82.815 86.065 83.245 86.850 ;
        RECT 83.265 86.125 88.775 86.935 ;
        RECT 88.785 86.125 94.295 86.935 ;
        RECT 94.305 86.125 99.815 86.935 ;
        RECT 99.825 86.125 105.335 86.935 ;
        RECT 105.345 86.125 108.095 86.935 ;
        RECT 108.575 86.065 109.005 86.850 ;
        RECT 109.025 86.125 111.775 86.935 ;
        RECT 112.245 86.125 113.615 86.935 ;
      LAYER nwell ;
        RECT 5.330 82.905 113.810 85.735 ;
      LAYER pwell ;
        RECT 5.525 81.705 6.895 82.515 ;
        RECT 6.905 81.705 12.415 82.515 ;
        RECT 12.425 81.705 17.935 82.515 ;
        RECT 18.415 81.790 18.845 82.575 ;
        RECT 18.865 81.705 20.695 82.515 ;
        RECT 22.525 82.385 23.445 82.605 ;
        RECT 29.525 82.505 30.445 82.615 ;
        RECT 28.110 82.385 30.445 82.505 ;
        RECT 32.185 82.385 33.105 82.605 ;
        RECT 39.185 82.505 40.105 82.615 ;
        RECT 37.770 82.385 40.105 82.505 ;
        RECT 21.165 81.705 30.445 82.385 ;
        RECT 30.825 81.705 40.105 82.385 ;
        RECT 40.955 81.705 42.305 82.615 ;
        RECT 42.325 81.705 44.155 82.515 ;
        RECT 44.175 81.790 44.605 82.575 ;
        RECT 44.625 81.705 46.455 82.515 ;
        RECT 46.925 81.705 50.400 82.615 ;
        RECT 50.605 81.705 56.115 82.515 ;
        RECT 56.125 81.705 59.795 82.515 ;
        RECT 59.805 81.705 61.635 82.385 ;
        RECT 61.645 81.705 67.155 82.515 ;
        RECT 67.165 81.705 69.915 82.515 ;
        RECT 69.935 81.790 70.365 82.575 ;
        RECT 70.395 81.705 71.745 82.615 ;
        RECT 72.225 81.705 73.595 82.485 ;
        RECT 74.965 82.385 75.885 82.605 ;
        RECT 81.965 82.505 82.885 82.615 ;
        RECT 94.065 82.525 95.015 82.615 ;
        RECT 80.550 82.385 82.885 82.505 ;
        RECT 73.605 81.705 82.885 82.385 ;
        RECT 83.265 81.705 88.775 82.515 ;
        RECT 88.785 81.705 92.455 82.515 ;
        RECT 93.085 81.705 95.015 82.525 ;
        RECT 95.695 81.790 96.125 82.575 ;
        RECT 96.155 81.705 97.505 82.615 ;
        RECT 97.525 81.705 101.195 82.515 ;
        RECT 103.485 82.385 104.405 82.605 ;
        RECT 110.485 82.505 111.405 82.615 ;
        RECT 109.070 82.385 111.405 82.505 ;
        RECT 102.125 81.705 111.405 82.385 ;
        RECT 112.245 81.705 113.615 82.515 ;
        RECT 5.665 81.495 5.835 81.705 ;
        RECT 7.045 81.495 7.215 81.705 ;
        RECT 9.800 81.545 9.920 81.655 ;
        RECT 11.185 81.495 11.355 81.685 ;
        RECT 12.565 81.495 12.735 81.705 ;
        RECT 13.025 81.495 13.195 81.685 ;
        RECT 14.680 81.495 14.850 81.685 ;
        RECT 18.080 81.545 18.200 81.655 ;
        RECT 18.545 81.495 18.715 81.685 ;
        RECT 19.005 81.515 19.175 81.705 ;
        RECT 20.840 81.545 20.960 81.655 ;
        RECT 21.305 81.515 21.475 81.705 ;
        RECT 22.235 81.540 22.395 81.650 ;
        RECT 24.065 81.495 24.235 81.685 ;
        RECT 24.800 81.495 24.970 81.685 ;
        RECT 29.585 81.495 29.755 81.685 ;
        RECT 30.045 81.495 30.215 81.685 ;
        RECT 30.965 81.515 31.135 81.705 ;
        RECT 31.880 81.545 32.000 81.655 ;
        RECT 32.620 81.495 32.790 81.685 ;
        RECT 36.485 81.495 36.655 81.685 ;
        RECT 40.175 81.540 40.335 81.650 ;
        RECT 40.620 81.545 40.740 81.655 ;
        RECT 41.085 81.515 41.255 81.705 ;
        RECT 42.005 81.495 42.175 81.685 ;
        RECT 42.465 81.655 42.635 81.705 ;
        RECT 42.460 81.545 42.635 81.655 ;
        RECT 42.465 81.515 42.635 81.545 ;
        RECT 43.200 81.495 43.370 81.685 ;
        RECT 44.765 81.515 44.935 81.705 ;
        RECT 47.070 81.685 47.240 81.705 ;
        RECT 46.600 81.545 46.720 81.655 ;
        RECT 47.065 81.515 47.240 81.685 ;
        RECT 50.745 81.515 50.915 81.705 ;
        RECT 47.065 81.495 47.235 81.515 ;
        RECT 52.585 81.495 52.755 81.685 ;
        RECT 56.265 81.515 56.435 81.705 ;
        RECT 57.645 81.495 57.815 81.685 ;
        RECT 61.325 81.515 61.495 81.705 ;
        RECT 61.785 81.515 61.955 81.705 ;
        RECT 63.165 81.495 63.335 81.685 ;
        RECT 67.305 81.515 67.475 81.705 ;
        RECT 68.685 81.495 68.855 81.685 ;
        RECT 71.445 81.515 71.615 81.705 ;
        RECT 71.900 81.545 72.020 81.655 ;
        RECT 72.365 81.515 72.535 81.705 ;
        RECT 73.745 81.515 73.915 81.705 ;
        RECT 74.215 81.540 74.375 81.650 ;
        RECT 75.400 81.495 75.570 81.685 ;
        RECT 80.185 81.495 80.355 81.685 ;
        RECT 80.645 81.495 80.815 81.685 ;
        RECT 82.480 81.545 82.600 81.655 ;
        RECT 83.405 81.495 83.575 81.705 ;
        RECT 88.925 81.515 89.095 81.705 ;
        RECT 93.085 81.685 93.235 81.705 ;
        RECT 89.845 81.495 90.015 81.685 ;
        RECT 91.225 81.495 91.395 81.685 ;
        RECT 92.600 81.545 92.720 81.655 ;
        RECT 93.065 81.515 93.235 81.685 ;
        RECT 95.360 81.545 95.480 81.655 ;
        RECT 97.205 81.515 97.375 81.705 ;
        RECT 97.665 81.515 97.835 81.705 ;
        RECT 101.355 81.550 101.515 81.660 ;
        RECT 102.265 81.515 102.435 81.705 ;
        RECT 104.290 81.495 104.460 81.685 ;
        RECT 105.945 81.495 106.115 81.685 ;
        RECT 107.325 81.495 107.495 81.685 ;
        RECT 107.795 81.540 107.955 81.650 ;
        RECT 110.085 81.495 110.255 81.685 ;
        RECT 110.545 81.495 110.715 81.685 ;
        RECT 111.920 81.545 112.040 81.655 ;
        RECT 113.305 81.495 113.475 81.705 ;
        RECT 5.525 80.685 6.895 81.495 ;
        RECT 6.905 80.685 9.655 81.495 ;
        RECT 10.125 80.715 11.495 81.495 ;
        RECT 11.505 80.715 12.875 81.495 ;
        RECT 12.885 80.685 14.255 81.495 ;
        RECT 14.265 80.815 18.165 81.495 ;
        RECT 14.265 80.585 15.195 80.815 ;
        RECT 18.405 80.685 22.075 81.495 ;
        RECT 23.005 80.715 24.375 81.495 ;
        RECT 24.385 80.815 28.285 81.495 ;
        RECT 24.385 80.585 25.315 80.815 ;
        RECT 28.535 80.585 29.885 81.495 ;
        RECT 29.905 80.685 31.275 81.495 ;
        RECT 31.295 80.625 31.725 81.410 ;
        RECT 32.205 80.815 36.105 81.495 ;
        RECT 32.205 80.585 33.135 80.815 ;
        RECT 36.345 80.685 40.015 81.495 ;
        RECT 40.945 80.715 42.315 81.495 ;
        RECT 42.785 80.815 46.685 81.495 ;
        RECT 42.785 80.585 43.715 80.815 ;
        RECT 46.925 80.685 52.435 81.495 ;
        RECT 52.445 80.685 56.115 81.495 ;
        RECT 57.055 80.625 57.485 81.410 ;
        RECT 57.505 80.685 63.015 81.495 ;
        RECT 63.025 80.685 68.535 81.495 ;
        RECT 68.545 80.685 74.055 81.495 ;
        RECT 74.985 80.815 78.885 81.495 ;
        RECT 74.985 80.585 75.915 80.815 ;
        RECT 79.135 80.585 80.485 81.495 ;
        RECT 80.505 80.685 82.335 81.495 ;
        RECT 82.815 80.625 83.245 81.410 ;
        RECT 83.265 80.685 88.775 81.495 ;
        RECT 89.705 80.715 91.075 81.495 ;
        RECT 91.085 80.815 100.365 81.495 ;
        RECT 100.975 80.815 104.875 81.495 ;
        RECT 92.445 80.595 93.365 80.815 ;
        RECT 98.030 80.695 100.365 80.815 ;
        RECT 99.445 80.585 100.365 80.695 ;
        RECT 103.945 80.585 104.875 80.815 ;
        RECT 104.885 80.715 106.255 81.495 ;
        RECT 106.265 80.715 107.635 81.495 ;
        RECT 108.575 80.625 109.005 81.410 ;
        RECT 109.035 80.585 110.385 81.495 ;
        RECT 110.415 80.585 111.765 81.495 ;
        RECT 112.245 80.685 113.615 81.495 ;
      LAYER nwell ;
        RECT 5.330 77.465 113.810 80.295 ;
      LAYER pwell ;
        RECT 5.525 76.265 6.895 77.075 ;
        RECT 6.905 76.265 8.735 77.075 ;
        RECT 10.105 76.945 11.025 77.165 ;
        RECT 17.105 77.065 18.025 77.175 ;
        RECT 15.690 76.945 18.025 77.065 ;
        RECT 8.745 76.265 18.025 76.945 ;
        RECT 18.415 76.350 18.845 77.135 ;
        RECT 18.875 76.265 20.225 77.175 ;
        RECT 20.245 76.265 22.075 77.075 ;
        RECT 23.890 76.975 24.835 77.175 ;
        RECT 26.650 76.975 27.595 77.175 ;
        RECT 22.085 76.295 24.835 76.975 ;
        RECT 24.845 76.295 27.595 76.975 ;
        RECT 5.665 76.055 5.835 76.265 ;
        RECT 7.045 76.055 7.215 76.265 ;
        RECT 8.885 76.075 9.055 76.265 ;
        RECT 16.980 76.055 17.150 76.245 ;
        RECT 19.925 76.075 20.095 76.265 ;
        RECT 20.385 76.075 20.555 76.265 ;
        RECT 20.845 76.055 21.015 76.245 ;
        RECT 22.230 76.075 22.400 76.295 ;
        RECT 23.890 76.265 24.835 76.295 ;
        RECT 24.990 76.075 25.160 76.295 ;
        RECT 26.650 76.265 27.595 76.295 ;
        RECT 27.605 76.265 33.115 77.075 ;
        RECT 33.125 76.265 38.635 77.075 ;
        RECT 38.645 76.265 41.395 77.075 ;
        RECT 41.415 76.265 42.765 77.175 ;
        RECT 42.785 76.265 44.155 77.075 ;
        RECT 44.175 76.350 44.605 77.135 ;
        RECT 44.625 76.265 50.135 77.075 ;
        RECT 52.425 76.945 53.345 77.165 ;
        RECT 59.425 77.065 60.345 77.175 ;
        RECT 58.010 76.945 60.345 77.065 ;
        RECT 51.065 76.265 60.345 76.945 ;
        RECT 60.725 76.945 61.655 77.175 ;
        RECT 60.725 76.265 64.625 76.945 ;
        RECT 65.060 76.265 68.535 77.175 ;
        RECT 68.555 76.265 69.905 77.175 ;
        RECT 69.935 76.350 70.365 77.135 ;
        RECT 70.385 76.265 75.895 77.075 ;
        RECT 76.825 76.265 78.195 77.045 ;
        RECT 78.665 76.975 79.610 77.175 ;
        RECT 89.445 77.085 90.395 77.175 ;
        RECT 91.745 77.085 92.695 77.175 ;
        RECT 78.665 76.295 81.415 76.975 ;
        RECT 78.665 76.265 79.610 76.295 ;
        RECT 25.900 76.055 26.070 76.245 ;
        RECT 26.365 76.055 26.535 76.245 ;
        RECT 27.745 76.075 27.915 76.265 ;
        RECT 30.045 76.055 30.215 76.245 ;
        RECT 31.890 76.055 32.060 76.245 ;
        RECT 33.265 76.075 33.435 76.265 ;
        RECT 35.565 76.055 35.735 76.245 ;
        RECT 37.400 76.105 37.520 76.215 ;
        RECT 37.865 76.055 38.035 76.245 ;
        RECT 38.785 76.075 38.955 76.265 ;
        RECT 41.545 76.075 41.715 76.265 ;
        RECT 42.925 76.075 43.095 76.265 ;
        RECT 44.765 76.075 44.935 76.265 ;
        RECT 51.205 76.245 51.375 76.265 ;
        RECT 47.520 76.105 47.640 76.215 ;
        RECT 50.295 76.110 50.455 76.220 ;
        RECT 51.200 76.075 51.375 76.245 ;
        RECT 51.200 76.055 51.370 76.075 ;
        RECT 5.525 75.245 6.895 76.055 ;
        RECT 6.905 75.375 16.185 76.055 ;
        RECT 8.265 75.155 9.185 75.375 ;
        RECT 13.850 75.255 16.185 75.375 ;
        RECT 15.265 75.145 16.185 75.255 ;
        RECT 16.565 75.375 20.465 76.055 ;
        RECT 16.565 75.145 17.495 75.375 ;
        RECT 20.705 75.245 22.535 76.055 ;
        RECT 22.740 75.145 26.215 76.055 ;
        RECT 26.225 75.245 29.895 76.055 ;
        RECT 29.905 75.245 31.275 76.055 ;
        RECT 31.295 75.185 31.725 75.970 ;
        RECT 31.745 75.145 35.220 76.055 ;
        RECT 35.425 75.245 37.255 76.055 ;
        RECT 37.725 75.375 47.005 76.055 ;
        RECT 39.085 75.155 40.005 75.375 ;
        RECT 44.670 75.255 47.005 75.375 ;
        RECT 46.085 75.145 47.005 75.255 ;
        RECT 48.040 75.145 51.515 76.055 ;
        RECT 51.670 76.025 51.840 76.245 ;
        RECT 55.345 76.055 55.515 76.245 ;
        RECT 55.805 76.055 55.975 76.245 ;
        RECT 57.645 76.055 57.815 76.245 ;
        RECT 60.405 76.055 60.575 76.245 ;
        RECT 61.140 76.075 61.310 76.265 ;
        RECT 68.220 76.075 68.390 76.265 ;
        RECT 69.605 76.075 69.775 76.265 ;
        RECT 70.340 76.055 70.510 76.245 ;
        RECT 70.525 76.075 70.695 76.265 ;
        RECT 74.215 76.100 74.375 76.210 ;
        RECT 76.055 76.110 76.215 76.220 ;
        RECT 76.965 76.075 77.135 76.265 ;
        RECT 78.340 76.105 78.460 76.215 ;
        RECT 78.530 76.055 78.700 76.245 ;
        RECT 79.270 76.055 79.440 76.245 ;
        RECT 81.100 76.075 81.270 76.295 ;
        RECT 81.425 76.265 86.935 77.075 ;
        RECT 86.945 76.265 88.775 77.075 ;
        RECT 89.445 76.265 91.375 77.085 ;
        RECT 91.745 76.265 93.675 77.085 ;
        RECT 93.845 76.265 95.675 77.075 ;
        RECT 95.695 76.350 96.125 77.135 ;
        RECT 96.145 76.945 97.075 77.175 ;
        RECT 102.105 76.945 103.025 77.165 ;
        RECT 109.105 77.065 110.025 77.175 ;
        RECT 107.690 76.945 110.025 77.065 ;
        RECT 96.145 76.265 100.045 76.945 ;
        RECT 100.745 76.265 110.025 76.945 ;
        RECT 110.405 76.265 112.235 77.075 ;
        RECT 112.245 76.265 113.615 77.075 ;
        RECT 81.565 76.075 81.735 76.265 ;
        RECT 84.325 76.055 84.495 76.245 ;
        RECT 84.785 76.055 84.955 76.245 ;
        RECT 53.330 76.025 54.275 76.055 ;
        RECT 51.525 75.345 54.275 76.025 ;
        RECT 53.330 75.145 54.275 75.345 ;
        RECT 54.285 75.275 55.655 76.055 ;
        RECT 55.675 75.145 57.025 76.055 ;
        RECT 57.055 75.185 57.485 75.970 ;
        RECT 57.505 75.245 60.255 76.055 ;
        RECT 60.265 75.375 69.545 76.055 ;
        RECT 61.625 75.155 62.545 75.375 ;
        RECT 67.210 75.255 69.545 75.375 ;
        RECT 68.625 75.145 69.545 75.255 ;
        RECT 69.925 75.375 73.825 76.055 ;
        RECT 75.215 75.375 79.115 76.055 ;
        RECT 69.925 75.145 70.855 75.375 ;
        RECT 78.185 75.145 79.115 75.375 ;
        RECT 79.125 75.145 82.600 76.055 ;
        RECT 82.815 75.185 83.245 75.970 ;
        RECT 83.275 75.145 84.625 76.055 ;
        RECT 84.645 75.245 86.475 76.055 ;
        RECT 86.630 76.025 86.800 76.245 ;
        RECT 87.085 76.075 87.255 76.265 ;
        RECT 91.225 76.245 91.375 76.265 ;
        RECT 93.525 76.245 93.675 76.265 ;
        RECT 93.985 76.245 94.155 76.265 ;
        RECT 88.920 76.105 89.040 76.215 ;
        RECT 89.385 76.055 89.555 76.245 ;
        RECT 91.225 76.075 91.400 76.245 ;
        RECT 93.525 76.075 93.695 76.245 ;
        RECT 93.985 76.075 94.160 76.245 ;
        RECT 96.560 76.075 96.730 76.265 ;
        RECT 88.290 76.025 89.235 76.055 ;
        RECT 86.485 75.345 89.235 76.025 ;
        RECT 88.290 75.145 89.235 75.345 ;
        RECT 89.245 75.245 91.075 76.055 ;
        RECT 91.230 76.025 91.400 76.075 ;
        RECT 92.890 76.025 93.835 76.055 ;
        RECT 93.990 76.025 94.160 76.075 ;
        RECT 95.650 76.025 96.595 76.055 ;
        RECT 96.750 76.025 96.920 76.245 ;
        RECT 99.505 76.055 99.675 76.245 ;
        RECT 100.420 76.105 100.540 76.215 ;
        RECT 100.885 76.075 101.055 76.265 ;
        RECT 103.195 76.100 103.355 76.210 ;
        RECT 107.510 76.055 107.680 76.245 ;
        RECT 108.240 76.105 108.360 76.215 ;
        RECT 109.165 76.055 109.335 76.245 ;
        RECT 110.545 76.075 110.715 76.265 ;
        RECT 111.920 76.105 112.040 76.215 ;
        RECT 113.305 76.055 113.475 76.265 ;
        RECT 98.410 76.025 99.355 76.055 ;
        RECT 91.085 75.345 93.835 76.025 ;
        RECT 93.845 75.345 96.595 76.025 ;
        RECT 96.605 75.345 99.355 76.025 ;
        RECT 92.890 75.145 93.835 75.345 ;
        RECT 95.650 75.145 96.595 75.345 ;
        RECT 98.410 75.145 99.355 75.345 ;
        RECT 99.365 75.245 103.035 76.055 ;
        RECT 104.195 75.375 108.095 76.055 ;
        RECT 107.165 75.145 108.095 75.375 ;
        RECT 108.575 75.185 109.005 75.970 ;
        RECT 109.025 75.245 111.775 76.055 ;
        RECT 112.245 75.245 113.615 76.055 ;
      LAYER nwell ;
        RECT 5.330 72.025 113.810 74.855 ;
      LAYER pwell ;
        RECT 5.525 70.825 6.895 71.635 ;
        RECT 6.905 70.825 10.575 71.635 ;
        RECT 10.585 70.825 11.955 71.635 ;
        RECT 11.975 70.825 13.325 71.735 ;
        RECT 13.345 70.825 17.015 71.635 ;
        RECT 17.025 70.825 18.395 71.635 ;
        RECT 18.415 70.910 18.845 71.695 ;
        RECT 18.865 70.825 20.695 71.635 ;
        RECT 20.705 70.825 24.180 71.735 ;
        RECT 24.580 70.825 28.055 71.735 ;
        RECT 29.870 71.535 30.815 71.735 ;
        RECT 33.550 71.535 34.495 71.735 ;
        RECT 28.065 70.855 30.815 71.535 ;
        RECT 31.745 70.855 34.495 71.535 ;
        RECT 35.865 71.505 36.785 71.725 ;
        RECT 42.865 71.625 43.785 71.735 ;
        RECT 41.450 71.505 43.785 71.625 ;
        RECT 5.665 70.615 5.835 70.825 ;
        RECT 7.045 70.615 7.215 70.825 ;
        RECT 10.725 70.635 10.895 70.825 ;
        RECT 12.560 70.665 12.680 70.775 ;
        RECT 13.025 70.635 13.195 70.825 ;
        RECT 13.300 70.615 13.470 70.805 ;
        RECT 13.485 70.635 13.655 70.825 ;
        RECT 17.165 70.635 17.335 70.825 ;
        RECT 19.005 70.635 19.175 70.825 ;
        RECT 5.525 69.805 6.895 70.615 ;
        RECT 6.905 69.805 12.415 70.615 ;
        RECT 12.885 69.935 16.785 70.615 ;
        RECT 17.945 70.585 18.890 70.615 ;
        RECT 20.380 70.585 20.550 70.805 ;
        RECT 20.850 70.615 21.020 70.825 ;
        RECT 24.535 70.660 24.695 70.770 ;
        RECT 27.740 70.635 27.910 70.825 ;
        RECT 28.210 70.635 28.380 70.855 ;
        RECT 29.870 70.825 30.815 70.855 ;
        RECT 28.660 70.615 28.830 70.805 ;
        RECT 29.125 70.615 29.295 70.805 ;
        RECT 30.975 70.775 31.135 70.780 ;
        RECT 30.960 70.670 31.135 70.775 ;
        RECT 30.960 70.665 31.080 70.670 ;
        RECT 12.885 69.705 13.815 69.935 ;
        RECT 17.945 69.905 20.695 70.585 ;
        RECT 17.945 69.705 18.890 69.905 ;
        RECT 20.705 69.705 24.180 70.615 ;
        RECT 25.500 69.705 28.975 70.615 ;
        RECT 28.985 69.805 30.815 70.615 ;
        RECT 31.890 70.585 32.060 70.855 ;
        RECT 33.550 70.825 34.495 70.855 ;
        RECT 34.505 70.825 43.785 71.505 ;
        RECT 44.175 70.910 44.605 71.695 ;
        RECT 44.625 71.505 45.555 71.735 ;
        RECT 44.625 70.825 48.525 71.505 ;
        RECT 48.960 70.825 52.435 71.735 ;
        RECT 52.445 70.825 55.195 71.635 ;
        RECT 55.665 70.825 58.405 71.505 ;
        RECT 58.620 70.825 62.095 71.735 ;
        RECT 62.300 70.825 65.775 71.735 ;
        RECT 65.980 70.825 69.455 71.735 ;
        RECT 69.935 70.910 70.365 71.695 ;
        RECT 70.385 70.825 71.755 71.605 ;
        RECT 72.880 70.825 76.355 71.735 ;
        RECT 78.185 71.505 79.105 71.725 ;
        RECT 85.185 71.625 86.105 71.735 ;
        RECT 93.605 71.645 94.555 71.735 ;
        RECT 83.770 71.505 86.105 71.625 ;
        RECT 76.825 70.825 86.105 71.505 ;
        RECT 86.485 70.825 91.995 71.635 ;
        RECT 92.625 70.825 94.555 71.645 ;
        RECT 95.695 70.910 96.125 71.695 ;
        RECT 96.145 70.825 101.655 71.635 ;
        RECT 101.665 70.825 107.175 71.635 ;
        RECT 107.185 70.825 110.855 71.635 ;
        RECT 110.865 70.825 112.235 71.635 ;
        RECT 112.245 70.825 113.615 71.635 ;
        RECT 34.645 70.615 34.815 70.825 ;
        RECT 36.480 70.665 36.600 70.775 ;
        RECT 37.865 70.615 38.035 70.805 ;
        RECT 38.335 70.660 38.495 70.770 ;
        RECT 39.520 70.615 39.690 70.805 ;
        RECT 44.305 70.615 44.475 70.805 ;
        RECT 44.765 70.615 44.935 70.805 ;
        RECT 45.040 70.635 45.210 70.825 ;
        RECT 46.145 70.615 46.315 70.805 ;
        RECT 49.820 70.665 49.940 70.775 ;
        RECT 33.550 70.585 34.495 70.615 ;
        RECT 31.295 69.745 31.725 70.530 ;
        RECT 31.745 69.905 34.495 70.585 ;
        RECT 33.550 69.705 34.495 69.905 ;
        RECT 34.505 69.805 36.335 70.615 ;
        RECT 36.805 69.835 38.175 70.615 ;
        RECT 39.105 69.935 43.005 70.615 ;
        RECT 39.105 69.705 40.035 69.935 ;
        RECT 43.245 69.835 44.615 70.615 ;
        RECT 44.635 69.705 45.985 70.615 ;
        RECT 46.005 69.805 49.675 70.615 ;
        RECT 50.290 70.585 50.460 70.805 ;
        RECT 52.120 70.635 52.290 70.825 ;
        RECT 52.585 70.635 52.755 70.825 ;
        RECT 55.345 70.775 55.515 70.805 ;
        RECT 55.340 70.665 55.515 70.775 ;
        RECT 55.345 70.615 55.515 70.665 ;
        RECT 55.805 70.615 55.975 70.825 ;
        RECT 57.645 70.615 57.815 70.805 ;
        RECT 60.405 70.615 60.575 70.805 ;
        RECT 60.860 70.665 60.980 70.775 ;
        RECT 61.780 70.635 61.950 70.825 ;
        RECT 64.085 70.615 64.255 70.805 ;
        RECT 64.545 70.615 64.715 70.805 ;
        RECT 65.460 70.635 65.630 70.825 ;
        RECT 67.300 70.665 67.420 70.775 ;
        RECT 67.765 70.615 67.935 70.805 ;
        RECT 69.140 70.635 69.310 70.825 ;
        RECT 69.600 70.665 69.720 70.775 ;
        RECT 71.445 70.635 71.615 70.825 ;
        RECT 71.915 70.670 72.075 70.780 ;
        RECT 76.040 70.635 76.210 70.825 ;
        RECT 76.500 70.665 76.620 70.775 ;
        RECT 76.965 70.635 77.135 70.825 ;
        RECT 51.950 70.585 52.895 70.615 ;
        RECT 50.145 69.905 52.895 70.585 ;
        RECT 52.915 69.935 55.655 70.615 ;
        RECT 51.950 69.705 52.895 69.905 ;
        RECT 55.665 69.805 57.035 70.615 ;
        RECT 57.055 69.745 57.485 70.530 ;
        RECT 57.505 69.805 58.875 70.615 ;
        RECT 58.885 69.935 60.715 70.615 ;
        RECT 58.885 69.705 60.230 69.935 ;
        RECT 61.185 69.705 64.395 70.615 ;
        RECT 64.405 69.805 67.155 70.615 ;
        RECT 67.625 69.935 76.815 70.615 ;
        RECT 72.135 69.715 73.065 69.935 ;
        RECT 75.895 69.705 76.815 69.935 ;
        RECT 76.825 70.585 77.770 70.615 ;
        RECT 79.260 70.585 79.430 70.805 ;
        RECT 79.725 70.615 79.895 70.805 ;
        RECT 82.480 70.665 82.600 70.775 ;
        RECT 83.405 70.615 83.575 70.805 ;
        RECT 86.625 70.635 86.795 70.825 ;
        RECT 92.625 70.805 92.775 70.825 ;
        RECT 88.925 70.615 89.095 70.805 ;
        RECT 92.140 70.665 92.260 70.775 ;
        RECT 92.605 70.635 92.775 70.805 ;
        RECT 93.520 70.615 93.690 70.805 ;
        RECT 93.985 70.615 94.155 70.805 ;
        RECT 94.915 70.670 95.075 70.780 ;
        RECT 96.285 70.635 96.455 70.825 ;
        RECT 99.500 70.665 99.620 70.775 ;
        RECT 99.965 70.615 100.135 70.805 ;
        RECT 101.345 70.615 101.515 70.805 ;
        RECT 101.805 70.635 101.975 70.825 ;
        RECT 103.185 70.615 103.355 70.805 ;
        RECT 104.560 70.665 104.680 70.775 ;
        RECT 105.945 70.615 106.115 70.805 ;
        RECT 106.405 70.615 106.575 70.805 ;
        RECT 107.325 70.635 107.495 70.825 ;
        RECT 108.240 70.665 108.360 70.775 ;
        RECT 109.165 70.615 109.335 70.805 ;
        RECT 111.005 70.635 111.175 70.825 ;
        RECT 111.920 70.665 112.040 70.775 ;
        RECT 113.305 70.615 113.475 70.825 ;
        RECT 76.825 69.905 79.575 70.585 ;
        RECT 76.825 69.705 77.770 69.905 ;
        RECT 79.585 69.805 82.335 70.615 ;
        RECT 82.815 69.745 83.245 70.530 ;
        RECT 83.265 69.805 88.775 70.615 ;
        RECT 88.785 69.805 90.155 70.615 ;
        RECT 90.360 69.705 93.835 70.615 ;
        RECT 93.845 69.805 99.355 70.615 ;
        RECT 99.825 69.835 101.195 70.615 ;
        RECT 101.205 69.805 103.035 70.615 ;
        RECT 103.045 69.835 104.415 70.615 ;
        RECT 104.895 69.705 106.245 70.615 ;
        RECT 106.265 69.805 108.095 70.615 ;
        RECT 108.575 69.745 109.005 70.530 ;
        RECT 109.025 69.805 111.775 70.615 ;
        RECT 112.245 69.805 113.615 70.615 ;
      LAYER nwell ;
        RECT 5.330 66.585 113.810 69.415 ;
      LAYER pwell ;
        RECT 5.525 65.385 6.895 66.195 ;
        RECT 6.905 65.385 9.655 66.195 ;
        RECT 9.665 65.385 11.035 66.165 ;
        RECT 11.045 65.385 12.415 66.165 ;
        RECT 12.435 65.385 13.785 66.295 ;
        RECT 14.265 66.065 15.195 66.295 ;
        RECT 14.265 65.385 18.165 66.065 ;
        RECT 18.415 65.470 18.845 66.255 ;
        RECT 18.865 65.385 21.615 66.195 ;
        RECT 21.820 65.385 25.295 66.295 ;
        RECT 25.305 65.385 27.135 66.195 ;
        RECT 27.800 65.385 31.275 66.295 ;
        RECT 31.285 65.385 34.035 66.195 ;
        RECT 38.555 66.065 39.485 66.285 ;
        RECT 42.315 66.065 43.235 66.295 ;
        RECT 34.045 65.385 43.235 66.065 ;
        RECT 44.175 65.470 44.605 66.255 ;
        RECT 44.625 65.385 50.135 66.195 ;
        RECT 50.800 65.385 54.275 66.295 ;
        RECT 54.775 65.385 57.495 66.295 ;
        RECT 57.505 66.065 58.850 66.295 ;
        RECT 57.505 65.385 59.335 66.065 ;
        RECT 59.345 65.385 68.450 66.065 ;
        RECT 68.545 65.385 69.915 66.195 ;
        RECT 69.935 65.470 70.365 66.255 ;
        RECT 70.385 65.385 72.215 66.195 ;
        RECT 72.695 65.385 74.045 66.295 ;
        RECT 74.065 65.385 79.575 66.195 ;
        RECT 79.585 65.385 83.255 66.195 ;
        RECT 84.380 65.385 87.855 66.295 ;
        RECT 87.865 65.385 90.615 66.195 ;
        RECT 90.820 65.385 94.295 66.295 ;
        RECT 94.315 65.385 95.665 66.295 ;
        RECT 95.695 65.470 96.125 66.255 ;
        RECT 96.340 65.385 99.815 66.295 ;
        RECT 101.185 66.065 102.105 66.285 ;
        RECT 108.185 66.185 109.105 66.295 ;
        RECT 106.770 66.065 109.105 66.185 ;
        RECT 99.825 65.385 109.105 66.065 ;
        RECT 109.495 65.385 110.845 66.295 ;
        RECT 110.865 65.385 112.235 66.195 ;
        RECT 112.245 65.385 113.615 66.195 ;
        RECT 5.665 65.175 5.835 65.385 ;
        RECT 7.045 65.175 7.215 65.385 ;
        RECT 10.725 65.195 10.895 65.385 ;
        RECT 12.105 65.195 12.275 65.385 ;
        RECT 13.485 65.195 13.655 65.385 ;
        RECT 13.940 65.225 14.060 65.335 ;
        RECT 14.680 65.195 14.850 65.385 ;
        RECT 17.625 65.175 17.795 65.365 ;
        RECT 18.085 65.175 18.255 65.365 ;
        RECT 19.005 65.195 19.175 65.385 ;
        RECT 20.850 65.175 21.020 65.365 ;
        RECT 24.980 65.195 25.150 65.385 ;
        RECT 25.445 65.195 25.615 65.385 ;
        RECT 27.280 65.225 27.400 65.335 ;
        RECT 27.740 65.175 27.910 65.365 ;
        RECT 28.205 65.175 28.375 65.365 ;
        RECT 30.960 65.195 31.130 65.385 ;
        RECT 31.425 65.195 31.595 65.385 ;
        RECT 31.890 65.175 32.060 65.365 ;
        RECT 34.185 65.195 34.355 65.385 ;
        RECT 35.565 65.175 35.735 65.365 ;
        RECT 39.245 65.175 39.415 65.365 ;
        RECT 40.625 65.175 40.795 65.365 ;
        RECT 43.395 65.230 43.555 65.340 ;
        RECT 44.765 65.195 44.935 65.385 ;
        RECT 46.145 65.175 46.315 65.365 ;
        RECT 49.835 65.220 49.995 65.330 ;
        RECT 50.280 65.225 50.400 65.335 ;
        RECT 50.750 65.175 50.920 65.365 ;
        RECT 53.960 65.195 54.130 65.385 ;
        RECT 54.420 65.330 54.540 65.335 ;
        RECT 54.420 65.225 54.595 65.330 ;
        RECT 54.435 65.220 54.595 65.225 ;
        RECT 56.725 65.175 56.895 65.365 ;
        RECT 57.185 65.195 57.355 65.385 ;
        RECT 57.640 65.225 57.760 65.335 ;
        RECT 59.025 65.195 59.195 65.385 ;
        RECT 59.485 65.175 59.655 65.385 ;
        RECT 59.945 65.175 60.115 65.365 ;
        RECT 61.785 65.175 61.955 65.365 ;
        RECT 63.625 65.175 63.795 65.365 ;
        RECT 66.385 65.175 66.555 65.365 ;
        RECT 66.845 65.175 67.015 65.365 ;
        RECT 68.685 65.195 68.855 65.385 ;
        RECT 70.525 65.195 70.695 65.385 ;
        RECT 72.360 65.225 72.480 65.335 ;
        RECT 72.825 65.195 72.995 65.385 ;
        RECT 73.740 65.175 73.910 65.365 ;
        RECT 74.205 65.175 74.375 65.385 ;
        RECT 79.725 65.175 79.895 65.385 ;
        RECT 82.480 65.225 82.600 65.335 ;
        RECT 83.410 65.175 83.580 65.365 ;
        RECT 87.085 65.175 87.255 65.365 ;
        RECT 87.540 65.195 87.710 65.385 ;
        RECT 88.005 65.195 88.175 65.385 ;
        RECT 88.465 65.175 88.635 65.365 ;
        RECT 89.845 65.175 90.015 65.365 ;
        RECT 93.980 65.195 94.150 65.385 ;
        RECT 94.445 65.195 94.615 65.385 ;
        RECT 99.500 65.195 99.670 65.385 ;
        RECT 99.780 65.175 99.950 65.365 ;
        RECT 99.965 65.195 100.135 65.385 ;
        RECT 103.920 65.175 104.090 65.365 ;
        RECT 107.795 65.220 107.955 65.330 ;
        RECT 109.165 65.175 109.335 65.365 ;
        RECT 109.625 65.195 109.795 65.385 ;
        RECT 111.005 65.195 111.175 65.385 ;
        RECT 111.920 65.225 112.040 65.335 ;
        RECT 113.305 65.175 113.475 65.385 ;
        RECT 5.525 64.365 6.895 65.175 ;
        RECT 6.905 64.495 16.185 65.175 ;
        RECT 8.265 64.275 9.185 64.495 ;
        RECT 13.850 64.375 16.185 64.495 ;
        RECT 15.265 64.265 16.185 64.375 ;
        RECT 16.575 64.265 17.925 65.175 ;
        RECT 17.945 64.365 20.695 65.175 ;
        RECT 20.705 64.265 24.180 65.175 ;
        RECT 24.580 64.265 28.055 65.175 ;
        RECT 28.065 64.365 30.815 65.175 ;
        RECT 31.295 64.305 31.725 65.090 ;
        RECT 31.745 64.265 35.220 65.175 ;
        RECT 35.425 64.365 39.095 65.175 ;
        RECT 39.115 64.265 40.465 65.175 ;
        RECT 40.485 64.365 45.995 65.175 ;
        RECT 46.005 64.365 49.675 65.175 ;
        RECT 50.605 64.265 54.080 65.175 ;
        RECT 55.205 64.495 57.035 65.175 ;
        RECT 55.205 64.265 56.550 64.495 ;
        RECT 57.055 64.305 57.485 65.090 ;
        RECT 57.965 64.495 59.795 65.175 ;
        RECT 59.805 64.495 61.635 65.175 ;
        RECT 61.645 64.495 63.475 65.175 ;
        RECT 63.485 64.495 65.315 65.175 ;
        RECT 57.965 64.265 59.310 64.495 ;
        RECT 60.290 64.265 61.635 64.495 ;
        RECT 62.130 64.265 63.475 64.495 ;
        RECT 63.970 64.265 65.315 64.495 ;
        RECT 65.325 64.395 66.695 65.175 ;
        RECT 66.705 64.365 70.375 65.175 ;
        RECT 70.580 64.265 74.055 65.175 ;
        RECT 74.065 64.365 79.575 65.175 ;
        RECT 79.585 64.365 82.335 65.175 ;
        RECT 82.815 64.305 83.245 65.090 ;
        RECT 83.265 64.265 86.740 65.175 ;
        RECT 86.945 64.365 88.315 65.175 ;
        RECT 88.325 64.395 89.695 65.175 ;
        RECT 89.705 64.495 98.985 65.175 ;
        RECT 91.065 64.275 91.985 64.495 ;
        RECT 96.650 64.375 98.985 64.495 ;
        RECT 98.065 64.265 98.985 64.375 ;
        RECT 99.365 64.495 103.265 65.175 ;
        RECT 103.505 64.495 107.405 65.175 ;
        RECT 99.365 64.265 100.295 64.495 ;
        RECT 103.505 64.265 104.435 64.495 ;
        RECT 108.575 64.305 109.005 65.090 ;
        RECT 109.025 64.365 111.775 65.175 ;
        RECT 112.245 64.365 113.615 65.175 ;
      LAYER nwell ;
        RECT 5.330 61.145 113.810 63.975 ;
      LAYER pwell ;
        RECT 5.525 59.945 6.895 60.755 ;
        RECT 12.335 60.625 13.265 60.845 ;
        RECT 16.095 60.625 17.015 60.855 ;
        RECT 7.825 59.945 17.015 60.625 ;
        RECT 17.025 59.945 18.395 60.755 ;
        RECT 18.415 60.030 18.845 60.815 ;
        RECT 18.865 59.945 20.695 60.755 ;
        RECT 21.360 59.945 24.835 60.855 ;
        RECT 24.845 59.945 30.355 60.755 ;
        RECT 30.365 59.945 35.875 60.755 ;
        RECT 35.885 59.945 41.395 60.755 ;
        RECT 41.405 59.945 44.155 60.755 ;
        RECT 44.175 60.030 44.605 60.815 ;
        RECT 45.985 60.625 46.905 60.845 ;
        RECT 52.985 60.745 53.905 60.855 ;
        RECT 51.570 60.625 53.905 60.745 ;
        RECT 44.625 59.945 53.905 60.625 ;
        RECT 54.285 59.945 57.760 60.855 ;
        RECT 57.965 59.945 59.795 60.755 ;
        RECT 60.290 60.625 61.635 60.855 ;
        RECT 62.130 60.625 63.475 60.855 ;
        RECT 59.805 59.945 61.635 60.625 ;
        RECT 61.645 59.945 63.475 60.625 ;
        RECT 64.405 60.625 65.335 60.855 ;
        RECT 64.405 59.945 68.305 60.625 ;
        RECT 68.545 59.945 69.915 60.725 ;
        RECT 69.935 60.030 70.365 60.815 ;
        RECT 70.385 59.945 75.895 60.755 ;
        RECT 76.100 59.945 79.575 60.855 ;
        RECT 79.585 59.945 83.060 60.855 ;
        RECT 83.265 59.945 86.740 60.855 ;
        RECT 86.945 59.945 90.615 60.755 ;
        RECT 90.625 60.625 91.555 60.855 ;
        RECT 90.625 59.945 94.525 60.625 ;
        RECT 95.695 60.030 96.125 60.815 ;
        RECT 96.145 59.945 101.655 60.755 ;
        RECT 103.485 60.625 104.405 60.845 ;
        RECT 110.485 60.745 111.405 60.855 ;
        RECT 109.070 60.625 111.405 60.745 ;
        RECT 102.125 59.945 111.405 60.625 ;
        RECT 112.245 59.945 113.615 60.755 ;
        RECT 5.665 59.735 5.835 59.945 ;
        RECT 7.045 59.735 7.215 59.925 ;
        RECT 7.965 59.755 8.135 59.945 ;
        RECT 12.565 59.735 12.735 59.925 ;
        RECT 16.240 59.735 16.410 59.925 ;
        RECT 16.705 59.735 16.875 59.925 ;
        RECT 17.165 59.755 17.335 59.945 ;
        RECT 19.005 59.755 19.175 59.945 ;
        RECT 20.840 59.785 20.960 59.895 ;
        RECT 22.225 59.735 22.395 59.925 ;
        RECT 24.520 59.755 24.690 59.945 ;
        RECT 24.985 59.755 25.155 59.945 ;
        RECT 25.900 59.785 26.020 59.895 ;
        RECT 26.640 59.735 26.810 59.925 ;
        RECT 30.505 59.755 30.675 59.945 ;
        RECT 31.885 59.735 32.055 59.925 ;
        RECT 34.920 59.735 35.090 59.925 ;
        RECT 36.025 59.755 36.195 59.945 ;
        RECT 38.785 59.735 38.955 59.925 ;
        RECT 41.545 59.755 41.715 59.945 ;
        RECT 42.465 59.735 42.635 59.925 ;
        RECT 43.845 59.735 44.015 59.925 ;
        RECT 44.765 59.755 44.935 59.945 ;
        RECT 45.500 59.735 45.670 59.925 ;
        RECT 49.360 59.785 49.480 59.895 ;
        RECT 49.830 59.735 50.000 59.925 ;
        RECT 53.505 59.735 53.675 59.925 ;
        RECT 54.430 59.755 54.600 59.945 ;
        RECT 57.655 59.780 57.815 59.890 ;
        RECT 58.105 59.755 58.275 59.945 ;
        RECT 59.945 59.735 60.115 59.945 ;
        RECT 60.405 59.735 60.575 59.925 ;
        RECT 61.785 59.755 61.955 59.945 ;
        RECT 63.635 59.790 63.795 59.900 ;
        RECT 64.820 59.755 64.990 59.945 ;
        RECT 68.685 59.755 68.855 59.945 ;
        RECT 69.880 59.735 70.050 59.925 ;
        RECT 70.525 59.755 70.695 59.945 ;
        RECT 73.740 59.785 73.860 59.895 ;
        RECT 77.610 59.735 77.780 59.925 ;
        RECT 78.345 59.735 78.515 59.925 ;
        RECT 79.260 59.755 79.430 59.945 ;
        RECT 79.730 59.755 79.900 59.945 ;
        RECT 82.035 59.780 82.195 59.890 ;
        RECT 83.410 59.755 83.580 59.945 ;
        RECT 86.620 59.735 86.790 59.925 ;
        RECT 87.085 59.735 87.255 59.945 ;
        RECT 91.040 59.755 91.210 59.945 ;
        RECT 92.605 59.735 92.775 59.925 ;
        RECT 94.915 59.790 95.075 59.900 ;
        RECT 96.285 59.755 96.455 59.945 ;
        RECT 98.125 59.735 98.295 59.925 ;
        RECT 101.160 59.735 101.330 59.925 ;
        RECT 101.800 59.785 101.920 59.895 ;
        RECT 102.265 59.755 102.435 59.945 ;
        RECT 105.945 59.735 106.115 59.925 ;
        RECT 106.405 59.735 106.575 59.925 ;
        RECT 108.240 59.785 108.360 59.895 ;
        RECT 109.165 59.735 109.335 59.925 ;
        RECT 111.920 59.785 112.040 59.895 ;
        RECT 113.305 59.735 113.475 59.945 ;
        RECT 5.525 58.925 6.895 59.735 ;
        RECT 6.905 58.925 12.415 59.735 ;
        RECT 12.425 58.925 13.795 59.735 ;
        RECT 13.945 58.825 16.555 59.735 ;
        RECT 16.565 58.925 22.075 59.735 ;
        RECT 22.085 58.925 25.755 59.735 ;
        RECT 26.225 59.055 30.125 59.735 ;
        RECT 26.225 58.825 27.155 59.055 ;
        RECT 31.295 58.865 31.725 59.650 ;
        RECT 31.745 58.925 34.495 59.735 ;
        RECT 34.505 59.055 38.405 59.735 ;
        RECT 34.505 58.825 35.435 59.055 ;
        RECT 38.645 58.925 42.315 59.735 ;
        RECT 42.325 58.955 43.695 59.735 ;
        RECT 43.715 58.825 45.065 59.735 ;
        RECT 45.085 59.055 48.985 59.735 ;
        RECT 45.085 58.825 46.015 59.055 ;
        RECT 49.685 58.825 53.160 59.735 ;
        RECT 53.365 58.925 57.035 59.735 ;
        RECT 57.055 58.865 57.485 59.650 ;
        RECT 58.425 59.055 60.255 59.735 ;
        RECT 60.265 59.055 69.455 59.735 ;
        RECT 58.425 58.825 59.770 59.055 ;
        RECT 64.775 58.835 65.705 59.055 ;
        RECT 68.535 58.825 69.455 59.055 ;
        RECT 69.465 59.055 73.365 59.735 ;
        RECT 74.295 59.055 78.195 59.735 ;
        RECT 69.465 58.825 70.395 59.055 ;
        RECT 77.265 58.825 78.195 59.055 ;
        RECT 78.205 58.925 81.875 59.735 ;
        RECT 82.815 58.865 83.245 59.650 ;
        RECT 83.460 58.825 86.935 59.735 ;
        RECT 86.945 58.925 92.455 59.735 ;
        RECT 92.465 58.925 97.975 59.735 ;
        RECT 97.985 58.925 100.735 59.735 ;
        RECT 100.745 59.055 104.645 59.735 ;
        RECT 100.745 58.825 101.675 59.055 ;
        RECT 104.895 58.825 106.245 59.735 ;
        RECT 106.265 58.925 108.095 59.735 ;
        RECT 108.575 58.865 109.005 59.650 ;
        RECT 109.025 58.925 111.775 59.735 ;
        RECT 112.245 58.925 113.615 59.735 ;
      LAYER nwell ;
        RECT 5.330 55.705 113.810 58.535 ;
      LAYER pwell ;
        RECT 5.525 54.505 6.895 55.315 ;
        RECT 6.905 54.505 10.575 55.315 ;
        RECT 11.045 54.505 12.415 55.285 ;
        RECT 12.885 54.505 15.495 55.415 ;
        RECT 15.645 54.505 17.015 55.315 ;
        RECT 17.025 54.505 18.395 55.285 ;
        RECT 18.415 54.590 18.845 55.375 ;
        RECT 18.865 55.185 19.795 55.415 ;
        RECT 24.365 55.185 25.285 55.405 ;
        RECT 31.365 55.305 32.285 55.415 ;
        RECT 29.950 55.185 32.285 55.305 ;
        RECT 34.025 55.185 34.945 55.405 ;
        RECT 41.025 55.305 41.945 55.415 ;
        RECT 39.610 55.185 41.945 55.305 ;
        RECT 18.865 54.505 22.765 55.185 ;
        RECT 23.005 54.505 32.285 55.185 ;
        RECT 32.665 54.505 41.945 55.185 ;
        RECT 42.325 54.505 44.155 55.315 ;
        RECT 44.175 54.590 44.605 55.375 ;
        RECT 44.625 54.505 46.455 55.315 ;
        RECT 46.925 54.505 48.295 55.285 ;
        RECT 48.305 55.185 49.235 55.415 ;
        RECT 52.445 55.185 53.375 55.415 ;
        RECT 48.305 54.505 52.205 55.185 ;
        RECT 52.445 54.505 56.345 55.185 ;
        RECT 56.585 54.505 60.255 55.315 ;
        RECT 60.265 55.185 61.610 55.415 ;
        RECT 60.265 54.505 62.095 55.185 ;
        RECT 62.105 54.505 64.855 55.315 ;
        RECT 64.875 54.505 66.225 55.415 ;
        RECT 66.245 54.505 68.855 55.415 ;
        RECT 69.935 54.590 70.365 55.375 ;
        RECT 74.895 55.185 75.825 55.405 ;
        RECT 78.655 55.185 79.575 55.415 ;
        RECT 70.385 54.505 79.575 55.185 ;
        RECT 79.585 54.505 80.955 55.285 ;
        RECT 84.165 55.185 85.095 55.415 ;
        RECT 81.195 54.505 85.095 55.185 ;
        RECT 85.105 54.505 86.475 55.285 ;
        RECT 86.485 54.505 87.855 55.315 ;
        RECT 87.865 54.505 89.235 55.285 ;
        RECT 89.245 55.185 90.175 55.415 ;
        RECT 89.245 54.505 93.145 55.185 ;
        RECT 93.385 54.505 95.215 55.315 ;
        RECT 95.695 54.590 96.125 55.375 ;
        RECT 97.065 54.505 98.435 55.285 ;
        RECT 98.445 54.505 99.815 55.285 ;
        RECT 101.185 55.185 102.105 55.405 ;
        RECT 108.185 55.305 109.105 55.415 ;
        RECT 106.770 55.185 109.105 55.305 ;
        RECT 99.825 54.505 109.105 55.185 ;
        RECT 109.495 54.505 110.845 55.415 ;
        RECT 110.865 54.505 112.235 55.315 ;
        RECT 112.245 54.505 113.615 55.315 ;
        RECT 5.665 54.295 5.835 54.505 ;
        RECT 7.045 54.295 7.215 54.505 ;
        RECT 8.425 54.295 8.595 54.485 ;
        RECT 10.720 54.345 10.840 54.455 ;
        RECT 12.105 54.315 12.275 54.505 ;
        RECT 12.560 54.345 12.680 54.455 ;
        RECT 13.030 54.315 13.200 54.505 ;
        RECT 15.785 54.315 15.955 54.505 ;
        RECT 17.165 54.315 17.335 54.505 ;
        RECT 17.620 54.345 17.740 54.455 ;
        RECT 18.085 54.295 18.255 54.485 ;
        RECT 19.280 54.315 19.450 54.505 ;
        RECT 23.145 54.315 23.315 54.505 ;
        RECT 28.205 54.295 28.375 54.485 ;
        RECT 29.585 54.295 29.755 54.485 ;
        RECT 30.045 54.295 30.215 54.485 ;
        RECT 32.805 54.295 32.975 54.505 ;
        RECT 33.265 54.295 33.435 54.485 ;
        RECT 35.565 54.295 35.735 54.485 ;
        RECT 36.025 54.295 36.195 54.485 ;
        RECT 37.405 54.295 37.575 54.485 ;
        RECT 38.785 54.295 38.955 54.485 ;
        RECT 42.465 54.315 42.635 54.505 ;
        RECT 43.385 54.295 43.555 54.485 ;
        RECT 44.765 54.295 44.935 54.505 ;
        RECT 46.600 54.345 46.720 54.455 ;
        RECT 47.985 54.315 48.155 54.505 ;
        RECT 48.720 54.315 48.890 54.505 ;
        RECT 52.860 54.315 53.030 54.505 ;
        RECT 56.725 54.295 56.895 54.505 ;
        RECT 57.645 54.295 57.815 54.485 ;
        RECT 59.490 54.295 59.660 54.485 ;
        RECT 61.785 54.315 61.955 54.505 ;
        RECT 62.245 54.295 62.415 54.505 ;
        RECT 65.000 54.345 65.120 54.455 ;
        RECT 65.470 54.295 65.640 54.485 ;
        RECT 65.925 54.315 66.095 54.505 ;
        RECT 66.390 54.315 66.560 54.505 ;
        RECT 68.225 54.295 68.395 54.485 ;
        RECT 69.155 54.350 69.315 54.460 ;
        RECT 70.525 54.315 70.695 54.505 ;
        RECT 70.985 54.295 71.155 54.485 ;
        RECT 80.645 54.315 80.815 54.505 ;
        RECT 81.105 54.295 81.275 54.485 ;
        RECT 81.565 54.295 81.735 54.485 ;
        RECT 83.405 54.295 83.575 54.485 ;
        RECT 84.510 54.315 84.680 54.505 ;
        RECT 86.165 54.315 86.335 54.505 ;
        RECT 86.625 54.315 86.795 54.505 ;
        RECT 88.925 54.315 89.095 54.505 ;
        RECT 89.660 54.315 89.830 54.505 ;
        RECT 93.525 54.295 93.695 54.505 ;
        RECT 95.365 54.455 95.535 54.485 ;
        RECT 93.980 54.345 94.100 54.455 ;
        RECT 95.360 54.345 95.535 54.455 ;
        RECT 95.365 54.295 95.535 54.345 ;
        RECT 95.825 54.295 95.995 54.485 ;
        RECT 96.295 54.350 96.455 54.460 ;
        RECT 97.205 54.315 97.375 54.505 ;
        RECT 98.585 54.455 98.755 54.505 ;
        RECT 98.580 54.345 98.755 54.455 ;
        RECT 98.585 54.315 98.755 54.345 ;
        RECT 99.045 54.295 99.215 54.485 ;
        RECT 99.965 54.315 100.135 54.505 ;
        RECT 109.165 54.295 109.335 54.485 ;
        RECT 109.625 54.315 109.795 54.505 ;
        RECT 111.005 54.315 111.175 54.505 ;
        RECT 111.920 54.345 112.040 54.455 ;
        RECT 113.305 54.295 113.475 54.505 ;
        RECT 5.525 53.485 6.895 54.295 ;
        RECT 6.905 53.485 8.275 54.295 ;
        RECT 8.285 53.615 17.475 54.295 ;
        RECT 17.945 53.615 27.135 54.295 ;
        RECT 12.795 53.395 13.725 53.615 ;
        RECT 16.555 53.385 17.475 53.615 ;
        RECT 22.455 53.395 23.385 53.615 ;
        RECT 26.215 53.385 27.135 53.615 ;
        RECT 27.145 53.515 28.515 54.295 ;
        RECT 28.535 53.385 29.885 54.295 ;
        RECT 29.905 53.485 31.275 54.295 ;
        RECT 31.295 53.425 31.725 54.210 ;
        RECT 31.755 53.385 33.105 54.295 ;
        RECT 33.125 53.485 34.495 54.295 ;
        RECT 34.505 53.515 35.875 54.295 ;
        RECT 35.885 53.485 37.255 54.295 ;
        RECT 37.275 53.385 38.625 54.295 ;
        RECT 38.645 53.485 42.315 54.295 ;
        RECT 43.255 53.385 44.605 54.295 ;
        RECT 44.625 53.615 53.905 54.295 ;
        RECT 54.295 53.615 57.035 54.295 ;
        RECT 45.985 53.395 46.905 53.615 ;
        RECT 51.570 53.495 53.905 53.615 ;
        RECT 52.985 53.385 53.905 53.495 ;
        RECT 57.055 53.425 57.485 54.210 ;
        RECT 57.505 53.485 59.335 54.295 ;
        RECT 59.345 53.385 61.955 54.295 ;
        RECT 62.105 53.615 64.845 54.295 ;
        RECT 65.325 53.385 67.935 54.295 ;
        RECT 68.085 53.485 70.835 54.295 ;
        RECT 70.855 53.385 72.205 54.295 ;
        RECT 72.225 53.615 81.415 54.295 ;
        RECT 72.225 53.385 73.145 53.615 ;
        RECT 75.975 53.395 76.905 53.615 ;
        RECT 81.425 53.485 82.795 54.295 ;
        RECT 82.815 53.425 83.245 54.210 ;
        RECT 83.265 53.615 92.455 54.295 ;
        RECT 87.775 53.395 88.705 53.615 ;
        RECT 91.535 53.385 92.455 53.615 ;
        RECT 92.475 53.385 93.825 54.295 ;
        RECT 94.315 53.385 95.665 54.295 ;
        RECT 95.685 53.485 98.435 54.295 ;
        RECT 98.905 53.615 108.185 54.295 ;
        RECT 100.265 53.395 101.185 53.615 ;
        RECT 105.850 53.495 108.185 53.615 ;
        RECT 107.265 53.385 108.185 53.495 ;
        RECT 108.575 53.425 109.005 54.210 ;
        RECT 109.025 53.485 111.775 54.295 ;
        RECT 112.245 53.485 113.615 54.295 ;
      LAYER nwell ;
        RECT 5.330 50.265 113.810 53.095 ;
      LAYER pwell ;
        RECT 5.525 49.065 6.895 49.875 ;
        RECT 12.865 49.745 13.795 49.975 ;
        RECT 7.825 49.065 9.655 49.745 ;
        RECT 9.895 49.065 13.795 49.745 ;
        RECT 13.805 49.745 14.735 49.975 ;
        RECT 13.805 49.065 17.705 49.745 ;
        RECT 18.415 49.150 18.845 49.935 ;
        RECT 28.525 49.745 29.455 49.975 ;
        RECT 19.410 49.065 28.515 49.745 ;
        RECT 28.525 49.065 32.425 49.745 ;
        RECT 32.665 49.065 35.415 49.875 ;
        RECT 35.425 49.065 36.795 49.845 ;
        RECT 36.805 49.745 37.735 49.975 ;
        RECT 36.805 49.065 40.705 49.745 ;
        RECT 40.945 49.065 42.775 49.875 ;
        RECT 42.785 49.065 44.155 49.845 ;
        RECT 44.175 49.150 44.605 49.935 ;
        RECT 45.985 49.745 46.905 49.965 ;
        RECT 52.985 49.865 53.905 49.975 ;
        RECT 51.570 49.745 53.905 49.865 ;
        RECT 44.625 49.065 53.905 49.745 ;
        RECT 54.285 49.065 57.035 49.875 ;
        RECT 57.535 49.065 60.255 49.975 ;
        RECT 60.265 49.065 61.635 49.875 ;
        RECT 61.655 49.065 64.395 49.745 ;
        RECT 64.405 49.065 69.915 49.875 ;
        RECT 69.935 49.150 70.365 49.935 ;
        RECT 70.385 49.065 75.895 49.875 ;
        RECT 76.835 49.065 78.185 49.975 ;
        RECT 78.205 49.065 81.875 49.875 ;
        RECT 81.885 49.065 83.255 49.875 ;
        RECT 83.460 49.065 86.935 49.975 ;
        RECT 86.945 49.065 92.455 49.875 ;
        RECT 92.465 49.065 95.215 49.875 ;
        RECT 95.695 49.150 96.125 49.935 ;
        RECT 96.145 49.065 99.815 49.875 ;
        RECT 99.825 49.065 101.195 49.875 ;
        RECT 101.205 49.745 102.135 49.975 ;
        RECT 101.205 49.065 105.105 49.745 ;
        RECT 105.345 49.065 110.855 49.875 ;
        RECT 110.865 49.065 112.235 49.875 ;
        RECT 112.245 49.065 113.615 49.875 ;
        RECT 5.665 48.855 5.835 49.065 ;
        RECT 7.045 48.855 7.215 49.045 ;
        RECT 7.965 48.875 8.135 49.065 ;
        RECT 13.210 48.875 13.380 49.065 ;
        RECT 14.220 48.875 14.390 49.065 ;
        RECT 17.165 48.855 17.335 49.045 ;
        RECT 18.085 49.015 18.255 49.045 ;
        RECT 17.620 48.905 17.740 49.015 ;
        RECT 18.080 48.905 18.255 49.015 ;
        RECT 19.000 48.905 19.120 49.015 ;
        RECT 18.085 48.855 18.255 48.905 ;
        RECT 19.470 48.855 19.640 49.045 ;
        RECT 28.205 48.875 28.375 49.065 ;
        RECT 28.940 48.875 29.110 49.065 ;
        RECT 30.515 48.900 30.675 49.010 ;
        RECT 31.885 48.855 32.055 49.045 ;
        RECT 32.805 48.875 32.975 49.065 ;
        RECT 33.265 48.855 33.435 49.045 ;
        RECT 36.485 48.875 36.655 49.065 ;
        RECT 37.220 48.875 37.390 49.065 ;
        RECT 41.085 48.875 41.255 49.065 ;
        RECT 42.925 48.875 43.095 49.065 ;
        RECT 43.385 48.855 43.555 49.045 ;
        RECT 43.845 48.855 44.015 49.045 ;
        RECT 44.765 48.875 44.935 49.065 ;
        RECT 47.535 48.900 47.695 49.010 ;
        RECT 48.445 48.855 48.615 49.045 ;
        RECT 49.825 48.855 49.995 49.045 ;
        RECT 54.425 48.875 54.595 49.065 ;
        RECT 55.345 48.855 55.515 49.045 ;
        RECT 57.180 48.905 57.300 49.015 ;
        RECT 57.645 48.855 57.815 49.045 ;
        RECT 59.945 48.875 60.115 49.065 ;
        RECT 60.405 48.875 60.575 49.065 ;
        RECT 60.865 48.855 61.035 49.045 ;
        RECT 61.325 48.855 61.495 49.045 ;
        RECT 63.165 48.855 63.335 49.045 ;
        RECT 64.085 48.875 64.255 49.065 ;
        RECT 64.545 48.875 64.715 49.065 ;
        RECT 68.685 48.855 68.855 49.045 ;
        RECT 70.525 48.875 70.695 49.065 ;
        RECT 72.360 48.905 72.480 49.015 ;
        RECT 72.825 48.855 72.995 49.045 ;
        RECT 76.055 48.910 76.215 49.020 ;
        RECT 77.885 48.875 78.055 49.065 ;
        RECT 78.345 48.875 78.515 49.065 ;
        RECT 78.800 48.855 78.970 49.045 ;
        RECT 79.265 48.855 79.435 49.045 ;
        RECT 82.025 48.875 82.195 49.065 ;
        RECT 83.405 48.855 83.575 49.045 ;
        RECT 86.165 48.855 86.335 49.045 ;
        RECT 86.620 48.875 86.790 49.065 ;
        RECT 87.085 48.875 87.255 49.065 ;
        RECT 92.605 48.875 92.775 49.065 ;
        RECT 95.370 49.015 95.540 49.045 ;
        RECT 95.360 48.905 95.540 49.015 ;
        RECT 95.370 48.855 95.540 48.905 ;
        RECT 96.285 48.875 96.455 49.065 ;
        RECT 99.965 48.875 100.135 49.065 ;
        RECT 101.620 48.875 101.790 49.065 ;
        RECT 105.485 48.875 105.655 49.065 ;
        RECT 106.405 48.855 106.575 49.045 ;
        RECT 108.240 48.905 108.360 49.015 ;
        RECT 109.165 48.855 109.335 49.045 ;
        RECT 111.005 48.875 111.175 49.065 ;
        RECT 111.920 48.905 112.040 49.015 ;
        RECT 113.305 48.855 113.475 49.065 ;
        RECT 5.525 48.045 6.895 48.855 ;
        RECT 6.905 48.045 8.275 48.855 ;
        RECT 8.285 48.175 17.475 48.855 ;
        RECT 8.285 47.945 9.205 48.175 ;
        RECT 12.035 47.955 12.965 48.175 ;
        RECT 17.945 48.075 19.315 48.855 ;
        RECT 19.325 47.945 30.335 48.855 ;
        RECT 31.295 47.985 31.725 48.770 ;
        RECT 31.745 48.045 33.115 48.855 ;
        RECT 33.125 48.175 42.315 48.855 ;
        RECT 37.635 47.955 38.565 48.175 ;
        RECT 41.395 47.945 42.315 48.175 ;
        RECT 42.335 47.945 43.685 48.855 ;
        RECT 43.705 48.045 47.375 48.855 ;
        RECT 48.315 47.945 49.665 48.855 ;
        RECT 49.685 48.045 55.195 48.855 ;
        RECT 55.205 48.045 57.035 48.855 ;
        RECT 57.055 47.985 57.485 48.770 ;
        RECT 57.505 48.045 59.335 48.855 ;
        RECT 59.345 48.175 61.175 48.855 ;
        RECT 61.185 48.175 63.015 48.855 ;
        RECT 59.345 47.945 60.690 48.175 ;
        RECT 61.670 47.945 63.015 48.175 ;
        RECT 63.025 48.045 68.535 48.855 ;
        RECT 68.545 48.045 72.215 48.855 ;
        RECT 72.685 48.045 74.775 48.855 ;
        RECT 75.640 47.945 79.115 48.855 ;
        RECT 79.125 48.045 82.795 48.855 ;
        RECT 82.815 47.985 83.245 48.770 ;
        RECT 83.265 48.045 86.015 48.855 ;
        RECT 86.025 48.175 95.215 48.855 ;
        RECT 90.535 47.955 91.465 48.175 ;
        RECT 94.295 47.945 95.215 48.175 ;
        RECT 95.225 47.945 106.235 48.855 ;
        RECT 106.265 48.045 108.095 48.855 ;
        RECT 108.575 47.985 109.005 48.770 ;
        RECT 109.025 48.045 111.775 48.855 ;
        RECT 112.245 48.045 113.615 48.855 ;
      LAYER nwell ;
        RECT 5.330 44.825 113.810 47.655 ;
      LAYER pwell ;
        RECT 5.525 43.625 6.895 44.435 ;
        RECT 6.905 43.625 12.415 44.435 ;
        RECT 12.425 43.625 16.095 44.435 ;
        RECT 17.035 43.625 18.385 44.535 ;
        RECT 18.415 43.710 18.845 44.495 ;
        RECT 18.875 43.625 20.225 44.535 ;
        RECT 20.245 43.625 21.615 44.405 ;
        RECT 26.135 44.305 27.065 44.525 ;
        RECT 29.895 44.305 30.815 44.535 ;
        RECT 21.625 43.625 30.815 44.305 ;
        RECT 30.835 43.625 32.185 44.535 ;
        RECT 32.205 43.625 37.715 44.435 ;
        RECT 38.600 43.625 39.555 44.305 ;
        RECT 39.565 43.625 43.235 44.435 ;
        RECT 44.175 43.710 44.605 44.495 ;
        RECT 44.765 43.625 47.375 44.535 ;
        RECT 48.040 43.625 51.515 44.535 ;
        RECT 51.525 43.625 55.195 44.435 ;
        RECT 55.205 43.625 56.575 44.435 ;
        RECT 56.585 44.305 57.930 44.535 ;
        RECT 58.910 44.305 60.255 44.535 ;
        RECT 56.585 43.625 58.415 44.305 ;
        RECT 58.425 43.625 60.255 44.305 ;
        RECT 60.265 44.305 61.610 44.535 ;
        RECT 62.590 44.305 63.935 44.535 ;
        RECT 64.430 44.305 65.775 44.535 ;
        RECT 60.265 43.625 62.095 44.305 ;
        RECT 62.105 43.625 63.935 44.305 ;
        RECT 63.945 43.625 65.775 44.305 ;
        RECT 65.785 43.625 69.455 44.435 ;
        RECT 69.935 43.710 70.365 44.495 ;
        RECT 70.385 43.625 72.215 44.435 ;
        RECT 72.685 43.625 81.790 44.305 ;
        RECT 81.885 43.625 85.360 44.535 ;
        RECT 85.565 43.625 89.040 44.535 ;
        RECT 89.245 43.625 92.720 44.535 ;
        RECT 92.925 43.625 95.675 44.435 ;
        RECT 95.695 43.710 96.125 44.495 ;
        RECT 96.145 43.625 105.250 44.305 ;
        RECT 105.345 43.625 110.855 44.435 ;
        RECT 110.865 43.625 112.235 44.435 ;
        RECT 112.245 43.625 113.615 44.435 ;
        RECT 5.665 43.415 5.835 43.625 ;
        RECT 7.045 43.415 7.215 43.625 ;
        RECT 12.565 43.415 12.735 43.625 ;
        RECT 16.255 43.460 16.415 43.580 ;
        RECT 18.085 43.435 18.255 43.625 ;
        RECT 19.925 43.435 20.095 43.625 ;
        RECT 20.380 43.415 20.550 43.605 ;
        RECT 21.305 43.435 21.475 43.625 ;
        RECT 21.765 43.435 21.935 43.625 ;
        RECT 31.885 43.605 32.055 43.625 ;
        RECT 24.060 43.415 24.230 43.605 ;
        RECT 24.525 43.415 24.695 43.605 ;
        RECT 29.580 43.415 29.750 43.605 ;
        RECT 30.045 43.415 30.215 43.605 ;
        RECT 31.885 43.435 32.060 43.605 ;
        RECT 32.345 43.435 32.515 43.625 ;
        RECT 31.890 43.415 32.060 43.435 ;
        RECT 35.565 43.415 35.735 43.605 ;
        RECT 36.945 43.415 37.115 43.605 ;
        RECT 37.860 43.465 37.980 43.575 ;
        RECT 38.325 43.435 38.495 43.605 ;
        RECT 39.705 43.435 39.875 43.625 ;
        RECT 47.060 43.605 47.230 43.625 ;
        RECT 43.395 43.470 43.555 43.580 ;
        RECT 47.060 43.435 47.235 43.605 ;
        RECT 47.520 43.570 47.640 43.575 ;
        RECT 47.520 43.465 47.695 43.570 ;
        RECT 47.535 43.460 47.695 43.465 ;
        RECT 51.200 43.435 51.370 43.625 ;
        RECT 51.665 43.605 51.835 43.625 ;
        RECT 55.345 43.605 55.515 43.625 ;
        RECT 51.660 43.435 51.835 43.605 ;
        RECT 55.340 43.435 55.515 43.605 ;
        RECT 47.065 43.415 47.235 43.435 ;
        RECT 51.660 43.415 51.830 43.435 ;
        RECT 55.340 43.415 55.510 43.435 ;
        RECT 55.805 43.415 55.975 43.605 ;
        RECT 58.105 43.435 58.275 43.625 ;
        RECT 58.565 43.435 58.735 43.625 ;
        RECT 59.945 43.415 60.115 43.605 ;
        RECT 60.405 43.415 60.575 43.605 ;
        RECT 61.785 43.415 61.955 43.625 ;
        RECT 62.245 43.435 62.415 43.625 ;
        RECT 64.085 43.435 64.255 43.625 ;
        RECT 64.540 43.465 64.660 43.575 ;
        RECT 65.005 43.415 65.175 43.605 ;
        RECT 65.925 43.435 66.095 43.625 ;
        RECT 69.600 43.465 69.720 43.575 ;
        RECT 70.525 43.435 70.695 43.625 ;
        RECT 72.360 43.465 72.480 43.575 ;
        RECT 72.825 43.435 72.995 43.625 ;
        RECT 74.480 43.415 74.650 43.605 ;
        RECT 78.350 43.415 78.520 43.605 ;
        RECT 82.030 43.435 82.200 43.625 ;
        RECT 83.405 43.415 83.575 43.605 ;
        RECT 85.710 43.435 85.880 43.625 ;
        RECT 89.390 43.435 89.560 43.625 ;
        RECT 92.610 43.415 92.780 43.605 ;
        RECT 93.065 43.435 93.235 43.625 ;
        RECT 96.285 43.415 96.455 43.625 ;
        RECT 105.485 43.415 105.655 43.625 ;
        RECT 106.865 43.415 107.035 43.605 ;
        RECT 109.165 43.415 109.335 43.605 ;
        RECT 111.005 43.435 111.175 43.625 ;
        RECT 111.920 43.465 112.040 43.575 ;
        RECT 113.305 43.415 113.475 43.625 ;
        RECT 5.525 42.605 6.895 43.415 ;
        RECT 6.905 42.605 12.415 43.415 ;
        RECT 12.425 42.605 16.095 43.415 ;
        RECT 17.220 42.505 20.695 43.415 ;
        RECT 20.900 42.505 24.375 43.415 ;
        RECT 24.385 42.605 26.215 43.415 ;
        RECT 26.420 42.505 29.895 43.415 ;
        RECT 29.905 42.605 31.275 43.415 ;
        RECT 31.295 42.545 31.725 43.330 ;
        RECT 31.745 42.505 35.220 43.415 ;
        RECT 35.435 42.505 36.785 43.415 ;
        RECT 36.805 42.605 38.175 43.415 ;
        RECT 38.270 42.735 47.375 43.415 ;
        RECT 48.500 42.505 51.975 43.415 ;
        RECT 52.180 42.505 55.655 43.415 ;
        RECT 55.665 42.605 57.035 43.415 ;
        RECT 57.055 42.545 57.485 43.330 ;
        RECT 57.535 42.505 60.255 43.415 ;
        RECT 60.265 42.605 61.635 43.415 ;
        RECT 61.645 42.735 64.385 43.415 ;
        RECT 64.865 42.735 74.055 43.415 ;
        RECT 69.375 42.515 70.305 42.735 ;
        RECT 73.135 42.505 74.055 42.735 ;
        RECT 74.065 42.735 77.965 43.415 ;
        RECT 74.065 42.505 74.995 42.735 ;
        RECT 78.205 42.505 81.680 43.415 ;
        RECT 82.815 42.545 83.245 43.330 ;
        RECT 83.265 42.735 92.455 43.415 ;
        RECT 87.775 42.515 88.705 42.735 ;
        RECT 91.535 42.505 92.455 42.735 ;
        RECT 92.465 42.505 95.940 43.415 ;
        RECT 96.145 42.735 105.335 43.415 ;
        RECT 100.655 42.515 101.585 42.735 ;
        RECT 104.415 42.505 105.335 42.735 ;
        RECT 105.355 42.505 106.705 43.415 ;
        RECT 106.725 42.605 108.555 43.415 ;
        RECT 108.575 42.545 109.005 43.330 ;
        RECT 109.025 42.605 111.775 43.415 ;
        RECT 112.245 42.605 113.615 43.415 ;
      LAYER nwell ;
        RECT 5.330 39.385 113.810 42.215 ;
      LAYER pwell ;
        RECT 5.525 38.185 6.895 38.995 ;
        RECT 6.905 38.185 10.575 38.995 ;
        RECT 11.505 38.185 12.875 38.965 ;
        RECT 12.885 38.185 14.255 38.965 ;
        RECT 14.275 38.185 15.625 39.095 ;
        RECT 15.655 38.185 17.005 39.095 ;
        RECT 17.025 38.185 18.395 38.995 ;
        RECT 18.415 38.270 18.845 39.055 ;
        RECT 18.865 38.185 22.535 38.995 ;
        RECT 22.740 38.185 26.215 39.095 ;
        RECT 26.225 38.185 29.700 39.095 ;
        RECT 34.875 38.865 35.805 39.085 ;
        RECT 38.635 38.865 39.555 39.095 ;
        RECT 30.365 38.185 39.555 38.865 ;
        RECT 40.485 38.185 41.855 38.965 ;
        RECT 41.865 38.185 43.695 38.995 ;
        RECT 44.175 38.270 44.605 39.055 ;
        RECT 44.625 38.865 45.555 39.095 ;
        RECT 44.625 38.185 48.525 38.865 ;
        RECT 48.960 38.185 52.435 39.095 ;
        RECT 52.455 38.185 55.195 38.865 ;
        RECT 55.205 38.185 57.955 38.995 ;
        RECT 58.180 38.415 60.935 39.095 ;
        RECT 58.665 38.185 60.935 38.415 ;
        RECT 62.245 38.185 64.855 39.095 ;
        RECT 64.875 38.185 66.225 39.095 ;
        RECT 66.245 38.185 67.615 38.965 ;
        RECT 67.625 38.185 68.995 38.965 ;
        RECT 69.935 38.270 70.365 39.055 ;
        RECT 70.395 38.185 71.745 39.095 ;
        RECT 72.225 38.865 73.155 39.095 ;
        RECT 72.225 38.185 76.125 38.865 ;
        RECT 76.365 38.185 78.195 38.995 ;
        RECT 78.400 38.185 81.875 39.095 ;
        RECT 85.545 38.865 86.475 39.095 ;
        RECT 82.575 38.185 86.475 38.865 ;
        RECT 86.485 38.185 87.855 38.965 ;
        RECT 88.060 38.185 91.535 39.095 ;
        RECT 94.745 38.865 95.675 39.095 ;
        RECT 91.775 38.185 95.675 38.865 ;
        RECT 95.695 38.270 96.125 39.055 ;
        RECT 96.605 38.865 97.525 39.095 ;
        RECT 100.355 38.865 101.285 39.085 ;
        RECT 96.605 38.185 105.795 38.865 ;
        RECT 105.805 38.185 111.315 38.995 ;
        RECT 112.245 38.185 113.615 38.995 ;
        RECT 5.665 37.975 5.835 38.185 ;
        RECT 7.045 37.975 7.215 38.185 ;
        RECT 8.425 37.975 8.595 38.165 ;
        RECT 10.735 38.030 10.895 38.140 ;
        RECT 12.565 37.995 12.735 38.185 ;
        RECT 13.945 37.995 14.115 38.185 ;
        RECT 15.325 37.995 15.495 38.185 ;
        RECT 16.705 37.995 16.875 38.185 ;
        RECT 17.165 37.995 17.335 38.185 ;
        RECT 17.900 37.975 18.070 38.165 ;
        RECT 19.005 37.995 19.175 38.185 ;
        RECT 21.765 37.975 21.935 38.165 ;
        RECT 24.800 37.975 24.970 38.165 ;
        RECT 25.900 37.995 26.070 38.185 ;
        RECT 26.370 37.995 26.540 38.185 ;
        RECT 28.660 38.025 28.780 38.135 ;
        RECT 29.125 37.975 29.295 38.165 ;
        RECT 30.040 38.025 30.160 38.135 ;
        RECT 30.505 37.995 30.675 38.185 ;
        RECT 32.160 37.975 32.330 38.165 ;
        RECT 36.025 37.975 36.195 38.165 ;
        RECT 37.860 38.025 37.980 38.135 ;
        RECT 38.325 37.975 38.495 38.165 ;
        RECT 39.715 38.030 39.875 38.140 ;
        RECT 41.545 37.995 41.715 38.185 ;
        RECT 42.005 37.995 42.175 38.185 ;
        RECT 43.840 38.025 43.960 38.135 ;
        RECT 45.040 37.995 45.210 38.185 ;
        RECT 47.525 37.975 47.695 38.165 ;
        RECT 48.905 37.975 49.075 38.165 ;
        RECT 52.120 37.995 52.290 38.185 ;
        RECT 54.425 37.975 54.595 38.165 ;
        RECT 54.885 37.995 55.055 38.185 ;
        RECT 55.345 37.995 55.515 38.185 ;
        RECT 60.865 38.165 60.935 38.185 ;
        RECT 57.655 38.020 57.815 38.130 ;
        RECT 58.565 37.975 58.735 38.165 ;
        RECT 60.865 37.995 61.035 38.165 ;
        RECT 61.335 38.030 61.495 38.140 ;
        RECT 64.085 37.975 64.255 38.165 ;
        RECT 64.540 37.995 64.710 38.185 ;
        RECT 65.925 37.995 66.095 38.185 ;
        RECT 66.385 37.995 66.555 38.185 ;
        RECT 67.765 37.975 67.935 38.165 ;
        RECT 68.685 37.995 68.855 38.185 ;
        RECT 69.145 37.975 69.315 38.165 ;
        RECT 71.445 37.995 71.615 38.185 ;
        RECT 71.900 38.025 72.020 38.135 ;
        RECT 72.640 37.995 72.810 38.185 ;
        RECT 76.505 37.995 76.675 38.185 ;
        RECT 79.265 37.975 79.435 38.165 ;
        RECT 79.725 37.975 79.895 38.165 ;
        RECT 81.560 37.995 81.730 38.185 ;
        RECT 82.020 38.025 82.140 38.135 ;
        RECT 82.480 38.025 82.600 38.135 ;
        RECT 83.405 37.975 83.575 38.165 ;
        RECT 85.890 37.995 86.060 38.185 ;
        RECT 87.095 38.020 87.255 38.130 ;
        RECT 87.545 37.995 87.715 38.185 ;
        RECT 88.005 37.975 88.175 38.165 ;
        RECT 89.395 38.020 89.555 38.130 ;
        RECT 91.220 37.995 91.390 38.185 ;
        RECT 93.520 37.975 93.690 38.165 ;
        RECT 93.985 37.975 94.155 38.165 ;
        RECT 95.090 37.995 95.260 38.185 ;
        RECT 95.365 37.975 95.535 38.165 ;
        RECT 96.280 38.025 96.400 38.135 ;
        RECT 100.150 37.975 100.320 38.165 ;
        RECT 100.885 37.975 101.055 38.165 ;
        RECT 103.185 37.975 103.355 38.165 ;
        RECT 103.645 37.975 103.815 38.165 ;
        RECT 105.485 37.995 105.655 38.185 ;
        RECT 105.945 37.995 106.115 38.185 ;
        RECT 107.325 37.975 107.495 38.165 ;
        RECT 109.165 37.975 109.335 38.165 ;
        RECT 111.475 38.030 111.635 38.140 ;
        RECT 111.920 38.025 112.040 38.135 ;
        RECT 113.305 37.975 113.475 38.185 ;
        RECT 5.525 37.165 6.895 37.975 ;
        RECT 6.905 37.165 8.275 37.975 ;
        RECT 8.285 37.295 17.475 37.975 ;
        RECT 12.795 37.075 13.725 37.295 ;
        RECT 16.555 37.065 17.475 37.295 ;
        RECT 17.485 37.295 21.385 37.975 ;
        RECT 17.485 37.065 18.415 37.295 ;
        RECT 21.625 37.165 24.375 37.975 ;
        RECT 24.385 37.295 28.285 37.975 ;
        RECT 24.385 37.065 25.315 37.295 ;
        RECT 28.985 37.195 30.355 37.975 ;
        RECT 31.295 37.105 31.725 37.890 ;
        RECT 31.745 37.295 35.645 37.975 ;
        RECT 31.745 37.065 32.675 37.295 ;
        RECT 35.885 37.165 37.715 37.975 ;
        RECT 38.185 37.295 47.375 37.975 ;
        RECT 42.695 37.075 43.625 37.295 ;
        RECT 46.455 37.065 47.375 37.295 ;
        RECT 47.395 37.065 48.745 37.975 ;
        RECT 48.765 37.165 54.275 37.975 ;
        RECT 54.285 37.165 57.035 37.975 ;
        RECT 57.055 37.105 57.485 37.890 ;
        RECT 58.425 37.745 62.850 37.975 ;
        RECT 58.425 37.065 63.790 37.745 ;
        RECT 63.945 37.165 67.615 37.975 ;
        RECT 67.625 37.165 68.995 37.975 ;
        RECT 69.005 37.295 78.195 37.975 ;
        RECT 73.515 37.075 74.445 37.295 ;
        RECT 77.275 37.065 78.195 37.295 ;
        RECT 78.215 37.065 79.565 37.975 ;
        RECT 79.585 37.165 82.335 37.975 ;
        RECT 82.815 37.105 83.245 37.890 ;
        RECT 83.265 37.165 86.935 37.975 ;
        RECT 87.875 37.065 89.225 37.975 ;
        RECT 90.360 37.065 93.835 37.975 ;
        RECT 93.845 37.195 95.215 37.975 ;
        RECT 95.225 37.165 96.595 37.975 ;
        RECT 96.835 37.295 100.735 37.975 ;
        RECT 99.805 37.065 100.735 37.295 ;
        RECT 100.745 37.195 102.115 37.975 ;
        RECT 102.135 37.065 103.485 37.975 ;
        RECT 103.505 37.165 107.175 37.975 ;
        RECT 107.185 37.165 108.555 37.975 ;
        RECT 108.575 37.105 109.005 37.890 ;
        RECT 109.025 37.165 111.775 37.975 ;
        RECT 112.245 37.165 113.615 37.975 ;
      LAYER nwell ;
        RECT 5.330 33.945 113.810 36.775 ;
      LAYER pwell ;
        RECT 5.525 32.745 6.895 33.555 ;
        RECT 6.905 32.745 8.735 33.555 ;
        RECT 13.255 33.425 14.185 33.645 ;
        RECT 17.015 33.425 17.935 33.655 ;
        RECT 8.745 32.745 17.935 33.425 ;
        RECT 18.415 32.830 18.845 33.615 ;
        RECT 18.865 33.425 19.795 33.655 ;
        RECT 28.435 33.425 29.365 33.645 ;
        RECT 32.195 33.425 33.115 33.655 ;
        RECT 18.865 32.745 22.765 33.425 ;
        RECT 23.925 32.745 33.115 33.425 ;
        RECT 33.135 32.745 34.485 33.655 ;
        RECT 34.505 32.745 40.015 33.555 ;
        RECT 40.025 32.745 41.395 33.555 ;
        RECT 41.405 32.745 42.775 33.525 ;
        RECT 42.785 32.745 44.155 33.555 ;
        RECT 44.175 32.830 44.605 33.615 ;
        RECT 44.625 33.425 45.555 33.655 ;
        RECT 44.625 32.745 48.525 33.425 ;
        RECT 48.765 32.745 54.275 33.555 ;
        RECT 54.285 32.745 57.035 33.555 ;
        RECT 57.055 33.425 60.055 33.655 ;
        RECT 57.055 33.335 61.635 33.425 ;
        RECT 57.045 32.975 61.635 33.335 ;
        RECT 57.045 32.785 57.975 32.975 ;
        RECT 57.055 32.745 57.975 32.785 ;
        RECT 60.065 32.745 61.635 32.975 ;
        RECT 61.885 32.975 64.640 33.655 ;
        RECT 61.885 32.745 64.155 32.975 ;
        RECT 64.865 32.745 68.535 33.555 ;
        RECT 68.545 32.745 69.915 33.555 ;
        RECT 69.935 32.830 70.365 33.615 ;
        RECT 70.385 32.745 75.895 33.555 ;
        RECT 79.565 33.425 80.495 33.655 ;
        RECT 76.595 32.745 80.495 33.425 ;
        RECT 80.515 32.745 81.865 33.655 ;
        RECT 81.885 32.745 87.395 33.555 ;
        RECT 87.405 32.745 88.775 33.555 ;
        RECT 88.785 33.425 89.715 33.655 ;
        RECT 88.785 32.745 92.685 33.425 ;
        RECT 93.385 32.745 94.755 33.525 ;
        RECT 95.695 32.830 96.125 33.615 ;
        RECT 96.145 33.425 97.075 33.655 ;
        RECT 96.145 32.745 100.045 33.425 ;
        RECT 100.285 32.745 105.795 33.555 ;
        RECT 105.805 32.745 111.315 33.555 ;
        RECT 112.245 32.745 113.615 33.555 ;
        RECT 5.665 32.535 5.835 32.745 ;
        RECT 7.045 32.535 7.215 32.745 ;
        RECT 8.885 32.555 9.055 32.745 ;
        RECT 12.565 32.535 12.735 32.725 ;
        RECT 16.245 32.535 16.415 32.725 ;
        RECT 18.080 32.585 18.200 32.695 ;
        RECT 19.280 32.555 19.450 32.745 ;
        RECT 21.030 32.535 21.200 32.725 ;
        RECT 21.765 32.535 21.935 32.725 ;
        RECT 23.155 32.590 23.315 32.700 ;
        RECT 24.065 32.555 24.235 32.745 ;
        RECT 24.525 32.535 24.695 32.725 ;
        RECT 25.905 32.535 26.075 32.725 ;
        RECT 31.885 32.535 32.055 32.725 ;
        RECT 34.185 32.555 34.355 32.745 ;
        RECT 34.645 32.555 34.815 32.745 ;
        RECT 37.405 32.535 37.575 32.725 ;
        RECT 39.245 32.535 39.415 32.725 ;
        RECT 40.165 32.555 40.335 32.745 ;
        RECT 42.465 32.555 42.635 32.745 ;
        RECT 42.925 32.555 43.095 32.745 ;
        RECT 45.040 32.555 45.210 32.745 ;
        RECT 48.905 32.555 49.075 32.745 ;
        RECT 49.180 32.535 49.350 32.725 ;
        RECT 53.045 32.535 53.215 32.725 ;
        RECT 54.425 32.535 54.595 32.745 ;
        RECT 60.405 32.555 60.575 32.725 ;
        RECT 60.405 32.535 60.475 32.555 ;
        RECT 60.865 32.535 61.035 32.725 ;
        RECT 61.325 32.555 61.495 32.745 ;
        RECT 61.885 32.725 61.955 32.745 ;
        RECT 61.785 32.555 61.955 32.725 ;
        RECT 65.005 32.555 65.175 32.745 ;
        RECT 66.385 32.535 66.555 32.725 ;
        RECT 68.685 32.555 68.855 32.745 ;
        RECT 69.140 32.585 69.260 32.695 ;
        RECT 69.880 32.535 70.050 32.725 ;
        RECT 70.525 32.555 70.695 32.745 ;
        RECT 73.745 32.535 73.915 32.725 ;
        RECT 76.040 32.585 76.160 32.695 ;
        RECT 79.910 32.555 80.080 32.745 ;
        RECT 80.645 32.555 80.815 32.745 ;
        RECT 82.025 32.555 82.195 32.745 ;
        RECT 83.415 32.580 83.575 32.690 ;
        RECT 84.600 32.535 84.770 32.725 ;
        RECT 87.545 32.555 87.715 32.745 ;
        RECT 89.200 32.555 89.370 32.745 ;
        RECT 89.385 32.535 89.555 32.725 ;
        RECT 89.855 32.580 90.015 32.690 ;
        RECT 90.765 32.535 90.935 32.725 ;
        RECT 92.145 32.535 92.315 32.725 ;
        RECT 93.060 32.585 93.180 32.695 ;
        RECT 94.445 32.555 94.615 32.745 ;
        RECT 94.915 32.590 95.075 32.700 ;
        RECT 96.560 32.555 96.730 32.745 ;
        RECT 100.425 32.555 100.595 32.745 ;
        RECT 102.265 32.535 102.435 32.725 ;
        RECT 102.725 32.535 102.895 32.725 ;
        RECT 105.945 32.555 106.115 32.745 ;
        RECT 108.240 32.585 108.360 32.695 ;
        RECT 109.165 32.535 109.335 32.725 ;
        RECT 111.475 32.590 111.635 32.700 ;
        RECT 111.920 32.585 112.040 32.695 ;
        RECT 113.305 32.535 113.475 32.745 ;
        RECT 5.525 31.725 6.895 32.535 ;
        RECT 6.905 31.725 12.415 32.535 ;
        RECT 12.425 31.725 16.095 32.535 ;
        RECT 16.105 31.725 17.475 32.535 ;
        RECT 17.715 31.855 21.615 32.535 ;
        RECT 20.685 31.625 21.615 31.855 ;
        RECT 21.625 31.725 24.375 32.535 ;
        RECT 24.385 31.755 25.755 32.535 ;
        RECT 25.765 31.725 31.275 32.535 ;
        RECT 31.295 31.665 31.725 32.450 ;
        RECT 31.745 31.725 37.255 32.535 ;
        RECT 37.265 31.725 39.095 32.535 ;
        RECT 39.105 31.855 48.385 32.535 ;
        RECT 40.465 31.635 41.385 31.855 ;
        RECT 46.050 31.735 48.385 31.855 ;
        RECT 47.465 31.625 48.385 31.735 ;
        RECT 48.765 31.855 52.665 32.535 ;
        RECT 48.765 31.625 49.695 31.855 ;
        RECT 52.915 31.625 54.265 32.535 ;
        RECT 54.285 31.725 57.035 32.535 ;
        RECT 57.055 31.665 57.485 32.450 ;
        RECT 58.205 32.305 60.475 32.535 ;
        RECT 57.720 31.625 60.475 32.305 ;
        RECT 60.725 31.725 66.235 32.535 ;
        RECT 66.245 31.725 68.995 32.535 ;
        RECT 69.465 31.855 73.365 32.535 ;
        RECT 73.605 31.855 82.795 32.535 ;
        RECT 69.465 31.625 70.395 31.855 ;
        RECT 78.115 31.635 79.045 31.855 ;
        RECT 81.875 31.625 82.795 31.855 ;
        RECT 82.815 31.665 83.245 32.450 ;
        RECT 84.185 31.855 88.085 32.535 ;
        RECT 84.185 31.625 85.115 31.855 ;
        RECT 88.325 31.755 89.695 32.535 ;
        RECT 90.635 31.625 91.985 32.535 ;
        RECT 92.005 31.855 101.195 32.535 ;
        RECT 96.515 31.635 97.445 31.855 ;
        RECT 100.275 31.625 101.195 31.855 ;
        RECT 101.215 31.625 102.565 32.535 ;
        RECT 102.585 31.725 108.095 32.535 ;
        RECT 108.575 31.665 109.005 32.450 ;
        RECT 109.025 31.725 111.775 32.535 ;
        RECT 112.245 31.725 113.615 32.535 ;
      LAYER nwell ;
        RECT 5.330 28.505 113.810 31.335 ;
      LAYER pwell ;
        RECT 5.525 27.305 6.895 28.115 ;
        RECT 6.905 27.305 8.735 28.115 ;
        RECT 13.715 27.985 14.645 28.205 ;
        RECT 17.475 27.985 18.395 28.215 ;
        RECT 9.205 27.305 18.395 27.985 ;
        RECT 18.415 27.390 18.845 28.175 ;
        RECT 18.865 27.305 20.235 28.085 ;
        RECT 20.245 27.305 22.075 28.115 ;
        RECT 22.545 27.985 23.475 28.215 ;
        RECT 22.545 27.305 26.445 27.985 ;
        RECT 26.685 27.305 30.355 28.115 ;
        RECT 30.365 27.985 31.295 28.215 ;
        RECT 34.875 28.105 35.795 28.215 ;
        RECT 34.875 27.985 37.210 28.105 ;
        RECT 41.875 27.985 42.795 28.205 ;
        RECT 30.365 27.305 34.265 27.985 ;
        RECT 34.875 27.305 44.155 27.985 ;
        RECT 44.175 27.390 44.605 28.175 ;
        RECT 44.635 27.305 45.985 28.215 ;
        RECT 46.015 27.305 47.365 28.215 ;
        RECT 52.355 27.985 53.285 28.205 ;
        RECT 56.115 27.985 57.035 28.215 ;
        RECT 58.625 27.985 61.625 28.215 ;
        RECT 47.845 27.305 57.035 27.985 ;
        RECT 57.045 27.895 61.625 27.985 ;
        RECT 57.045 27.535 61.635 27.895 ;
        RECT 57.045 27.305 58.615 27.535 ;
        RECT 60.705 27.345 61.635 27.535 ;
        RECT 60.705 27.305 61.625 27.345 ;
        RECT 61.645 27.305 67.155 28.115 ;
        RECT 67.165 27.305 68.535 28.115 ;
        RECT 68.545 27.305 69.915 28.085 ;
        RECT 69.935 27.390 70.365 28.175 ;
        RECT 74.895 27.985 75.825 28.205 ;
        RECT 78.655 27.985 79.575 28.215 ;
        RECT 70.385 27.305 79.575 27.985 ;
        RECT 79.585 27.305 80.955 28.085 ;
        RECT 80.975 27.305 82.325 28.215 ;
        RECT 82.345 27.305 83.715 28.085 ;
        RECT 83.725 27.305 85.555 28.115 ;
        RECT 87.385 27.985 88.305 28.205 ;
        RECT 94.385 28.105 95.305 28.215 ;
        RECT 92.970 27.985 95.305 28.105 ;
        RECT 86.025 27.305 95.305 27.985 ;
        RECT 95.695 27.390 96.125 28.175 ;
        RECT 96.145 27.305 101.655 28.115 ;
        RECT 101.665 27.305 107.175 28.115 ;
        RECT 107.185 27.305 110.855 28.115 ;
        RECT 110.865 27.305 112.235 28.115 ;
        RECT 112.245 27.305 113.615 28.115 ;
        RECT 5.665 27.095 5.835 27.305 ;
        RECT 7.045 27.095 7.215 27.305 ;
        RECT 8.880 27.145 9.000 27.255 ;
        RECT 9.345 27.115 9.515 27.305 ;
        RECT 12.565 27.095 12.735 27.285 ;
        RECT 16.240 27.145 16.360 27.255 ;
        RECT 17.625 27.095 17.795 27.285 ;
        RECT 18.085 27.095 18.255 27.285 ;
        RECT 19.925 27.115 20.095 27.305 ;
        RECT 20.385 27.115 20.555 27.305 ;
        RECT 22.220 27.145 22.340 27.255 ;
        RECT 22.960 27.115 23.130 27.305 ;
        RECT 26.825 27.115 26.995 27.305 ;
        RECT 28.205 27.095 28.375 27.285 ;
        RECT 28.665 27.095 28.835 27.285 ;
        RECT 30.045 27.095 30.215 27.285 ;
        RECT 30.780 27.115 30.950 27.305 ;
        RECT 40.625 27.095 40.795 27.285 ;
        RECT 42.005 27.095 42.175 27.285 ;
        RECT 42.465 27.095 42.635 27.285 ;
        RECT 43.845 27.115 44.015 27.305 ;
        RECT 45.685 27.115 45.855 27.305 ;
        RECT 47.065 27.115 47.235 27.305 ;
        RECT 47.520 27.145 47.640 27.255 ;
        RECT 47.985 27.095 48.155 27.305 ;
        RECT 54.425 27.095 54.595 27.285 ;
        RECT 54.885 27.095 55.055 27.285 ;
        RECT 56.720 27.145 56.840 27.255 ;
        RECT 57.185 27.115 57.355 27.305 ;
        RECT 57.645 27.095 57.815 27.285 ;
        RECT 61.325 27.095 61.495 27.285 ;
        RECT 61.785 27.115 61.955 27.305 ;
        RECT 63.165 27.095 63.335 27.285 ;
        RECT 67.305 27.115 67.475 27.305 ;
        RECT 68.685 27.095 68.855 27.305 ;
        RECT 70.525 27.115 70.695 27.305 ;
        RECT 72.360 27.145 72.480 27.255 ;
        RECT 72.825 27.095 72.995 27.285 ;
        RECT 74.205 27.095 74.375 27.285 ;
        RECT 79.725 27.095 79.895 27.285 ;
        RECT 80.645 27.115 80.815 27.305 ;
        RECT 81.105 27.115 81.275 27.305 ;
        RECT 82.485 27.255 82.655 27.305 ;
        RECT 82.480 27.145 82.655 27.255 ;
        RECT 82.485 27.115 82.655 27.145 ;
        RECT 83.405 27.095 83.575 27.285 ;
        RECT 83.865 27.115 84.035 27.305 ;
        RECT 85.700 27.145 85.820 27.255 ;
        RECT 86.165 27.115 86.335 27.305 ;
        RECT 88.925 27.095 89.095 27.285 ;
        RECT 94.445 27.095 94.615 27.285 ;
        RECT 96.285 27.115 96.455 27.305 ;
        RECT 99.965 27.095 100.135 27.285 ;
        RECT 101.805 27.115 101.975 27.305 ;
        RECT 105.485 27.095 105.655 27.285 ;
        RECT 107.325 27.115 107.495 27.305 ;
        RECT 108.240 27.145 108.360 27.255 ;
        RECT 109.165 27.095 109.335 27.285 ;
        RECT 111.005 27.115 111.175 27.305 ;
        RECT 111.920 27.145 112.040 27.255 ;
        RECT 113.305 27.095 113.475 27.305 ;
        RECT 5.525 26.285 6.895 27.095 ;
        RECT 6.905 26.285 12.415 27.095 ;
        RECT 12.425 26.285 16.095 27.095 ;
        RECT 16.575 26.185 17.925 27.095 ;
        RECT 17.945 26.415 27.135 27.095 ;
        RECT 22.455 26.195 23.385 26.415 ;
        RECT 26.215 26.185 27.135 26.415 ;
        RECT 27.155 26.185 28.505 27.095 ;
        RECT 28.525 26.285 29.895 27.095 ;
        RECT 29.905 26.315 31.275 27.095 ;
        RECT 31.295 26.225 31.725 27.010 ;
        RECT 31.745 26.415 40.935 27.095 ;
        RECT 31.745 26.185 32.665 26.415 ;
        RECT 35.495 26.195 36.425 26.415 ;
        RECT 40.945 26.315 42.315 27.095 ;
        RECT 42.325 26.285 47.835 27.095 ;
        RECT 47.845 26.285 53.355 27.095 ;
        RECT 53.375 26.185 54.725 27.095 ;
        RECT 54.745 26.285 56.575 27.095 ;
        RECT 57.055 26.225 57.485 27.010 ;
        RECT 57.505 26.415 61.175 27.095 ;
        RECT 61.185 26.415 63.015 27.095 ;
        RECT 60.245 26.185 61.175 26.415 ;
        RECT 63.025 26.285 68.535 27.095 ;
        RECT 68.545 26.285 72.215 27.095 ;
        RECT 72.695 26.185 74.045 27.095 ;
        RECT 74.065 26.285 79.575 27.095 ;
        RECT 79.585 26.285 82.335 27.095 ;
        RECT 82.815 26.225 83.245 27.010 ;
        RECT 83.265 26.285 88.775 27.095 ;
        RECT 88.785 26.285 94.295 27.095 ;
        RECT 94.305 26.285 99.815 27.095 ;
        RECT 99.825 26.285 105.335 27.095 ;
        RECT 105.345 26.285 108.095 27.095 ;
        RECT 108.575 26.225 109.005 27.010 ;
        RECT 109.025 26.285 111.775 27.095 ;
        RECT 112.245 26.285 113.615 27.095 ;
      LAYER nwell ;
        RECT 5.330 23.065 113.810 25.895 ;
      LAYER pwell ;
        RECT 5.525 21.865 6.895 22.675 ;
        RECT 6.905 21.865 12.415 22.675 ;
        RECT 12.425 21.865 17.935 22.675 ;
        RECT 18.415 21.950 18.845 22.735 ;
        RECT 18.865 21.865 20.695 22.675 ;
        RECT 20.705 21.865 22.075 22.645 ;
        RECT 22.085 21.865 27.595 22.675 ;
        RECT 27.605 21.865 31.275 22.675 ;
        RECT 31.285 21.865 32.655 22.675 ;
        RECT 32.675 21.865 34.025 22.775 ;
        RECT 34.045 21.865 39.555 22.675 ;
        RECT 39.565 21.865 43.235 22.675 ;
        RECT 44.175 21.950 44.605 22.735 ;
        RECT 44.625 21.865 50.135 22.675 ;
        RECT 50.145 21.865 53.815 22.675 ;
        RECT 56.715 22.545 57.645 22.775 ;
        RECT 53.825 21.865 55.655 22.545 ;
        RECT 55.810 21.865 57.645 22.545 ;
        RECT 57.965 21.865 60.255 22.775 ;
        RECT 60.265 22.575 61.210 22.775 ;
        RECT 62.545 22.575 63.475 22.775 ;
        RECT 60.265 22.095 63.475 22.575 ;
        RECT 60.265 21.895 63.335 22.095 ;
        RECT 60.265 21.865 61.210 21.895 ;
        RECT 5.665 21.655 5.835 21.865 ;
        RECT 7.045 21.655 7.215 21.865 ;
        RECT 12.565 21.655 12.735 21.865 ;
        RECT 18.085 21.815 18.255 21.845 ;
        RECT 18.080 21.705 18.255 21.815 ;
        RECT 18.085 21.655 18.255 21.705 ;
        RECT 19.005 21.675 19.175 21.865 ;
        RECT 21.765 21.675 21.935 21.865 ;
        RECT 22.225 21.675 22.395 21.865 ;
        RECT 23.605 21.655 23.775 21.845 ;
        RECT 27.745 21.675 27.915 21.865 ;
        RECT 29.125 21.655 29.295 21.845 ;
        RECT 30.960 21.705 31.080 21.815 ;
        RECT 31.425 21.675 31.595 21.865 ;
        RECT 31.885 21.655 32.055 21.845 ;
        RECT 32.805 21.675 32.975 21.865 ;
        RECT 34.185 21.675 34.355 21.865 ;
        RECT 37.405 21.655 37.575 21.845 ;
        RECT 39.705 21.675 39.875 21.865 ;
        RECT 42.925 21.655 43.095 21.845 ;
        RECT 43.395 21.710 43.555 21.820 ;
        RECT 44.765 21.675 44.935 21.865 ;
        RECT 48.445 21.655 48.615 21.845 ;
        RECT 50.285 21.675 50.455 21.865 ;
        RECT 50.745 21.655 50.915 21.845 ;
        RECT 52.585 21.655 52.755 21.845 ;
        RECT 53.965 21.675 54.135 21.865 ;
        RECT 55.810 21.845 55.975 21.865 ;
        RECT 55.805 21.655 55.975 21.845 ;
        RECT 56.275 21.700 56.435 21.810 ;
        RECT 58.110 21.675 58.280 21.865 ;
        RECT 58.570 21.655 58.740 21.845 ;
        RECT 5.525 20.845 6.895 21.655 ;
        RECT 6.905 20.845 12.415 21.655 ;
        RECT 12.425 20.845 17.935 21.655 ;
        RECT 17.945 20.845 23.455 21.655 ;
        RECT 23.465 20.845 28.975 21.655 ;
        RECT 28.985 20.845 30.815 21.655 ;
        RECT 31.295 20.785 31.725 21.570 ;
        RECT 31.745 20.845 37.255 21.655 ;
        RECT 37.265 20.845 42.775 21.655 ;
        RECT 42.785 20.845 48.295 21.655 ;
        RECT 48.305 20.845 49.675 21.655 ;
        RECT 49.685 20.875 51.055 21.655 ;
        RECT 51.065 20.975 52.895 21.655 ;
        RECT 51.065 20.745 52.410 20.975 ;
        RECT 52.905 20.745 56.015 21.655 ;
        RECT 57.055 20.785 57.485 21.570 ;
        RECT 57.505 20.745 58.855 21.655 ;
        RECT 58.885 21.625 59.830 21.655 ;
        RECT 61.785 21.625 61.955 21.845 ;
        RECT 62.245 21.655 62.415 21.845 ;
        RECT 63.165 21.675 63.335 21.895 ;
        RECT 63.485 21.865 66.405 22.775 ;
        RECT 66.705 21.865 69.455 22.675 ;
        RECT 69.935 21.950 70.365 22.735 ;
        RECT 70.385 21.865 75.895 22.675 ;
        RECT 75.905 21.865 77.735 22.675 ;
        RECT 78.205 22.545 79.125 22.775 ;
        RECT 81.955 22.545 82.885 22.765 ;
        RECT 78.205 21.865 87.395 22.545 ;
        RECT 87.405 21.865 92.915 22.675 ;
        RECT 92.925 21.865 95.675 22.675 ;
        RECT 95.695 21.950 96.125 22.735 ;
        RECT 96.145 21.865 101.655 22.675 ;
        RECT 101.665 21.865 107.175 22.675 ;
        RECT 107.185 21.865 110.855 22.675 ;
        RECT 110.865 21.865 112.235 22.675 ;
        RECT 112.245 21.865 113.615 22.675 ;
        RECT 63.630 21.675 63.800 21.865 ;
        RECT 65.465 21.655 65.635 21.845 ;
        RECT 66.845 21.675 67.015 21.865 ;
        RECT 69.600 21.705 69.720 21.815 ;
        RECT 70.525 21.675 70.695 21.865 ;
        RECT 75.125 21.655 75.295 21.845 ;
        RECT 76.045 21.675 76.215 21.865 ;
        RECT 77.880 21.705 78.000 21.815 ;
        RECT 80.645 21.655 80.815 21.845 ;
        RECT 82.480 21.705 82.600 21.815 ;
        RECT 83.405 21.655 83.575 21.845 ;
        RECT 87.085 21.675 87.255 21.865 ;
        RECT 87.545 21.675 87.715 21.865 ;
        RECT 88.925 21.655 89.095 21.845 ;
        RECT 93.065 21.675 93.235 21.865 ;
        RECT 94.445 21.655 94.615 21.845 ;
        RECT 96.285 21.675 96.455 21.865 ;
        RECT 99.965 21.655 100.135 21.845 ;
        RECT 101.805 21.675 101.975 21.865 ;
        RECT 105.485 21.655 105.655 21.845 ;
        RECT 107.325 21.675 107.495 21.865 ;
        RECT 108.240 21.705 108.360 21.815 ;
        RECT 109.165 21.655 109.335 21.845 ;
        RECT 111.005 21.675 111.175 21.865 ;
        RECT 111.920 21.705 112.040 21.815 ;
        RECT 113.305 21.655 113.475 21.865 ;
        RECT 58.885 21.425 61.955 21.625 ;
        RECT 58.885 20.945 62.095 21.425 ;
        RECT 58.885 20.745 59.830 20.945 ;
        RECT 61.165 20.745 62.095 20.945 ;
        RECT 62.205 20.745 65.315 21.655 ;
        RECT 65.325 20.975 74.935 21.655 ;
        RECT 69.835 20.755 70.765 20.975 ;
        RECT 73.595 20.745 74.935 20.975 ;
        RECT 74.985 20.845 80.495 21.655 ;
        RECT 80.505 20.845 82.335 21.655 ;
        RECT 82.815 20.785 83.245 21.570 ;
        RECT 83.265 20.845 88.775 21.655 ;
        RECT 88.785 20.845 94.295 21.655 ;
        RECT 94.305 20.845 99.815 21.655 ;
        RECT 99.825 20.845 105.335 21.655 ;
        RECT 105.345 20.845 108.095 21.655 ;
        RECT 108.575 20.785 109.005 21.570 ;
        RECT 109.025 20.845 111.775 21.655 ;
        RECT 112.245 20.845 113.615 21.655 ;
      LAYER nwell ;
        RECT 5.330 17.625 113.810 20.455 ;
      LAYER pwell ;
        RECT 5.525 16.425 6.895 17.235 ;
        RECT 6.905 16.425 12.415 17.235 ;
        RECT 12.425 16.425 17.935 17.235 ;
        RECT 18.415 16.510 18.845 17.295 ;
        RECT 18.865 16.425 24.375 17.235 ;
        RECT 24.385 16.425 29.895 17.235 ;
        RECT 29.905 16.425 35.415 17.235 ;
        RECT 35.425 16.425 40.935 17.235 ;
        RECT 40.945 16.425 43.695 17.235 ;
        RECT 44.175 16.510 44.605 17.295 ;
        RECT 44.625 16.425 46.455 17.235 ;
        RECT 46.475 16.425 47.825 17.335 ;
        RECT 52.355 17.105 53.285 17.325 ;
        RECT 56.115 17.105 57.035 17.335 ;
        RECT 47.845 16.425 57.035 17.105 ;
        RECT 57.045 17.105 57.965 17.335 ;
        RECT 63.855 17.105 64.785 17.325 ;
        RECT 67.505 17.105 69.715 17.335 ;
        RECT 57.045 16.425 59.335 17.105 ;
        RECT 59.345 16.425 69.715 17.105 ;
        RECT 69.935 16.510 70.365 17.295 ;
        RECT 70.395 16.425 71.745 17.335 ;
        RECT 71.775 16.425 73.125 17.335 ;
        RECT 73.145 16.425 78.655 17.235 ;
        RECT 78.665 16.425 84.175 17.235 ;
        RECT 84.185 16.425 89.695 17.235 ;
        RECT 89.705 16.425 95.215 17.235 ;
        RECT 95.695 16.510 96.125 17.295 ;
        RECT 96.145 16.425 101.655 17.235 ;
        RECT 101.665 16.425 107.175 17.235 ;
        RECT 107.185 16.425 110.855 17.235 ;
        RECT 110.865 16.425 112.235 17.235 ;
        RECT 112.245 16.425 113.615 17.235 ;
        RECT 5.665 16.215 5.835 16.425 ;
        RECT 7.045 16.215 7.215 16.425 ;
        RECT 12.565 16.215 12.735 16.425 ;
        RECT 18.085 16.375 18.255 16.405 ;
        RECT 18.080 16.265 18.255 16.375 ;
        RECT 18.085 16.215 18.255 16.265 ;
        RECT 19.005 16.235 19.175 16.425 ;
        RECT 23.605 16.215 23.775 16.405 ;
        RECT 24.525 16.235 24.695 16.425 ;
        RECT 29.125 16.215 29.295 16.405 ;
        RECT 30.045 16.235 30.215 16.425 ;
        RECT 30.960 16.265 31.080 16.375 ;
        RECT 31.885 16.215 32.055 16.405 ;
        RECT 35.565 16.235 35.735 16.425 ;
        RECT 37.405 16.215 37.575 16.405 ;
        RECT 41.085 16.235 41.255 16.425 ;
        RECT 42.925 16.215 43.095 16.405 ;
        RECT 43.840 16.265 43.960 16.375 ;
        RECT 44.765 16.235 44.935 16.425 ;
        RECT 45.680 16.265 45.800 16.375 ;
        RECT 46.145 16.215 46.315 16.405 ;
        RECT 46.605 16.235 46.775 16.425 ;
        RECT 47.985 16.235 48.155 16.425 ;
        RECT 56.265 16.215 56.435 16.405 ;
        RECT 56.720 16.265 56.840 16.375 ;
        RECT 57.645 16.215 57.815 16.405 ;
        RECT 59.025 16.235 59.195 16.425 ;
        RECT 59.485 16.235 59.655 16.425 ;
        RECT 60.405 16.215 60.575 16.405 ;
        RECT 63.625 16.215 63.795 16.405 ;
        RECT 64.085 16.215 64.255 16.405 ;
        RECT 69.605 16.215 69.775 16.405 ;
        RECT 71.445 16.235 71.615 16.425 ;
        RECT 71.905 16.235 72.075 16.425 ;
        RECT 73.285 16.235 73.455 16.425 ;
        RECT 75.125 16.215 75.295 16.405 ;
        RECT 78.805 16.235 78.975 16.425 ;
        RECT 80.645 16.215 80.815 16.405 ;
        RECT 82.480 16.265 82.600 16.375 ;
        RECT 83.405 16.215 83.575 16.405 ;
        RECT 84.325 16.235 84.495 16.425 ;
        RECT 88.925 16.215 89.095 16.405 ;
        RECT 89.845 16.235 90.015 16.425 ;
        RECT 94.445 16.215 94.615 16.405 ;
        RECT 95.360 16.265 95.480 16.375 ;
        RECT 96.285 16.235 96.455 16.425 ;
        RECT 99.965 16.215 100.135 16.405 ;
        RECT 101.805 16.235 101.975 16.425 ;
        RECT 105.485 16.215 105.655 16.405 ;
        RECT 107.325 16.235 107.495 16.425 ;
        RECT 108.240 16.265 108.360 16.375 ;
        RECT 109.165 16.215 109.335 16.405 ;
        RECT 111.005 16.235 111.175 16.425 ;
        RECT 111.920 16.265 112.040 16.375 ;
        RECT 113.305 16.215 113.475 16.425 ;
        RECT 5.525 15.405 6.895 16.215 ;
        RECT 6.905 15.405 12.415 16.215 ;
        RECT 12.425 15.405 17.935 16.215 ;
        RECT 17.945 15.405 23.455 16.215 ;
        RECT 23.465 15.405 28.975 16.215 ;
        RECT 28.985 15.405 30.815 16.215 ;
        RECT 31.295 15.345 31.725 16.130 ;
        RECT 31.745 15.405 37.255 16.215 ;
        RECT 37.265 15.405 42.775 16.215 ;
        RECT 42.785 15.405 45.535 16.215 ;
        RECT 46.005 15.535 55.195 16.215 ;
        RECT 50.515 15.315 51.445 15.535 ;
        RECT 54.275 15.305 55.195 15.535 ;
        RECT 55.215 15.305 56.565 16.215 ;
        RECT 57.055 15.345 57.485 16.130 ;
        RECT 57.505 15.405 60.255 16.215 ;
        RECT 60.265 15.535 62.555 16.215 ;
        RECT 61.635 15.305 62.555 15.535 ;
        RECT 62.565 15.435 63.935 16.215 ;
        RECT 63.945 15.405 69.455 16.215 ;
        RECT 69.465 15.405 74.975 16.215 ;
        RECT 74.985 15.405 80.495 16.215 ;
        RECT 80.505 15.405 82.335 16.215 ;
        RECT 82.815 15.345 83.245 16.130 ;
        RECT 83.265 15.405 88.775 16.215 ;
        RECT 88.785 15.405 94.295 16.215 ;
        RECT 94.305 15.405 99.815 16.215 ;
        RECT 99.825 15.405 105.335 16.215 ;
        RECT 105.345 15.405 108.095 16.215 ;
        RECT 108.575 15.345 109.005 16.130 ;
        RECT 109.025 15.405 111.775 16.215 ;
        RECT 112.245 15.405 113.615 16.215 ;
      LAYER nwell ;
        RECT 5.330 12.185 113.810 15.015 ;
      LAYER pwell ;
        RECT 5.525 10.985 6.895 11.795 ;
        RECT 6.905 10.985 12.415 11.795 ;
        RECT 12.425 10.985 17.935 11.795 ;
        RECT 18.415 11.070 18.845 11.855 ;
        RECT 18.865 10.985 24.375 11.795 ;
        RECT 24.385 10.985 29.895 11.795 ;
        RECT 29.905 10.985 31.275 11.795 ;
        RECT 31.295 11.070 31.725 11.855 ;
        RECT 31.745 10.985 37.255 11.795 ;
        RECT 37.265 10.985 42.775 11.795 ;
        RECT 42.785 10.985 44.155 11.795 ;
        RECT 44.175 11.070 44.605 11.855 ;
        RECT 44.625 10.985 50.135 11.795 ;
        RECT 50.145 10.985 55.655 11.795 ;
        RECT 55.665 10.985 57.035 11.795 ;
        RECT 57.055 11.070 57.485 11.855 ;
        RECT 57.505 10.985 63.015 11.795 ;
        RECT 63.025 10.985 68.535 11.795 ;
        RECT 68.545 10.985 69.915 11.795 ;
        RECT 69.935 11.070 70.365 11.855 ;
        RECT 70.385 10.985 75.895 11.795 ;
        RECT 75.905 10.985 81.415 11.795 ;
        RECT 81.425 10.985 82.795 11.795 ;
        RECT 82.815 11.070 83.245 11.855 ;
        RECT 83.265 10.985 88.775 11.795 ;
        RECT 88.785 10.985 94.295 11.795 ;
        RECT 94.305 10.985 95.675 11.795 ;
        RECT 95.695 11.070 96.125 11.855 ;
        RECT 96.145 10.985 101.655 11.795 ;
        RECT 101.665 10.985 107.175 11.795 ;
        RECT 107.185 10.985 108.555 11.795 ;
        RECT 108.575 11.070 109.005 11.855 ;
        RECT 109.025 10.985 111.775 11.795 ;
        RECT 112.245 10.985 113.615 11.795 ;
        RECT 5.665 10.795 5.835 10.985 ;
        RECT 7.045 10.795 7.215 10.985 ;
        RECT 12.565 10.795 12.735 10.985 ;
        RECT 18.080 10.825 18.200 10.935 ;
        RECT 19.005 10.795 19.175 10.985 ;
        RECT 24.525 10.795 24.695 10.985 ;
        RECT 30.045 10.795 30.215 10.985 ;
        RECT 31.885 10.795 32.055 10.985 ;
        RECT 37.405 10.795 37.575 10.985 ;
        RECT 42.925 10.795 43.095 10.985 ;
        RECT 44.765 10.795 44.935 10.985 ;
        RECT 50.285 10.795 50.455 10.985 ;
        RECT 55.805 10.795 55.975 10.985 ;
        RECT 57.645 10.795 57.815 10.985 ;
        RECT 63.165 10.795 63.335 10.985 ;
        RECT 68.685 10.795 68.855 10.985 ;
        RECT 70.525 10.795 70.695 10.985 ;
        RECT 76.045 10.795 76.215 10.985 ;
        RECT 81.565 10.795 81.735 10.985 ;
        RECT 83.405 10.795 83.575 10.985 ;
        RECT 88.925 10.795 89.095 10.985 ;
        RECT 94.445 10.795 94.615 10.985 ;
        RECT 96.285 10.795 96.455 10.985 ;
        RECT 101.805 10.795 101.975 10.985 ;
        RECT 107.325 10.795 107.495 10.985 ;
        RECT 109.165 10.795 109.335 10.985 ;
        RECT 111.920 10.825 112.040 10.935 ;
        RECT 113.305 10.795 113.475 10.985 ;
      LAYER li1 ;
        RECT 5.520 116.875 113.620 117.045 ;
        RECT 5.605 115.785 6.815 116.875 ;
        RECT 5.605 115.075 6.125 115.615 ;
        RECT 6.295 115.245 6.815 115.785 ;
        RECT 7.065 115.945 7.245 116.705 ;
        RECT 7.425 116.115 7.755 116.875 ;
        RECT 7.065 115.775 7.740 115.945 ;
        RECT 7.925 115.800 8.195 116.705 ;
        RECT 8.365 116.440 13.710 116.875 ;
        RECT 7.570 115.630 7.740 115.775 ;
        RECT 7.005 115.225 7.345 115.595 ;
        RECT 7.570 115.300 7.845 115.630 ;
        RECT 5.605 114.325 6.815 115.075 ;
        RECT 7.570 115.045 7.740 115.300 ;
        RECT 7.075 114.875 7.740 115.045 ;
        RECT 8.015 115.000 8.195 115.800 ;
        RECT 7.075 114.495 7.245 114.875 ;
        RECT 7.425 114.325 7.755 114.705 ;
        RECT 7.935 114.495 8.195 115.000 ;
        RECT 9.950 114.870 10.290 115.700 ;
        RECT 11.770 115.190 12.120 116.440 ;
        RECT 13.885 115.785 17.395 116.875 ;
        RECT 13.885 115.095 15.535 115.615 ;
        RECT 15.705 115.265 17.395 115.785 ;
        RECT 18.485 115.710 18.775 116.875 ;
        RECT 18.945 116.440 24.290 116.875 ;
        RECT 24.465 116.440 29.810 116.875 ;
        RECT 8.365 114.325 13.710 114.870 ;
        RECT 13.885 114.325 17.395 115.095 ;
        RECT 18.485 114.325 18.775 115.050 ;
        RECT 20.530 114.870 20.870 115.700 ;
        RECT 22.350 115.190 22.700 116.440 ;
        RECT 26.050 114.870 26.390 115.700 ;
        RECT 27.870 115.190 28.220 116.440 ;
        RECT 29.985 115.785 31.195 116.875 ;
        RECT 29.985 115.075 30.505 115.615 ;
        RECT 30.675 115.245 31.195 115.785 ;
        RECT 31.365 115.710 31.655 116.875 ;
        RECT 31.830 115.685 32.085 116.565 ;
        RECT 32.255 115.735 32.560 116.875 ;
        RECT 32.900 116.495 33.230 116.875 ;
        RECT 33.410 116.325 33.580 116.615 ;
        RECT 33.750 116.415 34.000 116.875 ;
        RECT 32.780 116.155 33.580 116.325 ;
        RECT 34.170 116.365 35.040 116.705 ;
        RECT 18.945 114.325 24.290 114.870 ;
        RECT 24.465 114.325 29.810 114.870 ;
        RECT 29.985 114.325 31.195 115.075 ;
        RECT 31.365 114.325 31.655 115.050 ;
        RECT 31.830 115.035 32.040 115.685 ;
        RECT 32.780 115.565 32.950 116.155 ;
        RECT 34.170 115.985 34.340 116.365 ;
        RECT 35.275 116.245 35.445 116.705 ;
        RECT 35.615 116.415 35.985 116.875 ;
        RECT 36.280 116.275 36.450 116.615 ;
        RECT 36.620 116.445 36.950 116.875 ;
        RECT 37.185 116.275 37.355 116.615 ;
        RECT 33.120 115.815 34.340 115.985 ;
        RECT 34.510 115.905 34.970 116.195 ;
        RECT 35.275 116.075 35.835 116.245 ;
        RECT 36.280 116.105 37.355 116.275 ;
        RECT 37.525 116.375 38.205 116.705 ;
        RECT 38.420 116.375 38.670 116.705 ;
        RECT 38.840 116.415 39.090 116.875 ;
        RECT 35.665 115.935 35.835 116.075 ;
        RECT 34.510 115.895 35.475 115.905 ;
        RECT 34.170 115.725 34.340 115.815 ;
        RECT 34.800 115.735 35.475 115.895 ;
        RECT 32.210 115.535 32.950 115.565 ;
        RECT 32.210 115.235 33.125 115.535 ;
        RECT 32.800 115.060 33.125 115.235 ;
        RECT 31.830 114.505 32.085 115.035 ;
        RECT 32.255 114.325 32.560 114.785 ;
        RECT 32.805 114.705 33.125 115.060 ;
        RECT 33.295 115.275 33.835 115.645 ;
        RECT 34.170 115.555 34.575 115.725 ;
        RECT 33.295 114.875 33.535 115.275 ;
        RECT 34.015 115.105 34.235 115.385 ;
        RECT 33.705 114.935 34.235 115.105 ;
        RECT 33.705 114.705 33.875 114.935 ;
        RECT 34.405 114.775 34.575 115.555 ;
        RECT 34.745 114.945 35.095 115.565 ;
        RECT 35.265 114.945 35.475 115.735 ;
        RECT 35.665 115.765 37.165 115.935 ;
        RECT 35.665 115.075 35.835 115.765 ;
        RECT 37.525 115.595 37.695 116.375 ;
        RECT 38.500 116.245 38.670 116.375 ;
        RECT 36.005 115.425 37.695 115.595 ;
        RECT 37.865 115.815 38.330 116.205 ;
        RECT 38.500 116.075 38.895 116.245 ;
        RECT 36.005 115.245 36.175 115.425 ;
        RECT 32.805 114.535 33.875 114.705 ;
        RECT 34.045 114.325 34.235 114.765 ;
        RECT 34.405 114.495 35.355 114.775 ;
        RECT 35.665 114.685 35.925 115.075 ;
        RECT 36.345 115.005 37.135 115.255 ;
        RECT 35.575 114.515 35.925 114.685 ;
        RECT 36.135 114.325 36.465 114.785 ;
        RECT 37.340 114.715 37.510 115.425 ;
        RECT 37.865 115.225 38.035 115.815 ;
        RECT 37.680 115.005 38.035 115.225 ;
        RECT 38.205 115.005 38.555 115.625 ;
        RECT 38.725 114.715 38.895 116.075 ;
        RECT 39.260 115.905 39.585 116.690 ;
        RECT 39.065 114.855 39.525 115.905 ;
        RECT 37.340 114.545 38.195 114.715 ;
        RECT 38.400 114.545 38.895 114.715 ;
        RECT 39.065 114.325 39.395 114.685 ;
        RECT 39.755 114.585 39.925 116.705 ;
        RECT 40.095 116.375 40.425 116.875 ;
        RECT 40.595 116.205 40.850 116.705 ;
        RECT 40.100 116.035 40.850 116.205 ;
        RECT 40.100 115.045 40.330 116.035 ;
        RECT 40.500 115.215 40.850 115.865 ;
        RECT 41.025 115.785 43.615 116.875 ;
        RECT 41.025 115.095 42.235 115.615 ;
        RECT 42.405 115.265 43.615 115.785 ;
        RECT 44.245 115.710 44.535 116.875 ;
        RECT 44.705 116.440 50.050 116.875 ;
        RECT 40.100 114.875 40.850 115.045 ;
        RECT 40.095 114.325 40.425 114.705 ;
        RECT 40.595 114.585 40.850 114.875 ;
        RECT 41.025 114.325 43.615 115.095 ;
        RECT 44.245 114.325 44.535 115.050 ;
        RECT 46.290 114.870 46.630 115.700 ;
        RECT 48.110 115.190 48.460 116.440 ;
        RECT 51.185 115.735 51.415 116.875 ;
        RECT 51.585 115.725 51.915 116.705 ;
        RECT 52.085 115.735 52.295 116.875 ;
        RECT 53.025 115.735 53.255 116.875 ;
        RECT 53.425 115.725 53.755 116.705 ;
        RECT 53.925 115.735 54.135 116.875 ;
        RECT 54.365 115.785 56.955 116.875 ;
        RECT 51.165 115.315 51.495 115.565 ;
        RECT 44.705 114.325 50.050 114.870 ;
        RECT 51.185 114.325 51.415 115.145 ;
        RECT 51.665 115.125 51.915 115.725 ;
        RECT 53.005 115.315 53.335 115.565 ;
        RECT 51.585 114.495 51.915 115.125 ;
        RECT 52.085 114.325 52.295 115.145 ;
        RECT 53.025 114.325 53.255 115.145 ;
        RECT 53.505 115.125 53.755 115.725 ;
        RECT 53.425 114.495 53.755 115.125 ;
        RECT 53.925 114.325 54.135 115.145 ;
        RECT 54.365 115.095 55.575 115.615 ;
        RECT 55.745 115.265 56.955 115.785 ;
        RECT 57.125 115.710 57.415 116.875 ;
        RECT 57.585 116.440 62.930 116.875 ;
        RECT 63.105 116.440 68.450 116.875 ;
        RECT 54.365 114.325 56.955 115.095 ;
        RECT 57.125 114.325 57.415 115.050 ;
        RECT 59.170 114.870 59.510 115.700 ;
        RECT 60.990 115.190 61.340 116.440 ;
        RECT 64.690 114.870 65.030 115.700 ;
        RECT 66.510 115.190 66.860 116.440 ;
        RECT 68.625 115.785 69.835 116.875 ;
        RECT 68.625 115.075 69.145 115.615 ;
        RECT 69.315 115.245 69.835 115.785 ;
        RECT 70.005 115.710 70.295 116.875 ;
        RECT 70.465 116.440 75.810 116.875 ;
        RECT 75.985 116.440 81.330 116.875 ;
        RECT 57.585 114.325 62.930 114.870 ;
        RECT 63.105 114.325 68.450 114.870 ;
        RECT 68.625 114.325 69.835 115.075 ;
        RECT 70.005 114.325 70.295 115.050 ;
        RECT 72.050 114.870 72.390 115.700 ;
        RECT 73.870 115.190 74.220 116.440 ;
        RECT 77.570 114.870 77.910 115.700 ;
        RECT 79.390 115.190 79.740 116.440 ;
        RECT 81.505 115.785 82.715 116.875 ;
        RECT 81.505 115.075 82.025 115.615 ;
        RECT 82.195 115.245 82.715 115.785 ;
        RECT 82.885 115.710 83.175 116.875 ;
        RECT 83.345 115.785 84.555 116.875 ;
        RECT 83.345 115.075 83.865 115.615 ;
        RECT 84.035 115.245 84.555 115.785 ;
        RECT 84.765 115.735 84.995 116.875 ;
        RECT 85.165 115.725 85.495 116.705 ;
        RECT 85.665 115.735 85.875 116.875 ;
        RECT 86.105 115.785 89.615 116.875 ;
        RECT 84.745 115.315 85.075 115.565 ;
        RECT 70.465 114.325 75.810 114.870 ;
        RECT 75.985 114.325 81.330 114.870 ;
        RECT 81.505 114.325 82.715 115.075 ;
        RECT 82.885 114.325 83.175 115.050 ;
        RECT 83.345 114.325 84.555 115.075 ;
        RECT 84.765 114.325 84.995 115.145 ;
        RECT 85.245 115.125 85.495 115.725 ;
        RECT 85.165 114.495 85.495 115.125 ;
        RECT 85.665 114.325 85.875 115.145 ;
        RECT 86.105 115.095 87.755 115.615 ;
        RECT 87.925 115.265 89.615 115.785 ;
        RECT 90.745 115.735 90.975 116.875 ;
        RECT 91.145 115.725 91.475 116.705 ;
        RECT 91.645 115.735 91.855 116.875 ;
        RECT 92.085 115.785 95.595 116.875 ;
        RECT 90.725 115.315 91.055 115.565 ;
        RECT 86.105 114.325 89.615 115.095 ;
        RECT 90.745 114.325 90.975 115.145 ;
        RECT 91.225 115.125 91.475 115.725 ;
        RECT 91.145 114.495 91.475 115.125 ;
        RECT 91.645 114.325 91.855 115.145 ;
        RECT 92.085 115.095 93.735 115.615 ;
        RECT 93.905 115.265 95.595 115.785 ;
        RECT 95.765 115.710 96.055 116.875 ;
        RECT 97.185 115.735 97.415 116.875 ;
        RECT 97.585 115.725 97.915 116.705 ;
        RECT 98.085 115.735 98.295 116.875 ;
        RECT 99.450 116.205 99.705 116.705 ;
        RECT 99.875 116.375 100.205 116.875 ;
        RECT 99.450 116.035 100.200 116.205 ;
        RECT 97.165 115.315 97.495 115.565 ;
        RECT 92.085 114.325 95.595 115.095 ;
        RECT 95.765 114.325 96.055 115.050 ;
        RECT 97.185 114.325 97.415 115.145 ;
        RECT 97.665 115.125 97.915 115.725 ;
        RECT 99.450 115.215 99.800 115.865 ;
        RECT 97.585 114.495 97.915 115.125 ;
        RECT 98.085 114.325 98.295 115.145 ;
        RECT 99.970 115.045 100.200 116.035 ;
        RECT 99.450 114.875 100.200 115.045 ;
        RECT 99.450 114.585 99.705 114.875 ;
        RECT 99.875 114.325 100.205 114.705 ;
        RECT 100.375 114.585 100.545 116.705 ;
        RECT 100.715 115.905 101.040 116.690 ;
        RECT 101.210 116.415 101.460 116.875 ;
        RECT 101.630 116.375 101.880 116.705 ;
        RECT 102.095 116.375 102.775 116.705 ;
        RECT 101.630 116.245 101.800 116.375 ;
        RECT 101.405 116.075 101.800 116.245 ;
        RECT 100.775 114.855 101.235 115.905 ;
        RECT 101.405 114.715 101.575 116.075 ;
        RECT 101.970 115.815 102.435 116.205 ;
        RECT 101.745 115.005 102.095 115.625 ;
        RECT 102.265 115.225 102.435 115.815 ;
        RECT 102.605 115.595 102.775 116.375 ;
        RECT 102.945 116.275 103.115 116.615 ;
        RECT 103.350 116.445 103.680 116.875 ;
        RECT 103.850 116.275 104.020 116.615 ;
        RECT 104.315 116.415 104.685 116.875 ;
        RECT 102.945 116.105 104.020 116.275 ;
        RECT 104.855 116.245 105.025 116.705 ;
        RECT 105.260 116.365 106.130 116.705 ;
        RECT 106.300 116.415 106.550 116.875 ;
        RECT 104.465 116.075 105.025 116.245 ;
        RECT 104.465 115.935 104.635 116.075 ;
        RECT 103.135 115.765 104.635 115.935 ;
        RECT 105.330 115.905 105.790 116.195 ;
        RECT 102.605 115.425 104.295 115.595 ;
        RECT 102.265 115.005 102.620 115.225 ;
        RECT 102.790 114.715 102.960 115.425 ;
        RECT 103.165 115.005 103.955 115.255 ;
        RECT 104.125 115.245 104.295 115.425 ;
        RECT 104.465 115.075 104.635 115.765 ;
        RECT 100.905 114.325 101.235 114.685 ;
        RECT 101.405 114.545 101.900 114.715 ;
        RECT 102.105 114.545 102.960 114.715 ;
        RECT 103.835 114.325 104.165 114.785 ;
        RECT 104.375 114.685 104.635 115.075 ;
        RECT 104.825 115.895 105.790 115.905 ;
        RECT 105.960 115.985 106.130 116.365 ;
        RECT 106.720 116.325 106.890 116.615 ;
        RECT 107.070 116.495 107.400 116.875 ;
        RECT 106.720 116.155 107.520 116.325 ;
        RECT 104.825 115.735 105.500 115.895 ;
        RECT 105.960 115.815 107.180 115.985 ;
        RECT 104.825 114.945 105.035 115.735 ;
        RECT 105.960 115.725 106.130 115.815 ;
        RECT 105.205 114.945 105.555 115.565 ;
        RECT 105.725 115.555 106.130 115.725 ;
        RECT 105.725 114.775 105.895 115.555 ;
        RECT 106.065 115.105 106.285 115.385 ;
        RECT 106.465 115.275 107.005 115.645 ;
        RECT 107.350 115.565 107.520 116.155 ;
        RECT 107.740 115.735 108.045 116.875 ;
        RECT 108.215 115.685 108.470 116.565 ;
        RECT 108.645 115.710 108.935 116.875 ;
        RECT 109.105 115.785 111.695 116.875 ;
        RECT 107.350 115.535 108.090 115.565 ;
        RECT 106.065 114.935 106.595 115.105 ;
        RECT 104.375 114.515 104.725 114.685 ;
        RECT 104.945 114.495 105.895 114.775 ;
        RECT 106.065 114.325 106.255 114.765 ;
        RECT 106.425 114.705 106.595 114.935 ;
        RECT 106.765 114.875 107.005 115.275 ;
        RECT 107.175 115.235 108.090 115.535 ;
        RECT 107.175 115.060 107.500 115.235 ;
        RECT 107.175 114.705 107.495 115.060 ;
        RECT 108.260 115.035 108.470 115.685 ;
        RECT 109.105 115.095 110.315 115.615 ;
        RECT 110.485 115.265 111.695 115.785 ;
        RECT 112.325 115.785 113.535 116.875 ;
        RECT 112.325 115.245 112.845 115.785 ;
        RECT 106.425 114.535 107.495 114.705 ;
        RECT 107.740 114.325 108.045 114.785 ;
        RECT 108.215 114.505 108.470 115.035 ;
        RECT 108.645 114.325 108.935 115.050 ;
        RECT 109.105 114.325 111.695 115.095 ;
        RECT 113.015 115.075 113.535 115.615 ;
        RECT 112.325 114.325 113.535 115.075 ;
        RECT 5.520 114.155 113.620 114.325 ;
        RECT 5.605 113.405 6.815 114.155 ;
        RECT 5.605 112.865 6.125 113.405 ;
        RECT 6.985 113.385 9.575 114.155 ;
        RECT 10.210 113.445 10.465 113.975 ;
        RECT 10.635 113.695 10.940 114.155 ;
        RECT 11.185 113.775 12.255 113.945 ;
        RECT 6.295 112.695 6.815 113.235 ;
        RECT 6.985 112.865 8.195 113.385 ;
        RECT 8.365 112.695 9.575 113.215 ;
        RECT 5.605 111.605 6.815 112.695 ;
        RECT 6.985 111.605 9.575 112.695 ;
        RECT 10.210 112.795 10.420 113.445 ;
        RECT 11.185 113.420 11.505 113.775 ;
        RECT 11.180 113.245 11.505 113.420 ;
        RECT 10.590 112.945 11.505 113.245 ;
        RECT 11.675 113.205 11.915 113.605 ;
        RECT 12.085 113.545 12.255 113.775 ;
        RECT 12.425 113.715 12.615 114.155 ;
        RECT 12.785 113.705 13.735 113.985 ;
        RECT 13.955 113.795 14.305 113.965 ;
        RECT 12.085 113.375 12.615 113.545 ;
        RECT 10.590 112.915 11.330 112.945 ;
        RECT 10.210 111.915 10.465 112.795 ;
        RECT 10.635 111.605 10.940 112.745 ;
        RECT 11.160 112.325 11.330 112.915 ;
        RECT 11.675 112.835 12.215 113.205 ;
        RECT 12.395 113.095 12.615 113.375 ;
        RECT 12.785 112.925 12.955 113.705 ;
        RECT 12.550 112.755 12.955 112.925 ;
        RECT 13.125 112.915 13.475 113.535 ;
        RECT 12.550 112.665 12.720 112.755 ;
        RECT 13.645 112.745 13.855 113.535 ;
        RECT 11.500 112.495 12.720 112.665 ;
        RECT 13.180 112.585 13.855 112.745 ;
        RECT 11.160 112.155 11.960 112.325 ;
        RECT 11.280 111.605 11.610 111.985 ;
        RECT 11.790 111.865 11.960 112.155 ;
        RECT 12.550 112.115 12.720 112.495 ;
        RECT 12.890 112.575 13.855 112.585 ;
        RECT 14.045 113.405 14.305 113.795 ;
        RECT 14.515 113.695 14.845 114.155 ;
        RECT 15.720 113.765 16.575 113.935 ;
        RECT 16.780 113.765 17.275 113.935 ;
        RECT 17.445 113.795 17.775 114.155 ;
        RECT 14.045 112.715 14.215 113.405 ;
        RECT 14.385 113.055 14.555 113.235 ;
        RECT 14.725 113.225 15.515 113.475 ;
        RECT 15.720 113.055 15.890 113.765 ;
        RECT 16.060 113.255 16.415 113.475 ;
        RECT 14.385 112.885 16.075 113.055 ;
        RECT 12.890 112.285 13.350 112.575 ;
        RECT 14.045 112.545 15.545 112.715 ;
        RECT 14.045 112.405 14.215 112.545 ;
        RECT 13.655 112.235 14.215 112.405 ;
        RECT 12.130 111.605 12.380 112.065 ;
        RECT 12.550 111.775 13.420 112.115 ;
        RECT 13.655 111.775 13.825 112.235 ;
        RECT 14.660 112.205 15.735 112.375 ;
        RECT 13.995 111.605 14.365 112.065 ;
        RECT 14.660 111.865 14.830 112.205 ;
        RECT 15.000 111.605 15.330 112.035 ;
        RECT 15.565 111.865 15.735 112.205 ;
        RECT 15.905 112.105 16.075 112.885 ;
        RECT 16.245 112.665 16.415 113.255 ;
        RECT 16.585 112.855 16.935 113.475 ;
        RECT 16.245 112.275 16.710 112.665 ;
        RECT 17.105 112.405 17.275 113.765 ;
        RECT 17.445 112.575 17.905 113.625 ;
        RECT 16.880 112.235 17.275 112.405 ;
        RECT 16.880 112.105 17.050 112.235 ;
        RECT 15.905 111.775 16.585 112.105 ;
        RECT 16.800 111.775 17.050 112.105 ;
        RECT 17.220 111.605 17.470 112.065 ;
        RECT 17.640 111.790 17.965 112.575 ;
        RECT 18.135 111.775 18.305 113.895 ;
        RECT 18.475 113.775 18.805 114.155 ;
        RECT 18.975 113.605 19.230 113.895 ;
        RECT 18.480 113.435 19.230 113.605 ;
        RECT 18.480 112.445 18.710 113.435 ;
        RECT 19.405 113.385 21.075 114.155 ;
        RECT 21.250 113.605 21.505 113.895 ;
        RECT 21.675 113.775 22.005 114.155 ;
        RECT 21.250 113.435 22.000 113.605 ;
        RECT 18.880 112.615 19.230 113.265 ;
        RECT 19.405 112.865 20.155 113.385 ;
        RECT 20.325 112.695 21.075 113.215 ;
        RECT 18.480 112.275 19.230 112.445 ;
        RECT 18.475 111.605 18.805 112.105 ;
        RECT 18.975 111.775 19.230 112.275 ;
        RECT 19.405 111.605 21.075 112.695 ;
        RECT 21.250 112.615 21.600 113.265 ;
        RECT 21.770 112.445 22.000 113.435 ;
        RECT 21.250 112.275 22.000 112.445 ;
        RECT 21.250 111.775 21.505 112.275 ;
        RECT 21.675 111.605 22.005 112.105 ;
        RECT 22.175 111.775 22.345 113.895 ;
        RECT 22.705 113.795 23.035 114.155 ;
        RECT 23.205 113.765 23.700 113.935 ;
        RECT 23.905 113.765 24.760 113.935 ;
        RECT 22.575 112.575 23.035 113.625 ;
        RECT 22.515 111.790 22.840 112.575 ;
        RECT 23.205 112.405 23.375 113.765 ;
        RECT 23.545 112.855 23.895 113.475 ;
        RECT 24.065 113.255 24.420 113.475 ;
        RECT 24.065 112.665 24.235 113.255 ;
        RECT 24.590 113.055 24.760 113.765 ;
        RECT 25.635 113.695 25.965 114.155 ;
        RECT 26.175 113.795 26.525 113.965 ;
        RECT 24.965 113.225 25.755 113.475 ;
        RECT 26.175 113.405 26.435 113.795 ;
        RECT 26.745 113.705 27.695 113.985 ;
        RECT 27.865 113.715 28.055 114.155 ;
        RECT 28.225 113.775 29.295 113.945 ;
        RECT 25.925 113.055 26.095 113.235 ;
        RECT 23.205 112.235 23.600 112.405 ;
        RECT 23.770 112.275 24.235 112.665 ;
        RECT 24.405 112.885 26.095 113.055 ;
        RECT 23.430 112.105 23.600 112.235 ;
        RECT 24.405 112.105 24.575 112.885 ;
        RECT 26.265 112.715 26.435 113.405 ;
        RECT 24.935 112.545 26.435 112.715 ;
        RECT 26.625 112.745 26.835 113.535 ;
        RECT 27.005 112.915 27.355 113.535 ;
        RECT 27.525 112.925 27.695 113.705 ;
        RECT 28.225 113.545 28.395 113.775 ;
        RECT 27.865 113.375 28.395 113.545 ;
        RECT 27.865 113.095 28.085 113.375 ;
        RECT 28.565 113.205 28.805 113.605 ;
        RECT 27.525 112.755 27.930 112.925 ;
        RECT 28.265 112.835 28.805 113.205 ;
        RECT 28.975 113.420 29.295 113.775 ;
        RECT 29.540 113.695 29.845 114.155 ;
        RECT 30.015 113.445 30.270 113.975 ;
        RECT 28.975 113.245 29.300 113.420 ;
        RECT 28.975 112.945 29.890 113.245 ;
        RECT 29.150 112.915 29.890 112.945 ;
        RECT 26.625 112.585 27.300 112.745 ;
        RECT 27.760 112.665 27.930 112.755 ;
        RECT 26.625 112.575 27.590 112.585 ;
        RECT 26.265 112.405 26.435 112.545 ;
        RECT 23.010 111.605 23.260 112.065 ;
        RECT 23.430 111.775 23.680 112.105 ;
        RECT 23.895 111.775 24.575 112.105 ;
        RECT 24.745 112.205 25.820 112.375 ;
        RECT 26.265 112.235 26.825 112.405 ;
        RECT 27.130 112.285 27.590 112.575 ;
        RECT 27.760 112.495 28.980 112.665 ;
        RECT 24.745 111.865 24.915 112.205 ;
        RECT 25.150 111.605 25.480 112.035 ;
        RECT 25.650 111.865 25.820 112.205 ;
        RECT 26.115 111.605 26.485 112.065 ;
        RECT 26.655 111.775 26.825 112.235 ;
        RECT 27.760 112.115 27.930 112.495 ;
        RECT 29.150 112.325 29.320 112.915 ;
        RECT 30.060 112.795 30.270 113.445 ;
        RECT 31.365 113.430 31.655 114.155 ;
        RECT 31.825 113.610 37.170 114.155 ;
        RECT 27.060 111.775 27.930 112.115 ;
        RECT 28.520 112.155 29.320 112.325 ;
        RECT 28.100 111.605 28.350 112.065 ;
        RECT 28.520 111.865 28.690 112.155 ;
        RECT 28.870 111.605 29.200 111.985 ;
        RECT 29.540 111.605 29.845 112.745 ;
        RECT 30.015 111.915 30.270 112.795 ;
        RECT 33.410 112.780 33.750 113.610 ;
        RECT 38.270 113.605 38.525 113.895 ;
        RECT 38.695 113.775 39.025 114.155 ;
        RECT 38.270 113.435 39.020 113.605 ;
        RECT 31.365 111.605 31.655 112.770 ;
        RECT 35.230 112.040 35.580 113.290 ;
        RECT 38.270 112.615 38.620 113.265 ;
        RECT 38.790 112.445 39.020 113.435 ;
        RECT 38.270 112.275 39.020 112.445 ;
        RECT 31.825 111.605 37.170 112.040 ;
        RECT 38.270 111.775 38.525 112.275 ;
        RECT 38.695 111.605 39.025 112.105 ;
        RECT 39.195 111.775 39.365 113.895 ;
        RECT 39.725 113.795 40.055 114.155 ;
        RECT 40.225 113.765 40.720 113.935 ;
        RECT 40.925 113.765 41.780 113.935 ;
        RECT 39.595 112.575 40.055 113.625 ;
        RECT 39.535 111.790 39.860 112.575 ;
        RECT 40.225 112.405 40.395 113.765 ;
        RECT 40.565 112.855 40.915 113.475 ;
        RECT 41.085 113.255 41.440 113.475 ;
        RECT 41.085 112.665 41.255 113.255 ;
        RECT 41.610 113.055 41.780 113.765 ;
        RECT 42.655 113.695 42.985 114.155 ;
        RECT 43.195 113.795 43.545 113.965 ;
        RECT 41.985 113.225 42.775 113.475 ;
        RECT 43.195 113.405 43.455 113.795 ;
        RECT 43.765 113.705 44.715 113.985 ;
        RECT 44.885 113.715 45.075 114.155 ;
        RECT 45.245 113.775 46.315 113.945 ;
        RECT 42.945 113.055 43.115 113.235 ;
        RECT 40.225 112.235 40.620 112.405 ;
        RECT 40.790 112.275 41.255 112.665 ;
        RECT 41.425 112.885 43.115 113.055 ;
        RECT 40.450 112.105 40.620 112.235 ;
        RECT 41.425 112.105 41.595 112.885 ;
        RECT 43.285 112.715 43.455 113.405 ;
        RECT 41.955 112.545 43.455 112.715 ;
        RECT 43.645 112.745 43.855 113.535 ;
        RECT 44.025 112.915 44.375 113.535 ;
        RECT 44.545 112.925 44.715 113.705 ;
        RECT 45.245 113.545 45.415 113.775 ;
        RECT 44.885 113.375 45.415 113.545 ;
        RECT 44.885 113.095 45.105 113.375 ;
        RECT 45.585 113.205 45.825 113.605 ;
        RECT 44.545 112.755 44.950 112.925 ;
        RECT 45.285 112.835 45.825 113.205 ;
        RECT 45.995 113.420 46.315 113.775 ;
        RECT 46.560 113.695 46.865 114.155 ;
        RECT 47.035 113.445 47.290 113.975 ;
        RECT 45.995 113.245 46.320 113.420 ;
        RECT 45.995 112.945 46.910 113.245 ;
        RECT 46.170 112.915 46.910 112.945 ;
        RECT 43.645 112.585 44.320 112.745 ;
        RECT 44.780 112.665 44.950 112.755 ;
        RECT 43.645 112.575 44.610 112.585 ;
        RECT 43.285 112.405 43.455 112.545 ;
        RECT 40.030 111.605 40.280 112.065 ;
        RECT 40.450 111.775 40.700 112.105 ;
        RECT 40.915 111.775 41.595 112.105 ;
        RECT 41.765 112.205 42.840 112.375 ;
        RECT 43.285 112.235 43.845 112.405 ;
        RECT 44.150 112.285 44.610 112.575 ;
        RECT 44.780 112.495 46.000 112.665 ;
        RECT 41.765 111.865 41.935 112.205 ;
        RECT 42.170 111.605 42.500 112.035 ;
        RECT 42.670 111.865 42.840 112.205 ;
        RECT 43.135 111.605 43.505 112.065 ;
        RECT 43.675 111.775 43.845 112.235 ;
        RECT 44.780 112.115 44.950 112.495 ;
        RECT 46.170 112.325 46.340 112.915 ;
        RECT 47.080 112.795 47.290 113.445 ;
        RECT 47.930 113.605 48.185 113.895 ;
        RECT 48.355 113.775 48.685 114.155 ;
        RECT 47.930 113.435 48.680 113.605 ;
        RECT 44.080 111.775 44.950 112.115 ;
        RECT 45.540 112.155 46.340 112.325 ;
        RECT 45.120 111.605 45.370 112.065 ;
        RECT 45.540 111.865 45.710 112.155 ;
        RECT 45.890 111.605 46.220 111.985 ;
        RECT 46.560 111.605 46.865 112.745 ;
        RECT 47.035 111.915 47.290 112.795 ;
        RECT 47.930 112.615 48.280 113.265 ;
        RECT 48.450 112.445 48.680 113.435 ;
        RECT 47.930 112.275 48.680 112.445 ;
        RECT 47.930 111.775 48.185 112.275 ;
        RECT 48.355 111.605 48.685 112.105 ;
        RECT 48.855 111.775 49.025 113.895 ;
        RECT 49.385 113.795 49.715 114.155 ;
        RECT 49.885 113.765 50.380 113.935 ;
        RECT 50.585 113.765 51.440 113.935 ;
        RECT 49.255 112.575 49.715 113.625 ;
        RECT 49.195 111.790 49.520 112.575 ;
        RECT 49.885 112.405 50.055 113.765 ;
        RECT 50.225 112.855 50.575 113.475 ;
        RECT 50.745 113.255 51.100 113.475 ;
        RECT 50.745 112.665 50.915 113.255 ;
        RECT 51.270 113.055 51.440 113.765 ;
        RECT 52.315 113.695 52.645 114.155 ;
        RECT 52.855 113.795 53.205 113.965 ;
        RECT 51.645 113.225 52.435 113.475 ;
        RECT 52.855 113.405 53.115 113.795 ;
        RECT 53.425 113.705 54.375 113.985 ;
        RECT 54.545 113.715 54.735 114.155 ;
        RECT 54.905 113.775 55.975 113.945 ;
        RECT 52.605 113.055 52.775 113.235 ;
        RECT 49.885 112.235 50.280 112.405 ;
        RECT 50.450 112.275 50.915 112.665 ;
        RECT 51.085 112.885 52.775 113.055 ;
        RECT 50.110 112.105 50.280 112.235 ;
        RECT 51.085 112.105 51.255 112.885 ;
        RECT 52.945 112.715 53.115 113.405 ;
        RECT 51.615 112.545 53.115 112.715 ;
        RECT 53.305 112.745 53.515 113.535 ;
        RECT 53.685 112.915 54.035 113.535 ;
        RECT 54.205 112.925 54.375 113.705 ;
        RECT 54.905 113.545 55.075 113.775 ;
        RECT 54.545 113.375 55.075 113.545 ;
        RECT 54.545 113.095 54.765 113.375 ;
        RECT 55.245 113.205 55.485 113.605 ;
        RECT 54.205 112.755 54.610 112.925 ;
        RECT 54.945 112.835 55.485 113.205 ;
        RECT 55.655 113.420 55.975 113.775 ;
        RECT 56.220 113.695 56.525 114.155 ;
        RECT 56.695 113.445 56.950 113.975 ;
        RECT 55.655 113.245 55.980 113.420 ;
        RECT 55.655 112.945 56.570 113.245 ;
        RECT 55.830 112.915 56.570 112.945 ;
        RECT 53.305 112.585 53.980 112.745 ;
        RECT 54.440 112.665 54.610 112.755 ;
        RECT 53.305 112.575 54.270 112.585 ;
        RECT 52.945 112.405 53.115 112.545 ;
        RECT 49.690 111.605 49.940 112.065 ;
        RECT 50.110 111.775 50.360 112.105 ;
        RECT 50.575 111.775 51.255 112.105 ;
        RECT 51.425 112.205 52.500 112.375 ;
        RECT 52.945 112.235 53.505 112.405 ;
        RECT 53.810 112.285 54.270 112.575 ;
        RECT 54.440 112.495 55.660 112.665 ;
        RECT 51.425 111.865 51.595 112.205 ;
        RECT 51.830 111.605 52.160 112.035 ;
        RECT 52.330 111.865 52.500 112.205 ;
        RECT 52.795 111.605 53.165 112.065 ;
        RECT 53.335 111.775 53.505 112.235 ;
        RECT 54.440 112.115 54.610 112.495 ;
        RECT 55.830 112.325 56.000 112.915 ;
        RECT 56.740 112.795 56.950 113.445 ;
        RECT 57.125 113.430 57.415 114.155 ;
        RECT 57.585 113.385 61.095 114.155 ;
        RECT 62.190 113.605 62.445 113.895 ;
        RECT 62.615 113.775 62.945 114.155 ;
        RECT 62.190 113.435 62.940 113.605 ;
        RECT 57.585 112.865 59.235 113.385 ;
        RECT 53.740 111.775 54.610 112.115 ;
        RECT 55.200 112.155 56.000 112.325 ;
        RECT 54.780 111.605 55.030 112.065 ;
        RECT 55.200 111.865 55.370 112.155 ;
        RECT 55.550 111.605 55.880 111.985 ;
        RECT 56.220 111.605 56.525 112.745 ;
        RECT 56.695 111.915 56.950 112.795 ;
        RECT 57.125 111.605 57.415 112.770 ;
        RECT 59.405 112.695 61.095 113.215 ;
        RECT 57.585 111.605 61.095 112.695 ;
        RECT 62.190 112.615 62.540 113.265 ;
        RECT 62.710 112.445 62.940 113.435 ;
        RECT 62.190 112.275 62.940 112.445 ;
        RECT 62.190 111.775 62.445 112.275 ;
        RECT 62.615 111.605 62.945 112.105 ;
        RECT 63.115 111.775 63.285 113.895 ;
        RECT 63.645 113.795 63.975 114.155 ;
        RECT 64.145 113.765 64.640 113.935 ;
        RECT 64.845 113.765 65.700 113.935 ;
        RECT 63.515 112.575 63.975 113.625 ;
        RECT 63.455 111.790 63.780 112.575 ;
        RECT 64.145 112.405 64.315 113.765 ;
        RECT 64.485 112.855 64.835 113.475 ;
        RECT 65.005 113.255 65.360 113.475 ;
        RECT 65.005 112.665 65.175 113.255 ;
        RECT 65.530 113.055 65.700 113.765 ;
        RECT 66.575 113.695 66.905 114.155 ;
        RECT 67.115 113.795 67.465 113.965 ;
        RECT 65.905 113.225 66.695 113.475 ;
        RECT 67.115 113.405 67.375 113.795 ;
        RECT 67.685 113.705 68.635 113.985 ;
        RECT 68.805 113.715 68.995 114.155 ;
        RECT 69.165 113.775 70.235 113.945 ;
        RECT 66.865 113.055 67.035 113.235 ;
        RECT 64.145 112.235 64.540 112.405 ;
        RECT 64.710 112.275 65.175 112.665 ;
        RECT 65.345 112.885 67.035 113.055 ;
        RECT 64.370 112.105 64.540 112.235 ;
        RECT 65.345 112.105 65.515 112.885 ;
        RECT 67.205 112.715 67.375 113.405 ;
        RECT 65.875 112.545 67.375 112.715 ;
        RECT 67.565 112.745 67.775 113.535 ;
        RECT 67.945 112.915 68.295 113.535 ;
        RECT 68.465 112.925 68.635 113.705 ;
        RECT 69.165 113.545 69.335 113.775 ;
        RECT 68.805 113.375 69.335 113.545 ;
        RECT 68.805 113.095 69.025 113.375 ;
        RECT 69.505 113.205 69.745 113.605 ;
        RECT 68.465 112.755 68.870 112.925 ;
        RECT 69.205 112.835 69.745 113.205 ;
        RECT 69.915 113.420 70.235 113.775 ;
        RECT 70.480 113.695 70.785 114.155 ;
        RECT 70.955 113.445 71.210 113.975 ;
        RECT 69.915 113.245 70.240 113.420 ;
        RECT 69.915 112.945 70.830 113.245 ;
        RECT 70.090 112.915 70.830 112.945 ;
        RECT 67.565 112.585 68.240 112.745 ;
        RECT 68.700 112.665 68.870 112.755 ;
        RECT 67.565 112.575 68.530 112.585 ;
        RECT 67.205 112.405 67.375 112.545 ;
        RECT 63.950 111.605 64.200 112.065 ;
        RECT 64.370 111.775 64.620 112.105 ;
        RECT 64.835 111.775 65.515 112.105 ;
        RECT 65.685 112.205 66.760 112.375 ;
        RECT 67.205 112.235 67.765 112.405 ;
        RECT 68.070 112.285 68.530 112.575 ;
        RECT 68.700 112.495 69.920 112.665 ;
        RECT 65.685 111.865 65.855 112.205 ;
        RECT 66.090 111.605 66.420 112.035 ;
        RECT 66.590 111.865 66.760 112.205 ;
        RECT 67.055 111.605 67.425 112.065 ;
        RECT 67.595 111.775 67.765 112.235 ;
        RECT 68.700 112.115 68.870 112.495 ;
        RECT 70.090 112.325 70.260 112.915 ;
        RECT 71.000 112.795 71.210 113.445 ;
        RECT 71.390 113.605 71.645 113.895 ;
        RECT 71.815 113.775 72.145 114.155 ;
        RECT 71.390 113.435 72.140 113.605 ;
        RECT 68.000 111.775 68.870 112.115 ;
        RECT 69.460 112.155 70.260 112.325 ;
        RECT 69.040 111.605 69.290 112.065 ;
        RECT 69.460 111.865 69.630 112.155 ;
        RECT 69.810 111.605 70.140 111.985 ;
        RECT 70.480 111.605 70.785 112.745 ;
        RECT 70.955 111.915 71.210 112.795 ;
        RECT 71.390 112.615 71.740 113.265 ;
        RECT 71.910 112.445 72.140 113.435 ;
        RECT 71.390 112.275 72.140 112.445 ;
        RECT 71.390 111.775 71.645 112.275 ;
        RECT 71.815 111.605 72.145 112.105 ;
        RECT 72.315 111.775 72.485 113.895 ;
        RECT 72.845 113.795 73.175 114.155 ;
        RECT 73.345 113.765 73.840 113.935 ;
        RECT 74.045 113.765 74.900 113.935 ;
        RECT 72.715 112.575 73.175 113.625 ;
        RECT 72.655 111.790 72.980 112.575 ;
        RECT 73.345 112.405 73.515 113.765 ;
        RECT 73.685 112.855 74.035 113.475 ;
        RECT 74.205 113.255 74.560 113.475 ;
        RECT 74.205 112.665 74.375 113.255 ;
        RECT 74.730 113.055 74.900 113.765 ;
        RECT 75.775 113.695 76.105 114.155 ;
        RECT 76.315 113.795 76.665 113.965 ;
        RECT 75.105 113.225 75.895 113.475 ;
        RECT 76.315 113.405 76.575 113.795 ;
        RECT 76.885 113.705 77.835 113.985 ;
        RECT 78.005 113.715 78.195 114.155 ;
        RECT 78.365 113.775 79.435 113.945 ;
        RECT 76.065 113.055 76.235 113.235 ;
        RECT 73.345 112.235 73.740 112.405 ;
        RECT 73.910 112.275 74.375 112.665 ;
        RECT 74.545 112.885 76.235 113.055 ;
        RECT 73.570 112.105 73.740 112.235 ;
        RECT 74.545 112.105 74.715 112.885 ;
        RECT 76.405 112.715 76.575 113.405 ;
        RECT 75.075 112.545 76.575 112.715 ;
        RECT 76.765 112.745 76.975 113.535 ;
        RECT 77.145 112.915 77.495 113.535 ;
        RECT 77.665 112.925 77.835 113.705 ;
        RECT 78.365 113.545 78.535 113.775 ;
        RECT 78.005 113.375 78.535 113.545 ;
        RECT 78.005 113.095 78.225 113.375 ;
        RECT 78.705 113.205 78.945 113.605 ;
        RECT 77.665 112.755 78.070 112.925 ;
        RECT 78.405 112.835 78.945 113.205 ;
        RECT 79.115 113.420 79.435 113.775 ;
        RECT 79.680 113.695 79.985 114.155 ;
        RECT 80.155 113.445 80.410 113.975 ;
        RECT 79.115 113.245 79.440 113.420 ;
        RECT 79.115 112.945 80.030 113.245 ;
        RECT 79.290 112.915 80.030 112.945 ;
        RECT 76.765 112.585 77.440 112.745 ;
        RECT 77.900 112.665 78.070 112.755 ;
        RECT 76.765 112.575 77.730 112.585 ;
        RECT 76.405 112.405 76.575 112.545 ;
        RECT 73.150 111.605 73.400 112.065 ;
        RECT 73.570 111.775 73.820 112.105 ;
        RECT 74.035 111.775 74.715 112.105 ;
        RECT 74.885 112.205 75.960 112.375 ;
        RECT 76.405 112.235 76.965 112.405 ;
        RECT 77.270 112.285 77.730 112.575 ;
        RECT 77.900 112.495 79.120 112.665 ;
        RECT 74.885 111.865 75.055 112.205 ;
        RECT 75.290 111.605 75.620 112.035 ;
        RECT 75.790 111.865 75.960 112.205 ;
        RECT 76.255 111.605 76.625 112.065 ;
        RECT 76.795 111.775 76.965 112.235 ;
        RECT 77.900 112.115 78.070 112.495 ;
        RECT 79.290 112.325 79.460 112.915 ;
        RECT 80.200 112.795 80.410 113.445 ;
        RECT 80.645 113.335 80.855 114.155 ;
        RECT 81.025 113.355 81.355 113.985 ;
        RECT 77.200 111.775 78.070 112.115 ;
        RECT 78.660 112.155 79.460 112.325 ;
        RECT 78.240 111.605 78.490 112.065 ;
        RECT 78.660 111.865 78.830 112.155 ;
        RECT 79.010 111.605 79.340 111.985 ;
        RECT 79.680 111.605 79.985 112.745 ;
        RECT 80.155 111.915 80.410 112.795 ;
        RECT 81.025 112.755 81.275 113.355 ;
        RECT 81.525 113.335 81.755 114.155 ;
        RECT 82.885 113.430 83.175 114.155 ;
        RECT 83.350 113.605 83.605 113.895 ;
        RECT 83.775 113.775 84.105 114.155 ;
        RECT 83.350 113.435 84.100 113.605 ;
        RECT 81.445 112.915 81.775 113.165 ;
        RECT 80.645 111.605 80.855 112.745 ;
        RECT 81.025 111.775 81.355 112.755 ;
        RECT 81.525 111.605 81.755 112.745 ;
        RECT 82.885 111.605 83.175 112.770 ;
        RECT 83.350 112.615 83.700 113.265 ;
        RECT 83.870 112.445 84.100 113.435 ;
        RECT 83.350 112.275 84.100 112.445 ;
        RECT 83.350 111.775 83.605 112.275 ;
        RECT 83.775 111.605 84.105 112.105 ;
        RECT 84.275 111.775 84.445 113.895 ;
        RECT 84.805 113.795 85.135 114.155 ;
        RECT 85.305 113.765 85.800 113.935 ;
        RECT 86.005 113.765 86.860 113.935 ;
        RECT 84.675 112.575 85.135 113.625 ;
        RECT 84.615 111.790 84.940 112.575 ;
        RECT 85.305 112.405 85.475 113.765 ;
        RECT 85.645 112.855 85.995 113.475 ;
        RECT 86.165 113.255 86.520 113.475 ;
        RECT 86.165 112.665 86.335 113.255 ;
        RECT 86.690 113.055 86.860 113.765 ;
        RECT 87.735 113.695 88.065 114.155 ;
        RECT 88.275 113.795 88.625 113.965 ;
        RECT 87.065 113.225 87.855 113.475 ;
        RECT 88.275 113.405 88.535 113.795 ;
        RECT 88.845 113.705 89.795 113.985 ;
        RECT 89.965 113.715 90.155 114.155 ;
        RECT 90.325 113.775 91.395 113.945 ;
        RECT 88.025 113.055 88.195 113.235 ;
        RECT 85.305 112.235 85.700 112.405 ;
        RECT 85.870 112.275 86.335 112.665 ;
        RECT 86.505 112.885 88.195 113.055 ;
        RECT 85.530 112.105 85.700 112.235 ;
        RECT 86.505 112.105 86.675 112.885 ;
        RECT 88.365 112.715 88.535 113.405 ;
        RECT 87.035 112.545 88.535 112.715 ;
        RECT 88.725 112.745 88.935 113.535 ;
        RECT 89.105 112.915 89.455 113.535 ;
        RECT 89.625 112.925 89.795 113.705 ;
        RECT 90.325 113.545 90.495 113.775 ;
        RECT 89.965 113.375 90.495 113.545 ;
        RECT 89.965 113.095 90.185 113.375 ;
        RECT 90.665 113.205 90.905 113.605 ;
        RECT 89.625 112.755 90.030 112.925 ;
        RECT 90.365 112.835 90.905 113.205 ;
        RECT 91.075 113.420 91.395 113.775 ;
        RECT 91.640 113.695 91.945 114.155 ;
        RECT 92.115 113.445 92.370 113.975 ;
        RECT 91.075 113.245 91.400 113.420 ;
        RECT 91.075 112.945 91.990 113.245 ;
        RECT 91.250 112.915 91.990 112.945 ;
        RECT 88.725 112.585 89.400 112.745 ;
        RECT 89.860 112.665 90.030 112.755 ;
        RECT 88.725 112.575 89.690 112.585 ;
        RECT 88.365 112.405 88.535 112.545 ;
        RECT 85.110 111.605 85.360 112.065 ;
        RECT 85.530 111.775 85.780 112.105 ;
        RECT 85.995 111.775 86.675 112.105 ;
        RECT 86.845 112.205 87.920 112.375 ;
        RECT 88.365 112.235 88.925 112.405 ;
        RECT 89.230 112.285 89.690 112.575 ;
        RECT 89.860 112.495 91.080 112.665 ;
        RECT 86.845 111.865 87.015 112.205 ;
        RECT 87.250 111.605 87.580 112.035 ;
        RECT 87.750 111.865 87.920 112.205 ;
        RECT 88.215 111.605 88.585 112.065 ;
        RECT 88.755 111.775 88.925 112.235 ;
        RECT 89.860 112.115 90.030 112.495 ;
        RECT 91.250 112.325 91.420 112.915 ;
        RECT 92.160 112.795 92.370 113.445 ;
        RECT 92.550 113.605 92.805 113.895 ;
        RECT 92.975 113.775 93.305 114.155 ;
        RECT 92.550 113.435 93.300 113.605 ;
        RECT 89.160 111.775 90.030 112.115 ;
        RECT 90.620 112.155 91.420 112.325 ;
        RECT 90.200 111.605 90.450 112.065 ;
        RECT 90.620 111.865 90.790 112.155 ;
        RECT 90.970 111.605 91.300 111.985 ;
        RECT 91.640 111.605 91.945 112.745 ;
        RECT 92.115 111.915 92.370 112.795 ;
        RECT 92.550 112.615 92.900 113.265 ;
        RECT 93.070 112.445 93.300 113.435 ;
        RECT 92.550 112.275 93.300 112.445 ;
        RECT 92.550 111.775 92.805 112.275 ;
        RECT 92.975 111.605 93.305 112.105 ;
        RECT 93.475 111.775 93.645 113.895 ;
        RECT 94.005 113.795 94.335 114.155 ;
        RECT 94.505 113.765 95.000 113.935 ;
        RECT 95.205 113.765 96.060 113.935 ;
        RECT 93.875 112.575 94.335 113.625 ;
        RECT 93.815 111.790 94.140 112.575 ;
        RECT 94.505 112.405 94.675 113.765 ;
        RECT 94.845 112.855 95.195 113.475 ;
        RECT 95.365 113.255 95.720 113.475 ;
        RECT 95.365 112.665 95.535 113.255 ;
        RECT 95.890 113.055 96.060 113.765 ;
        RECT 96.935 113.695 97.265 114.155 ;
        RECT 97.475 113.795 97.825 113.965 ;
        RECT 96.265 113.225 97.055 113.475 ;
        RECT 97.475 113.405 97.735 113.795 ;
        RECT 98.045 113.705 98.995 113.985 ;
        RECT 99.165 113.715 99.355 114.155 ;
        RECT 99.525 113.775 100.595 113.945 ;
        RECT 97.225 113.055 97.395 113.235 ;
        RECT 94.505 112.235 94.900 112.405 ;
        RECT 95.070 112.275 95.535 112.665 ;
        RECT 95.705 112.885 97.395 113.055 ;
        RECT 94.730 112.105 94.900 112.235 ;
        RECT 95.705 112.105 95.875 112.885 ;
        RECT 97.565 112.715 97.735 113.405 ;
        RECT 96.235 112.545 97.735 112.715 ;
        RECT 97.925 112.745 98.135 113.535 ;
        RECT 98.305 112.915 98.655 113.535 ;
        RECT 98.825 112.925 98.995 113.705 ;
        RECT 99.525 113.545 99.695 113.775 ;
        RECT 99.165 113.375 99.695 113.545 ;
        RECT 99.165 113.095 99.385 113.375 ;
        RECT 99.865 113.205 100.105 113.605 ;
        RECT 98.825 112.755 99.230 112.925 ;
        RECT 99.565 112.835 100.105 113.205 ;
        RECT 100.275 113.420 100.595 113.775 ;
        RECT 100.840 113.695 101.145 114.155 ;
        RECT 101.315 113.445 101.570 113.975 ;
        RECT 100.275 113.245 100.600 113.420 ;
        RECT 100.275 112.945 101.190 113.245 ;
        RECT 100.450 112.915 101.190 112.945 ;
        RECT 97.925 112.585 98.600 112.745 ;
        RECT 99.060 112.665 99.230 112.755 ;
        RECT 97.925 112.575 98.890 112.585 ;
        RECT 97.565 112.405 97.735 112.545 ;
        RECT 94.310 111.605 94.560 112.065 ;
        RECT 94.730 111.775 94.980 112.105 ;
        RECT 95.195 111.775 95.875 112.105 ;
        RECT 96.045 112.205 97.120 112.375 ;
        RECT 97.565 112.235 98.125 112.405 ;
        RECT 98.430 112.285 98.890 112.575 ;
        RECT 99.060 112.495 100.280 112.665 ;
        RECT 96.045 111.865 96.215 112.205 ;
        RECT 96.450 111.605 96.780 112.035 ;
        RECT 96.950 111.865 97.120 112.205 ;
        RECT 97.415 111.605 97.785 112.065 ;
        RECT 97.955 111.775 98.125 112.235 ;
        RECT 99.060 112.115 99.230 112.495 ;
        RECT 100.450 112.325 100.620 112.915 ;
        RECT 101.360 112.795 101.570 113.445 ;
        RECT 98.360 111.775 99.230 112.115 ;
        RECT 99.820 112.155 100.620 112.325 ;
        RECT 99.400 111.605 99.650 112.065 ;
        RECT 99.820 111.865 99.990 112.155 ;
        RECT 100.170 111.605 100.500 111.985 ;
        RECT 100.840 111.605 101.145 112.745 ;
        RECT 101.315 111.915 101.570 112.795 ;
        RECT 101.745 113.480 102.005 113.985 ;
        RECT 102.185 113.775 102.515 114.155 ;
        RECT 102.695 113.605 102.865 113.985 ;
        RECT 101.745 112.680 101.915 113.480 ;
        RECT 102.200 113.435 102.865 113.605 ;
        RECT 102.200 113.180 102.370 113.435 ;
        RECT 103.185 113.335 103.395 114.155 ;
        RECT 103.565 113.355 103.895 113.985 ;
        RECT 102.085 112.850 102.370 113.180 ;
        RECT 102.605 112.885 102.935 113.255 ;
        RECT 102.200 112.705 102.370 112.850 ;
        RECT 103.565 112.755 103.815 113.355 ;
        RECT 104.065 113.335 104.295 114.155 ;
        RECT 104.505 113.385 106.175 114.155 ;
        RECT 103.985 112.915 104.315 113.165 ;
        RECT 104.505 112.865 105.255 113.385 ;
        RECT 106.845 113.335 107.075 114.155 ;
        RECT 107.245 113.355 107.575 113.985 ;
        RECT 101.745 111.775 102.015 112.680 ;
        RECT 102.200 112.535 102.865 112.705 ;
        RECT 102.185 111.605 102.515 112.365 ;
        RECT 102.695 111.775 102.865 112.535 ;
        RECT 103.185 111.605 103.395 112.745 ;
        RECT 103.565 111.775 103.895 112.755 ;
        RECT 104.065 111.605 104.295 112.745 ;
        RECT 105.425 112.695 106.175 113.215 ;
        RECT 106.825 112.915 107.155 113.165 ;
        RECT 107.325 112.755 107.575 113.355 ;
        RECT 107.745 113.335 107.955 114.155 ;
        RECT 108.645 113.430 108.935 114.155 ;
        RECT 109.105 113.385 111.695 114.155 ;
        RECT 112.325 113.405 113.535 114.155 ;
        RECT 109.105 112.865 110.315 113.385 ;
        RECT 104.505 111.605 106.175 112.695 ;
        RECT 106.845 111.605 107.075 112.745 ;
        RECT 107.245 111.775 107.575 112.755 ;
        RECT 107.745 111.605 107.955 112.745 ;
        RECT 108.645 111.605 108.935 112.770 ;
        RECT 110.485 112.695 111.695 113.215 ;
        RECT 109.105 111.605 111.695 112.695 ;
        RECT 112.325 112.695 112.845 113.235 ;
        RECT 113.015 112.865 113.535 113.405 ;
        RECT 112.325 111.605 113.535 112.695 ;
        RECT 5.520 111.435 113.620 111.605 ;
        RECT 5.605 110.345 6.815 111.435 ;
        RECT 6.985 110.345 8.195 111.435 ;
        RECT 5.605 109.635 6.125 110.175 ;
        RECT 6.295 109.805 6.815 110.345 ;
        RECT 6.985 109.635 7.505 110.175 ;
        RECT 7.675 109.805 8.195 110.345 ;
        RECT 8.370 110.245 8.625 111.125 ;
        RECT 8.795 110.295 9.100 111.435 ;
        RECT 9.440 111.055 9.770 111.435 ;
        RECT 9.950 110.885 10.120 111.175 ;
        RECT 10.290 110.975 10.540 111.435 ;
        RECT 9.320 110.715 10.120 110.885 ;
        RECT 10.710 110.925 11.580 111.265 ;
        RECT 5.605 108.885 6.815 109.635 ;
        RECT 6.985 108.885 8.195 109.635 ;
        RECT 8.370 109.595 8.580 110.245 ;
        RECT 9.320 110.125 9.490 110.715 ;
        RECT 10.710 110.545 10.880 110.925 ;
        RECT 11.815 110.805 11.985 111.265 ;
        RECT 12.155 110.975 12.525 111.435 ;
        RECT 12.820 110.835 12.990 111.175 ;
        RECT 13.160 111.005 13.490 111.435 ;
        RECT 13.725 110.835 13.895 111.175 ;
        RECT 9.660 110.375 10.880 110.545 ;
        RECT 11.050 110.465 11.510 110.755 ;
        RECT 11.815 110.635 12.375 110.805 ;
        RECT 12.820 110.665 13.895 110.835 ;
        RECT 14.065 110.935 14.745 111.265 ;
        RECT 14.960 110.935 15.210 111.265 ;
        RECT 15.380 110.975 15.630 111.435 ;
        RECT 12.205 110.495 12.375 110.635 ;
        RECT 11.050 110.455 12.015 110.465 ;
        RECT 10.710 110.285 10.880 110.375 ;
        RECT 11.340 110.295 12.015 110.455 ;
        RECT 8.750 110.095 9.490 110.125 ;
        RECT 8.750 109.795 9.665 110.095 ;
        RECT 9.340 109.620 9.665 109.795 ;
        RECT 8.370 109.065 8.625 109.595 ;
        RECT 8.795 108.885 9.100 109.345 ;
        RECT 9.345 109.265 9.665 109.620 ;
        RECT 9.835 109.835 10.375 110.205 ;
        RECT 10.710 110.115 11.115 110.285 ;
        RECT 9.835 109.435 10.075 109.835 ;
        RECT 10.555 109.665 10.775 109.945 ;
        RECT 10.245 109.495 10.775 109.665 ;
        RECT 10.245 109.265 10.415 109.495 ;
        RECT 10.945 109.335 11.115 110.115 ;
        RECT 11.285 109.505 11.635 110.125 ;
        RECT 11.805 109.505 12.015 110.295 ;
        RECT 12.205 110.325 13.705 110.495 ;
        RECT 12.205 109.635 12.375 110.325 ;
        RECT 14.065 110.155 14.235 110.935 ;
        RECT 15.040 110.805 15.210 110.935 ;
        RECT 12.545 109.985 14.235 110.155 ;
        RECT 14.405 110.375 14.870 110.765 ;
        RECT 15.040 110.635 15.435 110.805 ;
        RECT 12.545 109.805 12.715 109.985 ;
        RECT 9.345 109.095 10.415 109.265 ;
        RECT 10.585 108.885 10.775 109.325 ;
        RECT 10.945 109.055 11.895 109.335 ;
        RECT 12.205 109.245 12.465 109.635 ;
        RECT 12.885 109.565 13.675 109.815 ;
        RECT 12.115 109.075 12.465 109.245 ;
        RECT 12.675 108.885 13.005 109.345 ;
        RECT 13.880 109.275 14.050 109.985 ;
        RECT 14.405 109.785 14.575 110.375 ;
        RECT 14.220 109.565 14.575 109.785 ;
        RECT 14.745 109.565 15.095 110.185 ;
        RECT 15.265 109.275 15.435 110.635 ;
        RECT 15.800 110.465 16.125 111.250 ;
        RECT 15.605 109.415 16.065 110.465 ;
        RECT 13.880 109.105 14.735 109.275 ;
        RECT 14.940 109.105 15.435 109.275 ;
        RECT 15.605 108.885 15.935 109.245 ;
        RECT 16.295 109.145 16.465 111.265 ;
        RECT 16.635 110.935 16.965 111.435 ;
        RECT 17.135 110.765 17.390 111.265 ;
        RECT 16.640 110.595 17.390 110.765 ;
        RECT 16.640 109.605 16.870 110.595 ;
        RECT 17.040 109.775 17.390 110.425 ;
        RECT 18.485 110.270 18.775 111.435 ;
        RECT 19.870 110.245 20.125 111.125 ;
        RECT 20.295 110.295 20.600 111.435 ;
        RECT 20.940 111.055 21.270 111.435 ;
        RECT 21.450 110.885 21.620 111.175 ;
        RECT 21.790 110.975 22.040 111.435 ;
        RECT 20.820 110.715 21.620 110.885 ;
        RECT 22.210 110.925 23.080 111.265 ;
        RECT 16.640 109.435 17.390 109.605 ;
        RECT 16.635 108.885 16.965 109.265 ;
        RECT 17.135 109.145 17.390 109.435 ;
        RECT 18.485 108.885 18.775 109.610 ;
        RECT 19.870 109.595 20.080 110.245 ;
        RECT 20.820 110.125 20.990 110.715 ;
        RECT 22.210 110.545 22.380 110.925 ;
        RECT 23.315 110.805 23.485 111.265 ;
        RECT 23.655 110.975 24.025 111.435 ;
        RECT 24.320 110.835 24.490 111.175 ;
        RECT 24.660 111.005 24.990 111.435 ;
        RECT 25.225 110.835 25.395 111.175 ;
        RECT 21.160 110.375 22.380 110.545 ;
        RECT 22.550 110.465 23.010 110.755 ;
        RECT 23.315 110.635 23.875 110.805 ;
        RECT 24.320 110.665 25.395 110.835 ;
        RECT 25.565 110.935 26.245 111.265 ;
        RECT 26.460 110.935 26.710 111.265 ;
        RECT 26.880 110.975 27.130 111.435 ;
        RECT 23.705 110.495 23.875 110.635 ;
        RECT 22.550 110.455 23.515 110.465 ;
        RECT 22.210 110.285 22.380 110.375 ;
        RECT 22.840 110.295 23.515 110.455 ;
        RECT 20.250 110.095 20.990 110.125 ;
        RECT 20.250 109.795 21.165 110.095 ;
        RECT 20.840 109.620 21.165 109.795 ;
        RECT 19.870 109.065 20.125 109.595 ;
        RECT 20.295 108.885 20.600 109.345 ;
        RECT 20.845 109.265 21.165 109.620 ;
        RECT 21.335 109.835 21.875 110.205 ;
        RECT 22.210 110.115 22.615 110.285 ;
        RECT 21.335 109.435 21.575 109.835 ;
        RECT 22.055 109.665 22.275 109.945 ;
        RECT 21.745 109.495 22.275 109.665 ;
        RECT 21.745 109.265 21.915 109.495 ;
        RECT 22.445 109.335 22.615 110.115 ;
        RECT 22.785 109.505 23.135 110.125 ;
        RECT 23.305 109.505 23.515 110.295 ;
        RECT 23.705 110.325 25.205 110.495 ;
        RECT 23.705 109.635 23.875 110.325 ;
        RECT 25.565 110.155 25.735 110.935 ;
        RECT 26.540 110.805 26.710 110.935 ;
        RECT 24.045 109.985 25.735 110.155 ;
        RECT 25.905 110.375 26.370 110.765 ;
        RECT 26.540 110.635 26.935 110.805 ;
        RECT 24.045 109.805 24.215 109.985 ;
        RECT 20.845 109.095 21.915 109.265 ;
        RECT 22.085 108.885 22.275 109.325 ;
        RECT 22.445 109.055 23.395 109.335 ;
        RECT 23.705 109.245 23.965 109.635 ;
        RECT 24.385 109.565 25.175 109.815 ;
        RECT 23.615 109.075 23.965 109.245 ;
        RECT 24.175 108.885 24.505 109.345 ;
        RECT 25.380 109.275 25.550 109.985 ;
        RECT 25.905 109.785 26.075 110.375 ;
        RECT 25.720 109.565 26.075 109.785 ;
        RECT 26.245 109.565 26.595 110.185 ;
        RECT 26.765 109.275 26.935 110.635 ;
        RECT 27.300 110.465 27.625 111.250 ;
        RECT 27.105 109.415 27.565 110.465 ;
        RECT 25.380 109.105 26.235 109.275 ;
        RECT 26.440 109.105 26.935 109.275 ;
        RECT 27.105 108.885 27.435 109.245 ;
        RECT 27.795 109.145 27.965 111.265 ;
        RECT 28.135 110.935 28.465 111.435 ;
        RECT 28.635 110.765 28.890 111.265 ;
        RECT 28.140 110.595 28.890 110.765 ;
        RECT 28.140 109.605 28.370 110.595 ;
        RECT 28.540 109.775 28.890 110.425 ;
        RECT 29.125 110.295 29.335 111.435 ;
        RECT 29.505 110.285 29.835 111.265 ;
        RECT 30.005 110.295 30.235 111.435 ;
        RECT 30.445 110.345 31.655 111.435 ;
        RECT 28.140 109.435 28.890 109.605 ;
        RECT 28.135 108.885 28.465 109.265 ;
        RECT 28.635 109.145 28.890 109.435 ;
        RECT 29.125 108.885 29.335 109.705 ;
        RECT 29.505 109.685 29.755 110.285 ;
        RECT 29.925 109.875 30.255 110.125 ;
        RECT 29.505 109.055 29.835 109.685 ;
        RECT 30.005 108.885 30.235 109.705 ;
        RECT 30.445 109.635 30.965 110.175 ;
        RECT 31.135 109.805 31.655 110.345 ;
        RECT 31.915 110.505 32.085 111.265 ;
        RECT 32.265 110.675 32.595 111.435 ;
        RECT 31.915 110.335 32.580 110.505 ;
        RECT 32.765 110.360 33.035 111.265 ;
        RECT 32.410 110.190 32.580 110.335 ;
        RECT 31.845 109.785 32.175 110.155 ;
        RECT 32.410 109.860 32.695 110.190 ;
        RECT 30.445 108.885 31.655 109.635 ;
        RECT 32.410 109.605 32.580 109.860 ;
        RECT 31.915 109.435 32.580 109.605 ;
        RECT 32.865 109.560 33.035 110.360 ;
        RECT 33.245 110.295 33.475 111.435 ;
        RECT 33.645 110.285 33.975 111.265 ;
        RECT 34.145 110.295 34.355 111.435 ;
        RECT 34.590 110.765 34.845 111.265 ;
        RECT 35.015 110.935 35.345 111.435 ;
        RECT 34.590 110.595 35.340 110.765 ;
        RECT 33.225 109.875 33.555 110.125 ;
        RECT 31.915 109.055 32.085 109.435 ;
        RECT 32.265 108.885 32.595 109.265 ;
        RECT 32.775 109.055 33.035 109.560 ;
        RECT 33.245 108.885 33.475 109.705 ;
        RECT 33.725 109.685 33.975 110.285 ;
        RECT 34.590 109.775 34.940 110.425 ;
        RECT 33.645 109.055 33.975 109.685 ;
        RECT 34.145 108.885 34.355 109.705 ;
        RECT 35.110 109.605 35.340 110.595 ;
        RECT 34.590 109.435 35.340 109.605 ;
        RECT 34.590 109.145 34.845 109.435 ;
        RECT 35.015 108.885 35.345 109.265 ;
        RECT 35.515 109.145 35.685 111.265 ;
        RECT 35.855 110.465 36.180 111.250 ;
        RECT 36.350 110.975 36.600 111.435 ;
        RECT 36.770 110.935 37.020 111.265 ;
        RECT 37.235 110.935 37.915 111.265 ;
        RECT 36.770 110.805 36.940 110.935 ;
        RECT 36.545 110.635 36.940 110.805 ;
        RECT 35.915 109.415 36.375 110.465 ;
        RECT 36.545 109.275 36.715 110.635 ;
        RECT 37.110 110.375 37.575 110.765 ;
        RECT 36.885 109.565 37.235 110.185 ;
        RECT 37.405 109.785 37.575 110.375 ;
        RECT 37.745 110.155 37.915 110.935 ;
        RECT 38.085 110.835 38.255 111.175 ;
        RECT 38.490 111.005 38.820 111.435 ;
        RECT 38.990 110.835 39.160 111.175 ;
        RECT 39.455 110.975 39.825 111.435 ;
        RECT 38.085 110.665 39.160 110.835 ;
        RECT 39.995 110.805 40.165 111.265 ;
        RECT 40.400 110.925 41.270 111.265 ;
        RECT 41.440 110.975 41.690 111.435 ;
        RECT 39.605 110.635 40.165 110.805 ;
        RECT 39.605 110.495 39.775 110.635 ;
        RECT 38.275 110.325 39.775 110.495 ;
        RECT 40.470 110.465 40.930 110.755 ;
        RECT 37.745 109.985 39.435 110.155 ;
        RECT 37.405 109.565 37.760 109.785 ;
        RECT 37.930 109.275 38.100 109.985 ;
        RECT 38.305 109.565 39.095 109.815 ;
        RECT 39.265 109.805 39.435 109.985 ;
        RECT 39.605 109.635 39.775 110.325 ;
        RECT 36.045 108.885 36.375 109.245 ;
        RECT 36.545 109.105 37.040 109.275 ;
        RECT 37.245 109.105 38.100 109.275 ;
        RECT 38.975 108.885 39.305 109.345 ;
        RECT 39.515 109.245 39.775 109.635 ;
        RECT 39.965 110.455 40.930 110.465 ;
        RECT 41.100 110.545 41.270 110.925 ;
        RECT 41.860 110.885 42.030 111.175 ;
        RECT 42.210 111.055 42.540 111.435 ;
        RECT 41.860 110.715 42.660 110.885 ;
        RECT 39.965 110.295 40.640 110.455 ;
        RECT 41.100 110.375 42.320 110.545 ;
        RECT 39.965 109.505 40.175 110.295 ;
        RECT 41.100 110.285 41.270 110.375 ;
        RECT 40.345 109.505 40.695 110.125 ;
        RECT 40.865 110.115 41.270 110.285 ;
        RECT 40.865 109.335 41.035 110.115 ;
        RECT 41.205 109.665 41.425 109.945 ;
        RECT 41.605 109.835 42.145 110.205 ;
        RECT 42.490 110.125 42.660 110.715 ;
        RECT 42.880 110.295 43.185 111.435 ;
        RECT 43.355 110.245 43.610 111.125 ;
        RECT 44.245 110.270 44.535 111.435 ;
        RECT 45.715 110.505 45.885 111.265 ;
        RECT 46.065 110.675 46.395 111.435 ;
        RECT 45.715 110.335 46.380 110.505 ;
        RECT 46.565 110.360 46.835 111.265 ;
        RECT 47.010 110.765 47.265 111.265 ;
        RECT 47.435 110.935 47.765 111.435 ;
        RECT 47.010 110.595 47.760 110.765 ;
        RECT 42.490 110.095 43.230 110.125 ;
        RECT 41.205 109.495 41.735 109.665 ;
        RECT 39.515 109.075 39.865 109.245 ;
        RECT 40.085 109.055 41.035 109.335 ;
        RECT 41.205 108.885 41.395 109.325 ;
        RECT 41.565 109.265 41.735 109.495 ;
        RECT 41.905 109.435 42.145 109.835 ;
        RECT 42.315 109.795 43.230 110.095 ;
        RECT 42.315 109.620 42.640 109.795 ;
        RECT 42.315 109.265 42.635 109.620 ;
        RECT 43.400 109.595 43.610 110.245 ;
        RECT 46.210 110.190 46.380 110.335 ;
        RECT 45.645 109.785 45.975 110.155 ;
        RECT 46.210 109.860 46.495 110.190 ;
        RECT 41.565 109.095 42.635 109.265 ;
        RECT 42.880 108.885 43.185 109.345 ;
        RECT 43.355 109.065 43.610 109.595 ;
        RECT 44.245 108.885 44.535 109.610 ;
        RECT 46.210 109.605 46.380 109.860 ;
        RECT 45.715 109.435 46.380 109.605 ;
        RECT 46.665 109.560 46.835 110.360 ;
        RECT 47.010 109.775 47.360 110.425 ;
        RECT 47.530 109.605 47.760 110.595 ;
        RECT 45.715 109.055 45.885 109.435 ;
        RECT 46.065 108.885 46.395 109.265 ;
        RECT 46.575 109.055 46.835 109.560 ;
        RECT 47.010 109.435 47.760 109.605 ;
        RECT 47.010 109.145 47.265 109.435 ;
        RECT 47.435 108.885 47.765 109.265 ;
        RECT 47.935 109.145 48.105 111.265 ;
        RECT 48.275 110.465 48.600 111.250 ;
        RECT 48.770 110.975 49.020 111.435 ;
        RECT 49.190 110.935 49.440 111.265 ;
        RECT 49.655 110.935 50.335 111.265 ;
        RECT 49.190 110.805 49.360 110.935 ;
        RECT 48.965 110.635 49.360 110.805 ;
        RECT 48.335 109.415 48.795 110.465 ;
        RECT 48.965 109.275 49.135 110.635 ;
        RECT 49.530 110.375 49.995 110.765 ;
        RECT 49.305 109.565 49.655 110.185 ;
        RECT 49.825 109.785 49.995 110.375 ;
        RECT 50.165 110.155 50.335 110.935 ;
        RECT 50.505 110.835 50.675 111.175 ;
        RECT 50.910 111.005 51.240 111.435 ;
        RECT 51.410 110.835 51.580 111.175 ;
        RECT 51.875 110.975 52.245 111.435 ;
        RECT 50.505 110.665 51.580 110.835 ;
        RECT 52.415 110.805 52.585 111.265 ;
        RECT 52.820 110.925 53.690 111.265 ;
        RECT 53.860 110.975 54.110 111.435 ;
        RECT 52.025 110.635 52.585 110.805 ;
        RECT 52.025 110.495 52.195 110.635 ;
        RECT 50.695 110.325 52.195 110.495 ;
        RECT 52.890 110.465 53.350 110.755 ;
        RECT 50.165 109.985 51.855 110.155 ;
        RECT 49.825 109.565 50.180 109.785 ;
        RECT 50.350 109.275 50.520 109.985 ;
        RECT 50.725 109.565 51.515 109.815 ;
        RECT 51.685 109.805 51.855 109.985 ;
        RECT 52.025 109.635 52.195 110.325 ;
        RECT 48.465 108.885 48.795 109.245 ;
        RECT 48.965 109.105 49.460 109.275 ;
        RECT 49.665 109.105 50.520 109.275 ;
        RECT 51.395 108.885 51.725 109.345 ;
        RECT 51.935 109.245 52.195 109.635 ;
        RECT 52.385 110.455 53.350 110.465 ;
        RECT 53.520 110.545 53.690 110.925 ;
        RECT 54.280 110.885 54.450 111.175 ;
        RECT 54.630 111.055 54.960 111.435 ;
        RECT 54.280 110.715 55.080 110.885 ;
        RECT 52.385 110.295 53.060 110.455 ;
        RECT 53.520 110.375 54.740 110.545 ;
        RECT 52.385 109.505 52.595 110.295 ;
        RECT 53.520 110.285 53.690 110.375 ;
        RECT 52.765 109.505 53.115 110.125 ;
        RECT 53.285 110.115 53.690 110.285 ;
        RECT 53.285 109.335 53.455 110.115 ;
        RECT 53.625 109.665 53.845 109.945 ;
        RECT 54.025 109.835 54.565 110.205 ;
        RECT 54.910 110.125 55.080 110.715 ;
        RECT 55.300 110.295 55.605 111.435 ;
        RECT 55.775 110.245 56.030 111.125 ;
        RECT 56.245 110.295 56.475 111.435 ;
        RECT 56.645 110.285 56.975 111.265 ;
        RECT 57.145 110.295 57.355 111.435 ;
        RECT 57.585 110.345 58.795 111.435 ;
        RECT 58.970 110.765 59.225 111.265 ;
        RECT 59.395 110.935 59.725 111.435 ;
        RECT 58.970 110.595 59.720 110.765 ;
        RECT 54.910 110.095 55.650 110.125 ;
        RECT 53.625 109.495 54.155 109.665 ;
        RECT 51.935 109.075 52.285 109.245 ;
        RECT 52.505 109.055 53.455 109.335 ;
        RECT 53.625 108.885 53.815 109.325 ;
        RECT 53.985 109.265 54.155 109.495 ;
        RECT 54.325 109.435 54.565 109.835 ;
        RECT 54.735 109.795 55.650 110.095 ;
        RECT 54.735 109.620 55.060 109.795 ;
        RECT 54.735 109.265 55.055 109.620 ;
        RECT 55.820 109.595 56.030 110.245 ;
        RECT 56.225 109.875 56.555 110.125 ;
        RECT 53.985 109.095 55.055 109.265 ;
        RECT 55.300 108.885 55.605 109.345 ;
        RECT 55.775 109.065 56.030 109.595 ;
        RECT 56.245 108.885 56.475 109.705 ;
        RECT 56.725 109.685 56.975 110.285 ;
        RECT 56.645 109.055 56.975 109.685 ;
        RECT 57.145 108.885 57.355 109.705 ;
        RECT 57.585 109.635 58.105 110.175 ;
        RECT 58.275 109.805 58.795 110.345 ;
        RECT 58.970 109.775 59.320 110.425 ;
        RECT 57.585 108.885 58.795 109.635 ;
        RECT 59.490 109.605 59.720 110.595 ;
        RECT 58.970 109.435 59.720 109.605 ;
        RECT 58.970 109.145 59.225 109.435 ;
        RECT 59.395 108.885 59.725 109.265 ;
        RECT 59.895 109.145 60.065 111.265 ;
        RECT 60.235 110.465 60.560 111.250 ;
        RECT 60.730 110.975 60.980 111.435 ;
        RECT 61.150 110.935 61.400 111.265 ;
        RECT 61.615 110.935 62.295 111.265 ;
        RECT 61.150 110.805 61.320 110.935 ;
        RECT 60.925 110.635 61.320 110.805 ;
        RECT 60.295 109.415 60.755 110.465 ;
        RECT 60.925 109.275 61.095 110.635 ;
        RECT 61.490 110.375 61.955 110.765 ;
        RECT 61.265 109.565 61.615 110.185 ;
        RECT 61.785 109.785 61.955 110.375 ;
        RECT 62.125 110.155 62.295 110.935 ;
        RECT 62.465 110.835 62.635 111.175 ;
        RECT 62.870 111.005 63.200 111.435 ;
        RECT 63.370 110.835 63.540 111.175 ;
        RECT 63.835 110.975 64.205 111.435 ;
        RECT 62.465 110.665 63.540 110.835 ;
        RECT 64.375 110.805 64.545 111.265 ;
        RECT 64.780 110.925 65.650 111.265 ;
        RECT 65.820 110.975 66.070 111.435 ;
        RECT 63.985 110.635 64.545 110.805 ;
        RECT 63.985 110.495 64.155 110.635 ;
        RECT 62.655 110.325 64.155 110.495 ;
        RECT 64.850 110.465 65.310 110.755 ;
        RECT 62.125 109.985 63.815 110.155 ;
        RECT 61.785 109.565 62.140 109.785 ;
        RECT 62.310 109.275 62.480 109.985 ;
        RECT 62.685 109.565 63.475 109.815 ;
        RECT 63.645 109.805 63.815 109.985 ;
        RECT 63.985 109.635 64.155 110.325 ;
        RECT 60.425 108.885 60.755 109.245 ;
        RECT 60.925 109.105 61.420 109.275 ;
        RECT 61.625 109.105 62.480 109.275 ;
        RECT 63.355 108.885 63.685 109.345 ;
        RECT 63.895 109.245 64.155 109.635 ;
        RECT 64.345 110.455 65.310 110.465 ;
        RECT 65.480 110.545 65.650 110.925 ;
        RECT 66.240 110.885 66.410 111.175 ;
        RECT 66.590 111.055 66.920 111.435 ;
        RECT 66.240 110.715 67.040 110.885 ;
        RECT 64.345 110.295 65.020 110.455 ;
        RECT 65.480 110.375 66.700 110.545 ;
        RECT 64.345 109.505 64.555 110.295 ;
        RECT 65.480 110.285 65.650 110.375 ;
        RECT 64.725 109.505 65.075 110.125 ;
        RECT 65.245 110.115 65.650 110.285 ;
        RECT 65.245 109.335 65.415 110.115 ;
        RECT 65.585 109.665 65.805 109.945 ;
        RECT 65.985 109.835 66.525 110.205 ;
        RECT 66.870 110.125 67.040 110.715 ;
        RECT 67.260 110.295 67.565 111.435 ;
        RECT 67.735 110.245 67.990 111.125 ;
        RECT 66.870 110.095 67.610 110.125 ;
        RECT 65.585 109.495 66.115 109.665 ;
        RECT 63.895 109.075 64.245 109.245 ;
        RECT 64.465 109.055 65.415 109.335 ;
        RECT 65.585 108.885 65.775 109.325 ;
        RECT 65.945 109.265 66.115 109.495 ;
        RECT 66.285 109.435 66.525 109.835 ;
        RECT 66.695 109.795 67.610 110.095 ;
        RECT 66.695 109.620 67.020 109.795 ;
        RECT 66.695 109.265 67.015 109.620 ;
        RECT 67.780 109.595 67.990 110.245 ;
        RECT 65.945 109.095 67.015 109.265 ;
        RECT 67.260 108.885 67.565 109.345 ;
        RECT 67.735 109.065 67.990 109.595 ;
        RECT 68.165 110.360 68.435 111.265 ;
        RECT 68.605 110.675 68.935 111.435 ;
        RECT 69.115 110.505 69.285 111.265 ;
        RECT 68.165 109.560 68.335 110.360 ;
        RECT 68.620 110.335 69.285 110.505 ;
        RECT 68.620 110.190 68.790 110.335 ;
        RECT 70.005 110.270 70.295 111.435 ;
        RECT 70.525 110.295 70.735 111.435 ;
        RECT 70.905 110.285 71.235 111.265 ;
        RECT 71.405 110.295 71.635 111.435 ;
        RECT 72.765 110.360 73.035 111.265 ;
        RECT 73.205 110.675 73.535 111.435 ;
        RECT 73.715 110.505 73.885 111.265 ;
        RECT 74.150 110.765 74.405 111.265 ;
        RECT 74.575 110.935 74.905 111.435 ;
        RECT 74.150 110.595 74.900 110.765 ;
        RECT 68.505 109.860 68.790 110.190 ;
        RECT 68.620 109.605 68.790 109.860 ;
        RECT 69.025 109.785 69.355 110.155 ;
        RECT 68.165 109.055 68.425 109.560 ;
        RECT 68.620 109.435 69.285 109.605 ;
        RECT 68.605 108.885 68.935 109.265 ;
        RECT 69.115 109.055 69.285 109.435 ;
        RECT 70.005 108.885 70.295 109.610 ;
        RECT 70.525 108.885 70.735 109.705 ;
        RECT 70.905 109.685 71.155 110.285 ;
        RECT 71.325 109.875 71.655 110.125 ;
        RECT 70.905 109.055 71.235 109.685 ;
        RECT 71.405 108.885 71.635 109.705 ;
        RECT 72.765 109.560 72.935 110.360 ;
        RECT 73.220 110.335 73.885 110.505 ;
        RECT 73.220 110.190 73.390 110.335 ;
        RECT 73.105 109.860 73.390 110.190 ;
        RECT 73.220 109.605 73.390 109.860 ;
        RECT 73.625 109.785 73.955 110.155 ;
        RECT 74.150 109.775 74.500 110.425 ;
        RECT 74.670 109.605 74.900 110.595 ;
        RECT 72.765 109.055 73.025 109.560 ;
        RECT 73.220 109.435 73.885 109.605 ;
        RECT 73.205 108.885 73.535 109.265 ;
        RECT 73.715 109.055 73.885 109.435 ;
        RECT 74.150 109.435 74.900 109.605 ;
        RECT 74.150 109.145 74.405 109.435 ;
        RECT 74.575 108.885 74.905 109.265 ;
        RECT 75.075 109.145 75.245 111.265 ;
        RECT 75.415 110.465 75.740 111.250 ;
        RECT 75.910 110.975 76.160 111.435 ;
        RECT 76.330 110.935 76.580 111.265 ;
        RECT 76.795 110.935 77.475 111.265 ;
        RECT 76.330 110.805 76.500 110.935 ;
        RECT 76.105 110.635 76.500 110.805 ;
        RECT 75.475 109.415 75.935 110.465 ;
        RECT 76.105 109.275 76.275 110.635 ;
        RECT 76.670 110.375 77.135 110.765 ;
        RECT 76.445 109.565 76.795 110.185 ;
        RECT 76.965 109.785 77.135 110.375 ;
        RECT 77.305 110.155 77.475 110.935 ;
        RECT 77.645 110.835 77.815 111.175 ;
        RECT 78.050 111.005 78.380 111.435 ;
        RECT 78.550 110.835 78.720 111.175 ;
        RECT 79.015 110.975 79.385 111.435 ;
        RECT 77.645 110.665 78.720 110.835 ;
        RECT 79.555 110.805 79.725 111.265 ;
        RECT 79.960 110.925 80.830 111.265 ;
        RECT 81.000 110.975 81.250 111.435 ;
        RECT 79.165 110.635 79.725 110.805 ;
        RECT 79.165 110.495 79.335 110.635 ;
        RECT 77.835 110.325 79.335 110.495 ;
        RECT 80.030 110.465 80.490 110.755 ;
        RECT 77.305 109.985 78.995 110.155 ;
        RECT 76.965 109.565 77.320 109.785 ;
        RECT 77.490 109.275 77.660 109.985 ;
        RECT 77.865 109.565 78.655 109.815 ;
        RECT 78.825 109.805 78.995 109.985 ;
        RECT 79.165 109.635 79.335 110.325 ;
        RECT 75.605 108.885 75.935 109.245 ;
        RECT 76.105 109.105 76.600 109.275 ;
        RECT 76.805 109.105 77.660 109.275 ;
        RECT 78.535 108.885 78.865 109.345 ;
        RECT 79.075 109.245 79.335 109.635 ;
        RECT 79.525 110.455 80.490 110.465 ;
        RECT 80.660 110.545 80.830 110.925 ;
        RECT 81.420 110.885 81.590 111.175 ;
        RECT 81.770 111.055 82.100 111.435 ;
        RECT 81.420 110.715 82.220 110.885 ;
        RECT 79.525 110.295 80.200 110.455 ;
        RECT 80.660 110.375 81.880 110.545 ;
        RECT 79.525 109.505 79.735 110.295 ;
        RECT 80.660 110.285 80.830 110.375 ;
        RECT 79.905 109.505 80.255 110.125 ;
        RECT 80.425 110.115 80.830 110.285 ;
        RECT 80.425 109.335 80.595 110.115 ;
        RECT 80.765 109.665 80.985 109.945 ;
        RECT 81.165 109.835 81.705 110.205 ;
        RECT 82.050 110.125 82.220 110.715 ;
        RECT 82.440 110.295 82.745 111.435 ;
        RECT 82.915 110.245 83.170 111.125 ;
        RECT 83.435 110.505 83.605 111.265 ;
        RECT 83.785 110.675 84.115 111.435 ;
        RECT 83.435 110.335 84.100 110.505 ;
        RECT 84.285 110.360 84.555 111.265 ;
        RECT 85.650 110.765 85.905 111.265 ;
        RECT 86.075 110.935 86.405 111.435 ;
        RECT 85.650 110.595 86.400 110.765 ;
        RECT 82.050 110.095 82.790 110.125 ;
        RECT 80.765 109.495 81.295 109.665 ;
        RECT 79.075 109.075 79.425 109.245 ;
        RECT 79.645 109.055 80.595 109.335 ;
        RECT 80.765 108.885 80.955 109.325 ;
        RECT 81.125 109.265 81.295 109.495 ;
        RECT 81.465 109.435 81.705 109.835 ;
        RECT 81.875 109.795 82.790 110.095 ;
        RECT 81.875 109.620 82.200 109.795 ;
        RECT 81.875 109.265 82.195 109.620 ;
        RECT 82.960 109.595 83.170 110.245 ;
        RECT 83.930 110.190 84.100 110.335 ;
        RECT 83.365 109.785 83.695 110.155 ;
        RECT 83.930 109.860 84.215 110.190 ;
        RECT 83.930 109.605 84.100 109.860 ;
        RECT 81.125 109.095 82.195 109.265 ;
        RECT 82.440 108.885 82.745 109.345 ;
        RECT 82.915 109.065 83.170 109.595 ;
        RECT 83.435 109.435 84.100 109.605 ;
        RECT 84.385 109.560 84.555 110.360 ;
        RECT 85.650 109.775 86.000 110.425 ;
        RECT 86.170 109.605 86.400 110.595 ;
        RECT 83.435 109.055 83.605 109.435 ;
        RECT 83.785 108.885 84.115 109.265 ;
        RECT 84.295 109.055 84.555 109.560 ;
        RECT 85.650 109.435 86.400 109.605 ;
        RECT 85.650 109.145 85.905 109.435 ;
        RECT 86.075 108.885 86.405 109.265 ;
        RECT 86.575 109.145 86.745 111.265 ;
        RECT 86.915 110.465 87.240 111.250 ;
        RECT 87.410 110.975 87.660 111.435 ;
        RECT 87.830 110.935 88.080 111.265 ;
        RECT 88.295 110.935 88.975 111.265 ;
        RECT 87.830 110.805 88.000 110.935 ;
        RECT 87.605 110.635 88.000 110.805 ;
        RECT 86.975 109.415 87.435 110.465 ;
        RECT 87.605 109.275 87.775 110.635 ;
        RECT 88.170 110.375 88.635 110.765 ;
        RECT 87.945 109.565 88.295 110.185 ;
        RECT 88.465 109.785 88.635 110.375 ;
        RECT 88.805 110.155 88.975 110.935 ;
        RECT 89.145 110.835 89.315 111.175 ;
        RECT 89.550 111.005 89.880 111.435 ;
        RECT 90.050 110.835 90.220 111.175 ;
        RECT 90.515 110.975 90.885 111.435 ;
        RECT 89.145 110.665 90.220 110.835 ;
        RECT 91.055 110.805 91.225 111.265 ;
        RECT 91.460 110.925 92.330 111.265 ;
        RECT 92.500 110.975 92.750 111.435 ;
        RECT 90.665 110.635 91.225 110.805 ;
        RECT 90.665 110.495 90.835 110.635 ;
        RECT 89.335 110.325 90.835 110.495 ;
        RECT 91.530 110.465 91.990 110.755 ;
        RECT 88.805 109.985 90.495 110.155 ;
        RECT 88.465 109.565 88.820 109.785 ;
        RECT 88.990 109.275 89.160 109.985 ;
        RECT 89.365 109.565 90.155 109.815 ;
        RECT 90.325 109.805 90.495 109.985 ;
        RECT 90.665 109.635 90.835 110.325 ;
        RECT 87.105 108.885 87.435 109.245 ;
        RECT 87.605 109.105 88.100 109.275 ;
        RECT 88.305 109.105 89.160 109.275 ;
        RECT 90.035 108.885 90.365 109.345 ;
        RECT 90.575 109.245 90.835 109.635 ;
        RECT 91.025 110.455 91.990 110.465 ;
        RECT 92.160 110.545 92.330 110.925 ;
        RECT 92.920 110.885 93.090 111.175 ;
        RECT 93.270 111.055 93.600 111.435 ;
        RECT 92.920 110.715 93.720 110.885 ;
        RECT 91.025 110.295 91.700 110.455 ;
        RECT 92.160 110.375 93.380 110.545 ;
        RECT 91.025 109.505 91.235 110.295 ;
        RECT 92.160 110.285 92.330 110.375 ;
        RECT 91.405 109.505 91.755 110.125 ;
        RECT 91.925 110.115 92.330 110.285 ;
        RECT 91.925 109.335 92.095 110.115 ;
        RECT 92.265 109.665 92.485 109.945 ;
        RECT 92.665 109.835 93.205 110.205 ;
        RECT 93.550 110.125 93.720 110.715 ;
        RECT 93.940 110.295 94.245 111.435 ;
        RECT 94.415 110.245 94.670 111.125 ;
        RECT 95.765 110.270 96.055 111.435 ;
        RECT 96.225 110.360 96.495 111.265 ;
        RECT 96.665 110.675 96.995 111.435 ;
        RECT 97.175 110.505 97.345 111.265 ;
        RECT 97.610 110.765 97.865 111.265 ;
        RECT 98.035 110.935 98.365 111.435 ;
        RECT 97.610 110.595 98.360 110.765 ;
        RECT 93.550 110.095 94.290 110.125 ;
        RECT 92.265 109.495 92.795 109.665 ;
        RECT 90.575 109.075 90.925 109.245 ;
        RECT 91.145 109.055 92.095 109.335 ;
        RECT 92.265 108.885 92.455 109.325 ;
        RECT 92.625 109.265 92.795 109.495 ;
        RECT 92.965 109.435 93.205 109.835 ;
        RECT 93.375 109.795 94.290 110.095 ;
        RECT 93.375 109.620 93.700 109.795 ;
        RECT 93.375 109.265 93.695 109.620 ;
        RECT 94.460 109.595 94.670 110.245 ;
        RECT 92.625 109.095 93.695 109.265 ;
        RECT 93.940 108.885 94.245 109.345 ;
        RECT 94.415 109.065 94.670 109.595 ;
        RECT 95.765 108.885 96.055 109.610 ;
        RECT 96.225 109.560 96.395 110.360 ;
        RECT 96.680 110.335 97.345 110.505 ;
        RECT 96.680 110.190 96.850 110.335 ;
        RECT 96.565 109.860 96.850 110.190 ;
        RECT 96.680 109.605 96.850 109.860 ;
        RECT 97.085 109.785 97.415 110.155 ;
        RECT 97.610 109.775 97.960 110.425 ;
        RECT 98.130 109.605 98.360 110.595 ;
        RECT 96.225 109.055 96.485 109.560 ;
        RECT 96.680 109.435 97.345 109.605 ;
        RECT 96.665 108.885 96.995 109.265 ;
        RECT 97.175 109.055 97.345 109.435 ;
        RECT 97.610 109.435 98.360 109.605 ;
        RECT 97.610 109.145 97.865 109.435 ;
        RECT 98.035 108.885 98.365 109.265 ;
        RECT 98.535 109.145 98.705 111.265 ;
        RECT 98.875 110.465 99.200 111.250 ;
        RECT 99.370 110.975 99.620 111.435 ;
        RECT 99.790 110.935 100.040 111.265 ;
        RECT 100.255 110.935 100.935 111.265 ;
        RECT 99.790 110.805 99.960 110.935 ;
        RECT 99.565 110.635 99.960 110.805 ;
        RECT 98.935 109.415 99.395 110.465 ;
        RECT 99.565 109.275 99.735 110.635 ;
        RECT 100.130 110.375 100.595 110.765 ;
        RECT 99.905 109.565 100.255 110.185 ;
        RECT 100.425 109.785 100.595 110.375 ;
        RECT 100.765 110.155 100.935 110.935 ;
        RECT 101.105 110.835 101.275 111.175 ;
        RECT 101.510 111.005 101.840 111.435 ;
        RECT 102.010 110.835 102.180 111.175 ;
        RECT 102.475 110.975 102.845 111.435 ;
        RECT 101.105 110.665 102.180 110.835 ;
        RECT 103.015 110.805 103.185 111.265 ;
        RECT 103.420 110.925 104.290 111.265 ;
        RECT 104.460 110.975 104.710 111.435 ;
        RECT 102.625 110.635 103.185 110.805 ;
        RECT 102.625 110.495 102.795 110.635 ;
        RECT 101.295 110.325 102.795 110.495 ;
        RECT 103.490 110.465 103.950 110.755 ;
        RECT 100.765 109.985 102.455 110.155 ;
        RECT 100.425 109.565 100.780 109.785 ;
        RECT 100.950 109.275 101.120 109.985 ;
        RECT 101.325 109.565 102.115 109.815 ;
        RECT 102.285 109.805 102.455 109.985 ;
        RECT 102.625 109.635 102.795 110.325 ;
        RECT 99.065 108.885 99.395 109.245 ;
        RECT 99.565 109.105 100.060 109.275 ;
        RECT 100.265 109.105 101.120 109.275 ;
        RECT 101.995 108.885 102.325 109.345 ;
        RECT 102.535 109.245 102.795 109.635 ;
        RECT 102.985 110.455 103.950 110.465 ;
        RECT 104.120 110.545 104.290 110.925 ;
        RECT 104.880 110.885 105.050 111.175 ;
        RECT 105.230 111.055 105.560 111.435 ;
        RECT 104.880 110.715 105.680 110.885 ;
        RECT 102.985 110.295 103.660 110.455 ;
        RECT 104.120 110.375 105.340 110.545 ;
        RECT 102.985 109.505 103.195 110.295 ;
        RECT 104.120 110.285 104.290 110.375 ;
        RECT 103.365 109.505 103.715 110.125 ;
        RECT 103.885 110.115 104.290 110.285 ;
        RECT 103.885 109.335 104.055 110.115 ;
        RECT 104.225 109.665 104.445 109.945 ;
        RECT 104.625 109.835 105.165 110.205 ;
        RECT 105.510 110.125 105.680 110.715 ;
        RECT 105.900 110.295 106.205 111.435 ;
        RECT 106.375 110.245 106.630 111.125 ;
        RECT 106.805 111.000 112.150 111.435 ;
        RECT 105.510 110.095 106.250 110.125 ;
        RECT 104.225 109.495 104.755 109.665 ;
        RECT 102.535 109.075 102.885 109.245 ;
        RECT 103.105 109.055 104.055 109.335 ;
        RECT 104.225 108.885 104.415 109.325 ;
        RECT 104.585 109.265 104.755 109.495 ;
        RECT 104.925 109.435 105.165 109.835 ;
        RECT 105.335 109.795 106.250 110.095 ;
        RECT 105.335 109.620 105.660 109.795 ;
        RECT 105.335 109.265 105.655 109.620 ;
        RECT 106.420 109.595 106.630 110.245 ;
        RECT 104.585 109.095 105.655 109.265 ;
        RECT 105.900 108.885 106.205 109.345 ;
        RECT 106.375 109.065 106.630 109.595 ;
        RECT 108.390 109.430 108.730 110.260 ;
        RECT 110.210 109.750 110.560 111.000 ;
        RECT 112.325 110.345 113.535 111.435 ;
        RECT 112.325 109.805 112.845 110.345 ;
        RECT 113.015 109.635 113.535 110.175 ;
        RECT 106.805 108.885 112.150 109.430 ;
        RECT 112.325 108.885 113.535 109.635 ;
        RECT 5.520 108.715 113.620 108.885 ;
        RECT 5.605 107.965 6.815 108.715 ;
        RECT 6.990 108.165 7.245 108.455 ;
        RECT 7.415 108.335 7.745 108.715 ;
        RECT 6.990 107.995 7.740 108.165 ;
        RECT 5.605 107.425 6.125 107.965 ;
        RECT 6.295 107.255 6.815 107.795 ;
        RECT 5.605 106.165 6.815 107.255 ;
        RECT 6.990 107.175 7.340 107.825 ;
        RECT 7.510 107.005 7.740 107.995 ;
        RECT 6.990 106.835 7.740 107.005 ;
        RECT 6.990 106.335 7.245 106.835 ;
        RECT 7.415 106.165 7.745 106.665 ;
        RECT 7.915 106.335 8.085 108.455 ;
        RECT 8.445 108.355 8.775 108.715 ;
        RECT 8.945 108.325 9.440 108.495 ;
        RECT 9.645 108.325 10.500 108.495 ;
        RECT 8.315 107.135 8.775 108.185 ;
        RECT 8.255 106.350 8.580 107.135 ;
        RECT 8.945 106.965 9.115 108.325 ;
        RECT 9.285 107.415 9.635 108.035 ;
        RECT 9.805 107.815 10.160 108.035 ;
        RECT 9.805 107.225 9.975 107.815 ;
        RECT 10.330 107.615 10.500 108.325 ;
        RECT 11.375 108.255 11.705 108.715 ;
        RECT 11.915 108.355 12.265 108.525 ;
        RECT 10.705 107.785 11.495 108.035 ;
        RECT 11.915 107.965 12.175 108.355 ;
        RECT 12.485 108.265 13.435 108.545 ;
        RECT 13.605 108.275 13.795 108.715 ;
        RECT 13.965 108.335 15.035 108.505 ;
        RECT 11.665 107.615 11.835 107.795 ;
        RECT 8.945 106.795 9.340 106.965 ;
        RECT 9.510 106.835 9.975 107.225 ;
        RECT 10.145 107.445 11.835 107.615 ;
        RECT 9.170 106.665 9.340 106.795 ;
        RECT 10.145 106.665 10.315 107.445 ;
        RECT 12.005 107.275 12.175 107.965 ;
        RECT 10.675 107.105 12.175 107.275 ;
        RECT 12.365 107.305 12.575 108.095 ;
        RECT 12.745 107.475 13.095 108.095 ;
        RECT 13.265 107.485 13.435 108.265 ;
        RECT 13.965 108.105 14.135 108.335 ;
        RECT 13.605 107.935 14.135 108.105 ;
        RECT 13.605 107.655 13.825 107.935 ;
        RECT 14.305 107.765 14.545 108.165 ;
        RECT 13.265 107.315 13.670 107.485 ;
        RECT 14.005 107.395 14.545 107.765 ;
        RECT 14.715 107.980 15.035 108.335 ;
        RECT 15.280 108.255 15.585 108.715 ;
        RECT 15.755 108.005 16.010 108.535 ;
        RECT 14.715 107.805 15.040 107.980 ;
        RECT 14.715 107.505 15.630 107.805 ;
        RECT 14.890 107.475 15.630 107.505 ;
        RECT 12.365 107.145 13.040 107.305 ;
        RECT 13.500 107.225 13.670 107.315 ;
        RECT 12.365 107.135 13.330 107.145 ;
        RECT 12.005 106.965 12.175 107.105 ;
        RECT 8.750 106.165 9.000 106.625 ;
        RECT 9.170 106.335 9.420 106.665 ;
        RECT 9.635 106.335 10.315 106.665 ;
        RECT 10.485 106.765 11.560 106.935 ;
        RECT 12.005 106.795 12.565 106.965 ;
        RECT 12.870 106.845 13.330 107.135 ;
        RECT 13.500 107.055 14.720 107.225 ;
        RECT 10.485 106.425 10.655 106.765 ;
        RECT 10.890 106.165 11.220 106.595 ;
        RECT 11.390 106.425 11.560 106.765 ;
        RECT 11.855 106.165 12.225 106.625 ;
        RECT 12.395 106.335 12.565 106.795 ;
        RECT 13.500 106.675 13.670 107.055 ;
        RECT 14.890 106.885 15.060 107.475 ;
        RECT 15.800 107.355 16.010 108.005 ;
        RECT 16.245 107.895 16.455 108.715 ;
        RECT 16.625 107.915 16.955 108.545 ;
        RECT 12.800 106.335 13.670 106.675 ;
        RECT 14.260 106.715 15.060 106.885 ;
        RECT 13.840 106.165 14.090 106.625 ;
        RECT 14.260 106.425 14.430 106.715 ;
        RECT 14.610 106.165 14.940 106.545 ;
        RECT 15.280 106.165 15.585 107.305 ;
        RECT 15.755 106.475 16.010 107.355 ;
        RECT 16.625 107.315 16.875 107.915 ;
        RECT 17.125 107.895 17.355 108.715 ;
        RECT 17.625 107.895 17.835 108.715 ;
        RECT 18.005 107.915 18.335 108.545 ;
        RECT 17.045 107.475 17.375 107.725 ;
        RECT 18.005 107.315 18.255 107.915 ;
        RECT 18.505 107.895 18.735 108.715 ;
        RECT 19.865 108.040 20.125 108.545 ;
        RECT 20.305 108.335 20.635 108.715 ;
        RECT 20.815 108.165 20.985 108.545 ;
        RECT 18.425 107.475 18.755 107.725 ;
        RECT 16.245 106.165 16.455 107.305 ;
        RECT 16.625 106.335 16.955 107.315 ;
        RECT 17.125 106.165 17.355 107.305 ;
        RECT 17.625 106.165 17.835 107.305 ;
        RECT 18.005 106.335 18.335 107.315 ;
        RECT 18.505 106.165 18.735 107.305 ;
        RECT 19.865 107.240 20.035 108.040 ;
        RECT 20.320 107.995 20.985 108.165 ;
        RECT 20.320 107.740 20.490 107.995 ;
        RECT 21.245 107.965 22.455 108.715 ;
        RECT 22.625 108.040 22.885 108.545 ;
        RECT 23.065 108.335 23.395 108.715 ;
        RECT 23.575 108.165 23.745 108.545 ;
        RECT 20.205 107.410 20.490 107.740 ;
        RECT 20.725 107.445 21.055 107.815 ;
        RECT 21.245 107.425 21.765 107.965 ;
        RECT 20.320 107.265 20.490 107.410 ;
        RECT 19.865 106.335 20.135 107.240 ;
        RECT 20.320 107.095 20.985 107.265 ;
        RECT 21.935 107.255 22.455 107.795 ;
        RECT 20.305 106.165 20.635 106.925 ;
        RECT 20.815 106.335 20.985 107.095 ;
        RECT 21.245 106.165 22.455 107.255 ;
        RECT 22.625 107.240 22.795 108.040 ;
        RECT 23.080 107.995 23.745 108.165 ;
        RECT 24.465 108.040 24.725 108.545 ;
        RECT 24.905 108.335 25.235 108.715 ;
        RECT 25.415 108.165 25.585 108.545 ;
        RECT 23.080 107.740 23.250 107.995 ;
        RECT 22.965 107.410 23.250 107.740 ;
        RECT 23.485 107.445 23.815 107.815 ;
        RECT 23.080 107.265 23.250 107.410 ;
        RECT 22.625 106.335 22.895 107.240 ;
        RECT 23.080 107.095 23.745 107.265 ;
        RECT 23.065 106.165 23.395 106.925 ;
        RECT 23.575 106.335 23.745 107.095 ;
        RECT 24.465 107.240 24.635 108.040 ;
        RECT 24.920 107.995 25.585 108.165 ;
        RECT 24.920 107.740 25.090 107.995 ;
        RECT 25.905 107.895 26.115 108.715 ;
        RECT 26.285 107.915 26.615 108.545 ;
        RECT 24.805 107.410 25.090 107.740 ;
        RECT 25.325 107.445 25.655 107.815 ;
        RECT 24.920 107.265 25.090 107.410 ;
        RECT 26.285 107.315 26.535 107.915 ;
        RECT 26.785 107.895 27.015 108.715 ;
        RECT 27.225 107.945 30.735 108.715 ;
        RECT 31.365 107.990 31.655 108.715 ;
        RECT 31.825 108.170 37.170 108.715 ;
        RECT 26.705 107.475 27.035 107.725 ;
        RECT 27.225 107.425 28.875 107.945 ;
        RECT 24.465 106.335 24.735 107.240 ;
        RECT 24.920 107.095 25.585 107.265 ;
        RECT 24.905 106.165 25.235 106.925 ;
        RECT 25.415 106.335 25.585 107.095 ;
        RECT 25.905 106.165 26.115 107.305 ;
        RECT 26.285 106.335 26.615 107.315 ;
        RECT 26.785 106.165 27.015 107.305 ;
        RECT 29.045 107.255 30.735 107.775 ;
        RECT 33.410 107.340 33.750 108.170 ;
        RECT 37.345 107.945 39.015 108.715 ;
        RECT 39.185 108.040 39.445 108.545 ;
        RECT 39.625 108.335 39.955 108.715 ;
        RECT 40.135 108.165 40.305 108.545 ;
        RECT 27.225 106.165 30.735 107.255 ;
        RECT 31.365 106.165 31.655 107.330 ;
        RECT 35.230 106.600 35.580 107.850 ;
        RECT 37.345 107.425 38.095 107.945 ;
        RECT 38.265 107.255 39.015 107.775 ;
        RECT 31.825 106.165 37.170 106.600 ;
        RECT 37.345 106.165 39.015 107.255 ;
        RECT 39.185 107.240 39.355 108.040 ;
        RECT 39.640 107.995 40.305 108.165 ;
        RECT 39.640 107.740 39.810 107.995 ;
        RECT 40.625 107.895 40.835 108.715 ;
        RECT 41.005 107.915 41.335 108.545 ;
        RECT 39.525 107.410 39.810 107.740 ;
        RECT 40.045 107.445 40.375 107.815 ;
        RECT 39.640 107.265 39.810 107.410 ;
        RECT 41.005 107.315 41.255 107.915 ;
        RECT 41.505 107.895 41.735 108.715 ;
        RECT 42.405 108.040 42.665 108.545 ;
        RECT 42.845 108.335 43.175 108.715 ;
        RECT 43.355 108.165 43.525 108.545 ;
        RECT 41.425 107.475 41.755 107.725 ;
        RECT 39.185 106.335 39.455 107.240 ;
        RECT 39.640 107.095 40.305 107.265 ;
        RECT 39.625 106.165 39.955 106.925 ;
        RECT 40.135 106.335 40.305 107.095 ;
        RECT 40.625 106.165 40.835 107.305 ;
        RECT 41.005 106.335 41.335 107.315 ;
        RECT 41.505 106.165 41.735 107.305 ;
        RECT 42.405 107.240 42.575 108.040 ;
        RECT 42.860 107.995 43.525 108.165 ;
        RECT 42.860 107.740 43.030 107.995 ;
        RECT 43.845 107.895 44.055 108.715 ;
        RECT 44.225 107.915 44.555 108.545 ;
        RECT 42.745 107.410 43.030 107.740 ;
        RECT 43.265 107.445 43.595 107.815 ;
        RECT 42.860 107.265 43.030 107.410 ;
        RECT 44.225 107.315 44.475 107.915 ;
        RECT 44.725 107.895 44.955 108.715 ;
        RECT 45.165 107.945 48.675 108.715 ;
        RECT 44.645 107.475 44.975 107.725 ;
        RECT 45.165 107.425 46.815 107.945 ;
        RECT 49.915 107.915 50.245 108.715 ;
        RECT 50.415 108.065 50.585 108.545 ;
        RECT 50.755 108.235 51.085 108.715 ;
        RECT 51.255 108.065 51.425 108.545 ;
        RECT 51.675 108.235 51.915 108.715 ;
        RECT 52.095 108.065 52.265 108.545 ;
        RECT 50.415 107.895 51.425 108.065 ;
        RECT 51.630 107.895 52.265 108.065 ;
        RECT 52.525 108.040 52.785 108.545 ;
        RECT 52.965 108.335 53.295 108.715 ;
        RECT 53.475 108.165 53.645 108.545 ;
        RECT 50.415 107.865 50.915 107.895 ;
        RECT 42.405 106.335 42.675 107.240 ;
        RECT 42.860 107.095 43.525 107.265 ;
        RECT 42.845 106.165 43.175 106.925 ;
        RECT 43.355 106.335 43.525 107.095 ;
        RECT 43.845 106.165 44.055 107.305 ;
        RECT 44.225 106.335 44.555 107.315 ;
        RECT 44.725 106.165 44.955 107.305 ;
        RECT 46.985 107.255 48.675 107.775 ;
        RECT 50.415 107.355 50.910 107.865 ;
        RECT 51.630 107.725 51.800 107.895 ;
        RECT 51.300 107.555 51.800 107.725 ;
        RECT 45.165 106.165 48.675 107.255 ;
        RECT 49.915 106.165 50.245 107.315 ;
        RECT 50.415 107.185 51.425 107.355 ;
        RECT 50.415 106.335 50.585 107.185 ;
        RECT 50.755 106.165 51.085 106.965 ;
        RECT 51.255 106.335 51.425 107.185 ;
        RECT 51.630 107.315 51.800 107.555 ;
        RECT 51.970 107.485 52.350 107.725 ;
        RECT 51.630 107.145 52.345 107.315 ;
        RECT 51.605 106.165 51.845 106.965 ;
        RECT 52.015 106.335 52.345 107.145 ;
        RECT 52.525 107.240 52.695 108.040 ;
        RECT 52.980 107.995 53.645 108.165 ;
        RECT 52.980 107.740 53.150 107.995 ;
        RECT 53.905 107.945 56.495 108.715 ;
        RECT 57.125 107.990 57.415 108.715 ;
        RECT 57.585 107.945 61.095 108.715 ;
        RECT 61.265 107.965 62.475 108.715 ;
        RECT 62.645 108.040 62.905 108.545 ;
        RECT 63.085 108.335 63.415 108.715 ;
        RECT 63.595 108.165 63.765 108.545 ;
        RECT 52.865 107.410 53.150 107.740 ;
        RECT 53.385 107.445 53.715 107.815 ;
        RECT 53.905 107.425 55.115 107.945 ;
        RECT 52.980 107.265 53.150 107.410 ;
        RECT 52.525 106.335 52.795 107.240 ;
        RECT 52.980 107.095 53.645 107.265 ;
        RECT 55.285 107.255 56.495 107.775 ;
        RECT 57.585 107.425 59.235 107.945 ;
        RECT 52.965 106.165 53.295 106.925 ;
        RECT 53.475 106.335 53.645 107.095 ;
        RECT 53.905 106.165 56.495 107.255 ;
        RECT 57.125 106.165 57.415 107.330 ;
        RECT 59.405 107.255 61.095 107.775 ;
        RECT 61.265 107.425 61.785 107.965 ;
        RECT 61.955 107.255 62.475 107.795 ;
        RECT 57.585 106.165 61.095 107.255 ;
        RECT 61.265 106.165 62.475 107.255 ;
        RECT 62.645 107.240 62.815 108.040 ;
        RECT 63.100 107.995 63.765 108.165 ;
        RECT 63.100 107.740 63.270 107.995 ;
        RECT 64.025 107.945 65.695 108.715 ;
        RECT 62.985 107.410 63.270 107.740 ;
        RECT 63.505 107.445 63.835 107.815 ;
        RECT 64.025 107.425 64.775 107.945 ;
        RECT 65.925 107.895 66.135 108.715 ;
        RECT 66.305 107.915 66.635 108.545 ;
        RECT 63.100 107.265 63.270 107.410 ;
        RECT 62.645 106.335 62.915 107.240 ;
        RECT 63.100 107.095 63.765 107.265 ;
        RECT 64.945 107.255 65.695 107.775 ;
        RECT 66.305 107.315 66.555 107.915 ;
        RECT 66.805 107.895 67.035 108.715 ;
        RECT 67.245 107.965 68.455 108.715 ;
        RECT 66.725 107.475 67.055 107.725 ;
        RECT 67.245 107.425 67.765 107.965 ;
        RECT 68.775 107.915 69.105 108.715 ;
        RECT 69.275 108.065 69.445 108.545 ;
        RECT 69.615 108.235 69.945 108.715 ;
        RECT 70.115 108.065 70.285 108.545 ;
        RECT 70.535 108.235 70.775 108.715 ;
        RECT 70.955 108.065 71.125 108.545 ;
        RECT 69.275 107.895 70.285 108.065 ;
        RECT 70.490 107.895 71.125 108.065 ;
        RECT 71.385 107.945 73.055 108.715 ;
        RECT 63.085 106.165 63.415 106.925 ;
        RECT 63.595 106.335 63.765 107.095 ;
        RECT 64.025 106.165 65.695 107.255 ;
        RECT 65.925 106.165 66.135 107.305 ;
        RECT 66.305 106.335 66.635 107.315 ;
        RECT 66.805 106.165 67.035 107.305 ;
        RECT 67.935 107.255 68.455 107.795 ;
        RECT 69.275 107.695 69.770 107.895 ;
        RECT 70.490 107.725 70.660 107.895 ;
        RECT 69.275 107.525 69.775 107.695 ;
        RECT 70.160 107.555 70.660 107.725 ;
        RECT 69.275 107.355 69.770 107.525 ;
        RECT 67.245 106.165 68.455 107.255 ;
        RECT 68.775 106.165 69.105 107.315 ;
        RECT 69.275 107.185 70.285 107.355 ;
        RECT 69.275 106.335 69.445 107.185 ;
        RECT 69.615 106.165 69.945 106.965 ;
        RECT 70.115 106.335 70.285 107.185 ;
        RECT 70.490 107.315 70.660 107.555 ;
        RECT 70.830 107.485 71.210 107.725 ;
        RECT 71.385 107.425 72.135 107.945 ;
        RECT 73.265 107.895 73.495 108.715 ;
        RECT 73.665 107.915 73.995 108.545 ;
        RECT 70.490 107.145 71.205 107.315 ;
        RECT 72.305 107.255 73.055 107.775 ;
        RECT 73.245 107.475 73.575 107.725 ;
        RECT 73.745 107.315 73.995 107.915 ;
        RECT 74.165 107.895 74.375 108.715 ;
        RECT 74.605 107.945 78.115 108.715 ;
        RECT 78.285 108.040 78.545 108.545 ;
        RECT 78.725 108.335 79.055 108.715 ;
        RECT 79.235 108.165 79.405 108.545 ;
        RECT 74.605 107.425 76.255 107.945 ;
        RECT 70.465 106.165 70.705 106.965 ;
        RECT 70.875 106.335 71.205 107.145 ;
        RECT 71.385 106.165 73.055 107.255 ;
        RECT 73.265 106.165 73.495 107.305 ;
        RECT 73.665 106.335 73.995 107.315 ;
        RECT 74.165 106.165 74.375 107.305 ;
        RECT 76.425 107.255 78.115 107.775 ;
        RECT 74.605 106.165 78.115 107.255 ;
        RECT 78.285 107.240 78.455 108.040 ;
        RECT 78.740 107.995 79.405 108.165 ;
        RECT 78.740 107.740 78.910 107.995 ;
        RECT 79.665 107.945 82.255 108.715 ;
        RECT 82.885 107.990 83.175 108.715 ;
        RECT 83.345 107.945 86.855 108.715 ;
        RECT 87.025 108.040 87.285 108.545 ;
        RECT 87.465 108.335 87.795 108.715 ;
        RECT 87.975 108.165 88.145 108.545 ;
        RECT 88.405 108.170 93.750 108.715 ;
        RECT 78.625 107.410 78.910 107.740 ;
        RECT 79.145 107.445 79.475 107.815 ;
        RECT 79.665 107.425 80.875 107.945 ;
        RECT 78.740 107.265 78.910 107.410 ;
        RECT 78.285 106.335 78.555 107.240 ;
        RECT 78.740 107.095 79.405 107.265 ;
        RECT 81.045 107.255 82.255 107.775 ;
        RECT 83.345 107.425 84.995 107.945 ;
        RECT 78.725 106.165 79.055 106.925 ;
        RECT 79.235 106.335 79.405 107.095 ;
        RECT 79.665 106.165 82.255 107.255 ;
        RECT 82.885 106.165 83.175 107.330 ;
        RECT 85.165 107.255 86.855 107.775 ;
        RECT 83.345 106.165 86.855 107.255 ;
        RECT 87.025 107.240 87.195 108.040 ;
        RECT 87.480 107.995 88.145 108.165 ;
        RECT 87.480 107.740 87.650 107.995 ;
        RECT 87.365 107.410 87.650 107.740 ;
        RECT 87.885 107.445 88.215 107.815 ;
        RECT 87.480 107.265 87.650 107.410 ;
        RECT 89.990 107.340 90.330 108.170 ;
        RECT 93.925 107.945 95.595 108.715 ;
        RECT 96.315 108.165 96.485 108.545 ;
        RECT 96.665 108.335 96.995 108.715 ;
        RECT 96.315 107.995 96.980 108.165 ;
        RECT 97.175 108.040 97.435 108.545 ;
        RECT 87.025 106.335 87.295 107.240 ;
        RECT 87.480 107.095 88.145 107.265 ;
        RECT 87.465 106.165 87.795 106.925 ;
        RECT 87.975 106.335 88.145 107.095 ;
        RECT 91.810 106.600 92.160 107.850 ;
        RECT 93.925 107.425 94.675 107.945 ;
        RECT 94.845 107.255 95.595 107.775 ;
        RECT 96.245 107.445 96.575 107.815 ;
        RECT 96.810 107.740 96.980 107.995 ;
        RECT 96.810 107.410 97.095 107.740 ;
        RECT 96.810 107.265 96.980 107.410 ;
        RECT 88.405 106.165 93.750 106.600 ;
        RECT 93.925 106.165 95.595 107.255 ;
        RECT 96.315 107.095 96.980 107.265 ;
        RECT 97.265 107.240 97.435 108.040 ;
        RECT 98.530 108.165 98.785 108.455 ;
        RECT 98.955 108.335 99.285 108.715 ;
        RECT 98.530 107.995 99.280 108.165 ;
        RECT 96.315 106.335 96.485 107.095 ;
        RECT 96.665 106.165 96.995 106.925 ;
        RECT 97.165 106.335 97.435 107.240 ;
        RECT 98.530 107.175 98.880 107.825 ;
        RECT 99.050 107.005 99.280 107.995 ;
        RECT 98.530 106.835 99.280 107.005 ;
        RECT 98.530 106.335 98.785 106.835 ;
        RECT 98.955 106.165 99.285 106.665 ;
        RECT 99.455 106.335 99.625 108.455 ;
        RECT 99.985 108.355 100.315 108.715 ;
        RECT 100.485 108.325 100.980 108.495 ;
        RECT 101.185 108.325 102.040 108.495 ;
        RECT 99.855 107.135 100.315 108.185 ;
        RECT 99.795 106.350 100.120 107.135 ;
        RECT 100.485 106.965 100.655 108.325 ;
        RECT 100.825 107.415 101.175 108.035 ;
        RECT 101.345 107.815 101.700 108.035 ;
        RECT 101.345 107.225 101.515 107.815 ;
        RECT 101.870 107.615 102.040 108.325 ;
        RECT 102.915 108.255 103.245 108.715 ;
        RECT 103.455 108.355 103.805 108.525 ;
        RECT 102.245 107.785 103.035 108.035 ;
        RECT 103.455 107.965 103.715 108.355 ;
        RECT 104.025 108.265 104.975 108.545 ;
        RECT 105.145 108.275 105.335 108.715 ;
        RECT 105.505 108.335 106.575 108.505 ;
        RECT 103.205 107.615 103.375 107.795 ;
        RECT 100.485 106.795 100.880 106.965 ;
        RECT 101.050 106.835 101.515 107.225 ;
        RECT 101.685 107.445 103.375 107.615 ;
        RECT 100.710 106.665 100.880 106.795 ;
        RECT 101.685 106.665 101.855 107.445 ;
        RECT 103.545 107.275 103.715 107.965 ;
        RECT 102.215 107.105 103.715 107.275 ;
        RECT 103.905 107.305 104.115 108.095 ;
        RECT 104.285 107.475 104.635 108.095 ;
        RECT 104.805 107.485 104.975 108.265 ;
        RECT 105.505 108.105 105.675 108.335 ;
        RECT 105.145 107.935 105.675 108.105 ;
        RECT 105.145 107.655 105.365 107.935 ;
        RECT 105.845 107.765 106.085 108.165 ;
        RECT 104.805 107.315 105.210 107.485 ;
        RECT 105.545 107.395 106.085 107.765 ;
        RECT 106.255 107.980 106.575 108.335 ;
        RECT 106.820 108.255 107.125 108.715 ;
        RECT 107.295 108.005 107.550 108.535 ;
        RECT 106.255 107.805 106.580 107.980 ;
        RECT 106.255 107.505 107.170 107.805 ;
        RECT 106.430 107.475 107.170 107.505 ;
        RECT 103.905 107.145 104.580 107.305 ;
        RECT 105.040 107.225 105.210 107.315 ;
        RECT 103.905 107.135 104.870 107.145 ;
        RECT 103.545 106.965 103.715 107.105 ;
        RECT 100.290 106.165 100.540 106.625 ;
        RECT 100.710 106.335 100.960 106.665 ;
        RECT 101.175 106.335 101.855 106.665 ;
        RECT 102.025 106.765 103.100 106.935 ;
        RECT 103.545 106.795 104.105 106.965 ;
        RECT 104.410 106.845 104.870 107.135 ;
        RECT 105.040 107.055 106.260 107.225 ;
        RECT 102.025 106.425 102.195 106.765 ;
        RECT 102.430 106.165 102.760 106.595 ;
        RECT 102.930 106.425 103.100 106.765 ;
        RECT 103.395 106.165 103.765 106.625 ;
        RECT 103.935 106.335 104.105 106.795 ;
        RECT 105.040 106.675 105.210 107.055 ;
        RECT 106.430 106.885 106.600 107.475 ;
        RECT 107.340 107.355 107.550 108.005 ;
        RECT 108.645 107.990 108.935 108.715 ;
        RECT 109.105 107.945 111.695 108.715 ;
        RECT 112.325 107.965 113.535 108.715 ;
        RECT 109.105 107.425 110.315 107.945 ;
        RECT 104.340 106.335 105.210 106.675 ;
        RECT 105.800 106.715 106.600 106.885 ;
        RECT 105.380 106.165 105.630 106.625 ;
        RECT 105.800 106.425 105.970 106.715 ;
        RECT 106.150 106.165 106.480 106.545 ;
        RECT 106.820 106.165 107.125 107.305 ;
        RECT 107.295 106.475 107.550 107.355 ;
        RECT 108.645 106.165 108.935 107.330 ;
        RECT 110.485 107.255 111.695 107.775 ;
        RECT 109.105 106.165 111.695 107.255 ;
        RECT 112.325 107.255 112.845 107.795 ;
        RECT 113.015 107.425 113.535 107.965 ;
        RECT 112.325 106.165 113.535 107.255 ;
        RECT 5.520 105.995 113.620 106.165 ;
        RECT 5.605 104.905 6.815 105.995 ;
        RECT 6.985 104.905 9.575 105.995 ;
        RECT 5.605 104.195 6.125 104.735 ;
        RECT 6.295 104.365 6.815 104.905 ;
        RECT 6.985 104.215 8.195 104.735 ;
        RECT 8.365 104.385 9.575 104.905 ;
        RECT 9.745 104.920 10.015 105.825 ;
        RECT 10.185 105.235 10.515 105.995 ;
        RECT 10.695 105.065 10.865 105.825 ;
        RECT 5.605 103.445 6.815 104.195 ;
        RECT 6.985 103.445 9.575 104.215 ;
        RECT 9.745 104.120 9.915 104.920 ;
        RECT 10.200 104.895 10.865 105.065 ;
        RECT 12.045 104.920 12.315 105.825 ;
        RECT 12.485 105.235 12.815 105.995 ;
        RECT 12.995 105.065 13.165 105.825 ;
        RECT 10.200 104.750 10.370 104.895 ;
        RECT 10.085 104.420 10.370 104.750 ;
        RECT 10.200 104.165 10.370 104.420 ;
        RECT 10.605 104.345 10.935 104.715 ;
        RECT 9.745 103.615 10.005 104.120 ;
        RECT 10.200 103.995 10.865 104.165 ;
        RECT 10.185 103.445 10.515 103.825 ;
        RECT 10.695 103.615 10.865 103.995 ;
        RECT 12.045 104.120 12.215 104.920 ;
        RECT 12.500 104.895 13.165 105.065 ;
        RECT 12.500 104.750 12.670 104.895 ;
        RECT 14.405 104.855 14.615 105.995 ;
        RECT 12.385 104.420 12.670 104.750 ;
        RECT 14.785 104.845 15.115 105.825 ;
        RECT 15.285 104.855 15.515 105.995 ;
        RECT 15.725 104.905 18.315 105.995 ;
        RECT 12.500 104.165 12.670 104.420 ;
        RECT 12.905 104.345 13.235 104.715 ;
        RECT 12.045 103.615 12.305 104.120 ;
        RECT 12.500 103.995 13.165 104.165 ;
        RECT 12.485 103.445 12.815 103.825 ;
        RECT 12.995 103.615 13.165 103.995 ;
        RECT 14.405 103.445 14.615 104.265 ;
        RECT 14.785 104.245 15.035 104.845 ;
        RECT 15.205 104.435 15.535 104.685 ;
        RECT 14.785 103.615 15.115 104.245 ;
        RECT 15.285 103.445 15.515 104.265 ;
        RECT 15.725 104.215 16.935 104.735 ;
        RECT 17.105 104.385 18.315 104.905 ;
        RECT 18.485 104.830 18.775 105.995 ;
        RECT 18.945 105.560 24.290 105.995 ;
        RECT 24.465 105.560 29.810 105.995 ;
        RECT 29.985 105.560 35.330 105.995 ;
        RECT 15.725 103.445 18.315 104.215 ;
        RECT 18.485 103.445 18.775 104.170 ;
        RECT 20.530 103.990 20.870 104.820 ;
        RECT 22.350 104.310 22.700 105.560 ;
        RECT 26.050 103.990 26.390 104.820 ;
        RECT 27.870 104.310 28.220 105.560 ;
        RECT 31.570 103.990 31.910 104.820 ;
        RECT 33.390 104.310 33.740 105.560 ;
        RECT 35.565 104.855 35.775 105.995 ;
        RECT 35.945 104.845 36.275 105.825 ;
        RECT 36.445 104.855 36.675 105.995 ;
        RECT 36.885 105.560 42.230 105.995 ;
        RECT 18.945 103.445 24.290 103.990 ;
        RECT 24.465 103.445 29.810 103.990 ;
        RECT 29.985 103.445 35.330 103.990 ;
        RECT 35.565 103.445 35.775 104.265 ;
        RECT 35.945 104.245 36.195 104.845 ;
        RECT 36.365 104.435 36.695 104.685 ;
        RECT 35.945 103.615 36.275 104.245 ;
        RECT 36.445 103.445 36.675 104.265 ;
        RECT 38.470 103.990 38.810 104.820 ;
        RECT 40.290 104.310 40.640 105.560 ;
        RECT 42.405 104.905 44.075 105.995 ;
        RECT 42.405 104.215 43.155 104.735 ;
        RECT 43.325 104.385 44.075 104.905 ;
        RECT 44.245 104.830 44.535 105.995 ;
        RECT 44.705 104.905 45.915 105.995 ;
        RECT 36.885 103.445 42.230 103.990 ;
        RECT 42.405 103.445 44.075 104.215 ;
        RECT 44.705 104.195 45.225 104.735 ;
        RECT 45.395 104.365 45.915 104.905 ;
        RECT 46.090 104.855 46.425 105.825 ;
        RECT 46.595 104.855 46.765 105.995 ;
        RECT 46.935 105.655 48.965 105.825 ;
        RECT 44.245 103.445 44.535 104.170 ;
        RECT 44.705 103.445 45.915 104.195 ;
        RECT 46.090 104.185 46.260 104.855 ;
        RECT 46.935 104.685 47.105 105.655 ;
        RECT 46.430 104.355 46.685 104.685 ;
        RECT 46.910 104.355 47.105 104.685 ;
        RECT 47.275 105.315 48.400 105.485 ;
        RECT 46.515 104.185 46.685 104.355 ;
        RECT 47.275 104.185 47.445 105.315 ;
        RECT 46.090 103.615 46.345 104.185 ;
        RECT 46.515 104.015 47.445 104.185 ;
        RECT 47.615 104.975 48.625 105.145 ;
        RECT 47.615 104.175 47.785 104.975 ;
        RECT 47.990 104.295 48.265 104.775 ;
        RECT 47.985 104.125 48.265 104.295 ;
        RECT 47.270 103.980 47.445 104.015 ;
        RECT 46.515 103.445 46.845 103.845 ;
        RECT 47.270 103.615 47.800 103.980 ;
        RECT 47.990 103.615 48.265 104.125 ;
        RECT 48.435 103.615 48.625 104.975 ;
        RECT 48.795 104.990 48.965 105.655 ;
        RECT 49.135 105.235 49.305 105.995 ;
        RECT 49.540 105.235 50.055 105.645 ;
        RECT 50.225 105.560 55.570 105.995 ;
        RECT 55.745 105.560 61.090 105.995 ;
        RECT 61.265 105.560 66.610 105.995 ;
        RECT 48.795 104.800 49.545 104.990 ;
        RECT 49.715 104.425 50.055 105.235 ;
        RECT 48.825 104.255 50.055 104.425 ;
        RECT 48.805 103.445 49.315 103.980 ;
        RECT 49.535 103.650 49.780 104.255 ;
        RECT 51.810 103.990 52.150 104.820 ;
        RECT 53.630 104.310 53.980 105.560 ;
        RECT 57.330 103.990 57.670 104.820 ;
        RECT 59.150 104.310 59.500 105.560 ;
        RECT 62.850 103.990 63.190 104.820 ;
        RECT 64.670 104.310 65.020 105.560 ;
        RECT 66.785 104.905 69.375 105.995 ;
        RECT 66.785 104.215 67.995 104.735 ;
        RECT 68.165 104.385 69.375 104.905 ;
        RECT 70.005 104.830 70.295 105.995 ;
        RECT 70.470 104.855 70.805 105.825 ;
        RECT 70.975 104.855 71.145 105.995 ;
        RECT 71.315 105.655 73.345 105.825 ;
        RECT 50.225 103.445 55.570 103.990 ;
        RECT 55.745 103.445 61.090 103.990 ;
        RECT 61.265 103.445 66.610 103.990 ;
        RECT 66.785 103.445 69.375 104.215 ;
        RECT 70.470 104.185 70.640 104.855 ;
        RECT 71.315 104.685 71.485 105.655 ;
        RECT 70.810 104.355 71.065 104.685 ;
        RECT 71.290 104.355 71.485 104.685 ;
        RECT 71.655 105.315 72.780 105.485 ;
        RECT 70.895 104.185 71.065 104.355 ;
        RECT 71.655 104.185 71.825 105.315 ;
        RECT 70.005 103.445 70.295 104.170 ;
        RECT 70.470 103.615 70.725 104.185 ;
        RECT 70.895 104.015 71.825 104.185 ;
        RECT 71.995 104.975 73.005 105.145 ;
        RECT 71.995 104.175 72.165 104.975 ;
        RECT 71.650 103.980 71.825 104.015 ;
        RECT 70.895 103.445 71.225 103.845 ;
        RECT 71.650 103.615 72.180 103.980 ;
        RECT 72.370 103.955 72.645 104.775 ;
        RECT 72.365 103.785 72.645 103.955 ;
        RECT 72.370 103.615 72.645 103.785 ;
        RECT 72.815 103.615 73.005 104.975 ;
        RECT 73.175 104.990 73.345 105.655 ;
        RECT 73.515 105.235 73.685 105.995 ;
        RECT 73.920 105.235 74.435 105.645 ;
        RECT 73.175 104.800 73.925 104.990 ;
        RECT 74.095 104.425 74.435 105.235 ;
        RECT 74.665 104.855 74.875 105.995 ;
        RECT 73.205 104.255 74.435 104.425 ;
        RECT 75.045 104.845 75.375 105.825 ;
        RECT 75.545 104.855 75.775 105.995 ;
        RECT 75.985 105.560 81.330 105.995 ;
        RECT 81.505 105.560 86.850 105.995 ;
        RECT 87.025 105.560 92.370 105.995 ;
        RECT 73.185 103.445 73.695 103.980 ;
        RECT 73.915 103.650 74.160 104.255 ;
        RECT 74.665 103.445 74.875 104.265 ;
        RECT 75.045 104.245 75.295 104.845 ;
        RECT 75.465 104.435 75.795 104.685 ;
        RECT 75.045 103.615 75.375 104.245 ;
        RECT 75.545 103.445 75.775 104.265 ;
        RECT 77.570 103.990 77.910 104.820 ;
        RECT 79.390 104.310 79.740 105.560 ;
        RECT 83.090 103.990 83.430 104.820 ;
        RECT 84.910 104.310 85.260 105.560 ;
        RECT 88.610 103.990 88.950 104.820 ;
        RECT 90.430 104.310 90.780 105.560 ;
        RECT 92.545 104.905 95.135 105.995 ;
        RECT 92.545 104.215 93.755 104.735 ;
        RECT 93.925 104.385 95.135 104.905 ;
        RECT 95.765 104.830 96.055 105.995 ;
        RECT 96.285 104.855 96.495 105.995 ;
        RECT 96.665 104.845 96.995 105.825 ;
        RECT 97.165 104.855 97.395 105.995 ;
        RECT 97.695 105.065 97.865 105.825 ;
        RECT 98.045 105.235 98.375 105.995 ;
        RECT 97.695 104.895 98.360 105.065 ;
        RECT 98.545 104.920 98.815 105.825 ;
        RECT 75.985 103.445 81.330 103.990 ;
        RECT 81.505 103.445 86.850 103.990 ;
        RECT 87.025 103.445 92.370 103.990 ;
        RECT 92.545 103.445 95.135 104.215 ;
        RECT 95.765 103.445 96.055 104.170 ;
        RECT 96.285 103.445 96.495 104.265 ;
        RECT 96.665 104.245 96.915 104.845 ;
        RECT 98.190 104.750 98.360 104.895 ;
        RECT 97.085 104.435 97.415 104.685 ;
        RECT 97.625 104.345 97.955 104.715 ;
        RECT 98.190 104.420 98.475 104.750 ;
        RECT 96.665 103.615 96.995 104.245 ;
        RECT 97.165 103.445 97.395 104.265 ;
        RECT 98.190 104.165 98.360 104.420 ;
        RECT 97.695 103.995 98.360 104.165 ;
        RECT 98.645 104.120 98.815 104.920 ;
        RECT 98.985 104.905 102.495 105.995 ;
        RECT 102.665 104.905 103.875 105.995 ;
        RECT 97.695 103.615 97.865 103.995 ;
        RECT 98.045 103.445 98.375 103.825 ;
        RECT 98.555 103.615 98.815 104.120 ;
        RECT 98.985 104.215 100.635 104.735 ;
        RECT 100.805 104.385 102.495 104.905 ;
        RECT 98.985 103.445 102.495 104.215 ;
        RECT 102.665 104.195 103.185 104.735 ;
        RECT 103.355 104.365 103.875 104.905 ;
        RECT 104.105 104.855 104.315 105.995 ;
        RECT 104.485 104.845 104.815 105.825 ;
        RECT 104.985 104.855 105.215 105.995 ;
        RECT 105.425 105.560 110.770 105.995 ;
        RECT 102.665 103.445 103.875 104.195 ;
        RECT 104.105 103.445 104.315 104.265 ;
        RECT 104.485 104.245 104.735 104.845 ;
        RECT 104.905 104.435 105.235 104.685 ;
        RECT 104.485 103.615 104.815 104.245 ;
        RECT 104.985 103.445 105.215 104.265 ;
        RECT 107.010 103.990 107.350 104.820 ;
        RECT 108.830 104.310 109.180 105.560 ;
        RECT 110.945 104.905 112.155 105.995 ;
        RECT 110.945 104.195 111.465 104.735 ;
        RECT 111.635 104.365 112.155 104.905 ;
        RECT 112.325 104.905 113.535 105.995 ;
        RECT 112.325 104.365 112.845 104.905 ;
        RECT 113.015 104.195 113.535 104.735 ;
        RECT 105.425 103.445 110.770 103.990 ;
        RECT 110.945 103.445 112.155 104.195 ;
        RECT 112.325 103.445 113.535 104.195 ;
        RECT 5.520 103.275 113.620 103.445 ;
        RECT 5.605 102.525 6.815 103.275 ;
        RECT 6.985 102.730 12.330 103.275 ;
        RECT 5.605 101.985 6.125 102.525 ;
        RECT 6.295 101.815 6.815 102.355 ;
        RECT 8.570 101.900 8.910 102.730 ;
        RECT 12.505 102.505 16.015 103.275 ;
        RECT 16.275 102.725 16.445 103.015 ;
        RECT 16.615 102.895 16.945 103.275 ;
        RECT 16.275 102.555 16.940 102.725 ;
        RECT 5.605 100.725 6.815 101.815 ;
        RECT 10.390 101.160 10.740 102.410 ;
        RECT 12.505 101.985 14.155 102.505 ;
        RECT 14.325 101.815 16.015 102.335 ;
        RECT 6.985 100.725 12.330 101.160 ;
        RECT 12.505 100.725 16.015 101.815 ;
        RECT 16.190 101.735 16.540 102.385 ;
        RECT 16.710 101.565 16.940 102.555 ;
        RECT 16.275 101.395 16.940 101.565 ;
        RECT 16.275 100.895 16.445 101.395 ;
        RECT 16.615 100.725 16.945 101.225 ;
        RECT 17.115 100.895 17.340 103.015 ;
        RECT 17.555 102.895 17.885 103.275 ;
        RECT 18.055 102.725 18.225 103.055 ;
        RECT 18.525 102.895 19.540 103.095 ;
        RECT 17.530 102.535 18.225 102.725 ;
        RECT 17.530 101.565 17.700 102.535 ;
        RECT 17.870 101.735 18.280 102.355 ;
        RECT 18.450 101.785 18.670 102.655 ;
        RECT 18.850 102.345 19.200 102.715 ;
        RECT 19.370 102.165 19.540 102.895 ;
        RECT 19.710 102.835 20.120 103.275 ;
        RECT 20.410 102.635 20.660 103.065 ;
        RECT 20.860 102.815 21.180 103.275 ;
        RECT 21.740 102.885 22.590 103.055 ;
        RECT 19.710 102.295 20.120 102.625 ;
        RECT 20.410 102.295 20.830 102.635 ;
        RECT 19.120 102.125 19.540 102.165 ;
        RECT 19.120 101.955 20.470 102.125 ;
        RECT 17.530 101.395 18.225 101.565 ;
        RECT 18.450 101.405 18.950 101.785 ;
        RECT 17.555 100.725 17.885 101.225 ;
        RECT 18.055 100.895 18.225 101.395 ;
        RECT 19.120 101.110 19.290 101.955 ;
        RECT 20.220 101.795 20.470 101.955 ;
        RECT 19.460 101.525 19.710 101.785 ;
        RECT 20.640 101.525 20.830 102.295 ;
        RECT 19.460 101.275 20.830 101.525 ;
        RECT 21.000 102.465 22.250 102.635 ;
        RECT 21.000 101.705 21.170 102.465 ;
        RECT 21.920 102.345 22.250 102.465 ;
        RECT 21.340 101.885 21.520 102.295 ;
        RECT 22.420 102.125 22.590 102.885 ;
        RECT 22.790 102.795 23.450 103.275 ;
        RECT 23.630 102.680 23.950 103.010 ;
        RECT 22.780 102.355 23.440 102.625 ;
        RECT 22.780 102.295 23.110 102.355 ;
        RECT 23.260 102.125 23.590 102.185 ;
        RECT 21.690 101.955 23.590 102.125 ;
        RECT 21.000 101.395 21.520 101.705 ;
        RECT 21.690 101.445 21.860 101.955 ;
        RECT 23.760 101.785 23.950 102.680 ;
        RECT 22.030 101.615 23.950 101.785 ;
        RECT 23.630 101.595 23.950 101.615 ;
        RECT 24.150 102.365 24.400 103.015 ;
        RECT 24.580 102.815 24.865 103.275 ;
        RECT 25.045 102.565 25.300 103.095 ;
        RECT 24.150 102.035 24.950 102.365 ;
        RECT 21.690 101.275 22.900 101.445 ;
        RECT 18.460 100.940 19.290 101.110 ;
        RECT 19.530 100.725 19.910 101.105 ;
        RECT 20.090 100.985 20.260 101.275 ;
        RECT 21.690 101.195 21.860 101.275 ;
        RECT 20.430 100.725 20.760 101.105 ;
        RECT 21.230 100.945 21.860 101.195 ;
        RECT 22.040 100.725 22.460 101.105 ;
        RECT 22.660 100.985 22.900 101.275 ;
        RECT 23.130 100.725 23.460 101.415 ;
        RECT 23.630 100.985 23.800 101.595 ;
        RECT 24.150 101.445 24.400 102.035 ;
        RECT 25.120 101.705 25.300 102.565 ;
        RECT 25.845 102.505 27.515 103.275 ;
        RECT 27.775 102.725 27.945 103.105 ;
        RECT 28.125 102.895 28.455 103.275 ;
        RECT 27.775 102.555 28.440 102.725 ;
        RECT 28.635 102.600 28.895 103.105 ;
        RECT 25.845 101.985 26.595 102.505 ;
        RECT 26.765 101.815 27.515 102.335 ;
        RECT 27.705 102.005 28.035 102.375 ;
        RECT 28.270 102.300 28.440 102.555 ;
        RECT 28.270 101.970 28.555 102.300 ;
        RECT 28.270 101.825 28.440 101.970 ;
        RECT 24.070 100.935 24.400 101.445 ;
        RECT 24.580 100.725 24.865 101.525 ;
        RECT 25.045 101.235 25.300 101.705 ;
        RECT 25.045 101.065 25.385 101.235 ;
        RECT 25.045 101.035 25.300 101.065 ;
        RECT 25.845 100.725 27.515 101.815 ;
        RECT 27.775 101.655 28.440 101.825 ;
        RECT 28.725 101.800 28.895 102.600 ;
        RECT 29.065 102.505 30.735 103.275 ;
        RECT 31.365 102.550 31.655 103.275 ;
        RECT 32.200 102.565 32.455 103.095 ;
        RECT 32.635 102.815 32.920 103.275 ;
        RECT 29.065 101.985 29.815 102.505 ;
        RECT 29.985 101.815 30.735 102.335 ;
        RECT 27.775 100.895 27.945 101.655 ;
        RECT 28.125 100.725 28.455 101.485 ;
        RECT 28.625 100.895 28.895 101.800 ;
        RECT 29.065 100.725 30.735 101.815 ;
        RECT 31.365 100.725 31.655 101.890 ;
        RECT 32.200 101.705 32.380 102.565 ;
        RECT 33.100 102.365 33.350 103.015 ;
        RECT 32.550 102.035 33.350 102.365 ;
        RECT 32.200 101.235 32.455 101.705 ;
        RECT 32.115 101.065 32.455 101.235 ;
        RECT 32.200 101.035 32.455 101.065 ;
        RECT 32.635 100.725 32.920 101.525 ;
        RECT 33.100 101.445 33.350 102.035 ;
        RECT 33.550 102.680 33.870 103.010 ;
        RECT 34.050 102.795 34.710 103.275 ;
        RECT 34.910 102.885 35.760 103.055 ;
        RECT 33.550 101.785 33.740 102.680 ;
        RECT 34.060 102.355 34.720 102.625 ;
        RECT 34.390 102.295 34.720 102.355 ;
        RECT 33.910 102.125 34.240 102.185 ;
        RECT 34.910 102.125 35.080 102.885 ;
        RECT 36.320 102.815 36.640 103.275 ;
        RECT 36.840 102.635 37.090 103.065 ;
        RECT 37.380 102.835 37.790 103.275 ;
        RECT 37.960 102.895 38.975 103.095 ;
        RECT 35.250 102.465 36.500 102.635 ;
        RECT 35.250 102.345 35.580 102.465 ;
        RECT 33.910 101.955 35.810 102.125 ;
        RECT 33.550 101.615 35.470 101.785 ;
        RECT 33.550 101.595 33.870 101.615 ;
        RECT 33.100 100.935 33.430 101.445 ;
        RECT 33.700 100.985 33.870 101.595 ;
        RECT 35.640 101.445 35.810 101.955 ;
        RECT 35.980 101.885 36.160 102.295 ;
        RECT 36.330 101.705 36.500 102.465 ;
        RECT 34.040 100.725 34.370 101.415 ;
        RECT 34.600 101.275 35.810 101.445 ;
        RECT 35.980 101.395 36.500 101.705 ;
        RECT 36.670 102.295 37.090 102.635 ;
        RECT 37.380 102.295 37.790 102.625 ;
        RECT 36.670 101.525 36.860 102.295 ;
        RECT 37.960 102.165 38.130 102.895 ;
        RECT 39.275 102.725 39.445 103.055 ;
        RECT 39.615 102.895 39.945 103.275 ;
        RECT 38.300 102.345 38.650 102.715 ;
        RECT 37.960 102.125 38.380 102.165 ;
        RECT 37.030 101.955 38.380 102.125 ;
        RECT 37.030 101.795 37.280 101.955 ;
        RECT 37.790 101.525 38.040 101.785 ;
        RECT 36.670 101.275 38.040 101.525 ;
        RECT 34.600 100.985 34.840 101.275 ;
        RECT 35.640 101.195 35.810 101.275 ;
        RECT 35.040 100.725 35.460 101.105 ;
        RECT 35.640 100.945 36.270 101.195 ;
        RECT 36.740 100.725 37.070 101.105 ;
        RECT 37.240 100.985 37.410 101.275 ;
        RECT 38.210 101.110 38.380 101.955 ;
        RECT 38.830 101.785 39.050 102.655 ;
        RECT 39.275 102.535 39.970 102.725 ;
        RECT 38.550 101.405 39.050 101.785 ;
        RECT 39.220 101.735 39.630 102.355 ;
        RECT 39.800 101.565 39.970 102.535 ;
        RECT 39.275 101.395 39.970 101.565 ;
        RECT 37.590 100.725 37.970 101.105 ;
        RECT 38.210 100.940 39.040 101.110 ;
        RECT 39.275 100.895 39.445 101.395 ;
        RECT 39.615 100.725 39.945 101.225 ;
        RECT 40.160 100.895 40.385 103.015 ;
        RECT 40.555 102.895 40.885 103.275 ;
        RECT 41.055 102.725 41.225 103.015 ;
        RECT 40.560 102.555 41.225 102.725 ;
        RECT 40.560 101.565 40.790 102.555 ;
        RECT 41.545 102.455 41.755 103.275 ;
        RECT 41.925 102.475 42.255 103.105 ;
        RECT 40.960 101.735 41.310 102.385 ;
        RECT 41.925 101.875 42.175 102.475 ;
        RECT 42.425 102.455 42.655 103.275 ;
        RECT 43.875 102.725 44.045 103.015 ;
        RECT 44.215 102.895 44.545 103.275 ;
        RECT 43.875 102.555 44.540 102.725 ;
        RECT 42.345 102.035 42.675 102.285 ;
        RECT 40.560 101.395 41.225 101.565 ;
        RECT 40.555 100.725 40.885 101.225 ;
        RECT 41.055 100.895 41.225 101.395 ;
        RECT 41.545 100.725 41.755 101.865 ;
        RECT 41.925 100.895 42.255 101.875 ;
        RECT 42.425 100.725 42.655 101.865 ;
        RECT 43.790 101.735 44.140 102.385 ;
        RECT 44.310 101.565 44.540 102.555 ;
        RECT 43.875 101.395 44.540 101.565 ;
        RECT 43.875 100.895 44.045 101.395 ;
        RECT 44.215 100.725 44.545 101.225 ;
        RECT 44.715 100.895 44.940 103.015 ;
        RECT 45.155 102.895 45.485 103.275 ;
        RECT 45.655 102.725 45.825 103.055 ;
        RECT 46.125 102.895 47.140 103.095 ;
        RECT 45.130 102.535 45.825 102.725 ;
        RECT 45.130 101.565 45.300 102.535 ;
        RECT 45.470 101.735 45.880 102.355 ;
        RECT 46.050 101.785 46.270 102.655 ;
        RECT 46.450 102.345 46.800 102.715 ;
        RECT 46.970 102.165 47.140 102.895 ;
        RECT 47.310 102.835 47.720 103.275 ;
        RECT 48.010 102.635 48.260 103.065 ;
        RECT 48.460 102.815 48.780 103.275 ;
        RECT 49.340 102.885 50.190 103.055 ;
        RECT 47.310 102.295 47.720 102.625 ;
        RECT 48.010 102.295 48.430 102.635 ;
        RECT 46.720 102.125 47.140 102.165 ;
        RECT 46.720 101.955 48.070 102.125 ;
        RECT 45.130 101.395 45.825 101.565 ;
        RECT 46.050 101.405 46.550 101.785 ;
        RECT 45.155 100.725 45.485 101.225 ;
        RECT 45.655 100.895 45.825 101.395 ;
        RECT 46.720 101.110 46.890 101.955 ;
        RECT 47.820 101.795 48.070 101.955 ;
        RECT 47.060 101.525 47.310 101.785 ;
        RECT 48.240 101.525 48.430 102.295 ;
        RECT 47.060 101.275 48.430 101.525 ;
        RECT 48.600 102.465 49.850 102.635 ;
        RECT 48.600 101.705 48.770 102.465 ;
        RECT 49.520 102.345 49.850 102.465 ;
        RECT 48.940 101.885 49.120 102.295 ;
        RECT 50.020 102.125 50.190 102.885 ;
        RECT 50.390 102.795 51.050 103.275 ;
        RECT 51.230 102.680 51.550 103.010 ;
        RECT 50.380 102.355 51.040 102.625 ;
        RECT 50.380 102.295 50.710 102.355 ;
        RECT 50.860 102.125 51.190 102.185 ;
        RECT 49.290 101.955 51.190 102.125 ;
        RECT 48.600 101.395 49.120 101.705 ;
        RECT 49.290 101.445 49.460 101.955 ;
        RECT 51.360 101.785 51.550 102.680 ;
        RECT 49.630 101.615 51.550 101.785 ;
        RECT 51.230 101.595 51.550 101.615 ;
        RECT 51.750 102.365 52.000 103.015 ;
        RECT 52.180 102.815 52.465 103.275 ;
        RECT 52.645 102.565 52.900 103.095 ;
        RECT 51.750 102.035 52.550 102.365 ;
        RECT 49.290 101.275 50.500 101.445 ;
        RECT 46.060 100.940 46.890 101.110 ;
        RECT 47.130 100.725 47.510 101.105 ;
        RECT 47.690 100.985 47.860 101.275 ;
        RECT 49.290 101.195 49.460 101.275 ;
        RECT 48.030 100.725 48.360 101.105 ;
        RECT 48.830 100.945 49.460 101.195 ;
        RECT 49.640 100.725 50.060 101.105 ;
        RECT 50.260 100.985 50.500 101.275 ;
        RECT 50.730 100.725 51.060 101.415 ;
        RECT 51.230 100.985 51.400 101.595 ;
        RECT 51.750 101.445 52.000 102.035 ;
        RECT 52.720 101.705 52.900 102.565 ;
        RECT 53.535 102.725 53.705 103.105 ;
        RECT 53.885 102.895 54.215 103.275 ;
        RECT 53.535 102.555 54.200 102.725 ;
        RECT 54.395 102.600 54.655 103.105 ;
        RECT 53.465 102.005 53.795 102.375 ;
        RECT 54.030 102.300 54.200 102.555 ;
        RECT 54.030 101.970 54.315 102.300 ;
        RECT 54.030 101.825 54.200 101.970 ;
        RECT 51.670 100.935 52.000 101.445 ;
        RECT 52.180 100.725 52.465 101.525 ;
        RECT 52.645 101.235 52.900 101.705 ;
        RECT 53.535 101.655 54.200 101.825 ;
        RECT 54.485 101.800 54.655 102.600 ;
        RECT 54.825 102.505 56.495 103.275 ;
        RECT 57.125 102.550 57.415 103.275 ;
        RECT 57.585 102.505 60.175 103.275 ;
        RECT 54.825 101.985 55.575 102.505 ;
        RECT 55.745 101.815 56.495 102.335 ;
        RECT 57.585 101.985 58.795 102.505 ;
        RECT 60.385 102.455 60.615 103.275 ;
        RECT 60.785 102.475 61.115 103.105 ;
        RECT 52.645 101.065 52.985 101.235 ;
        RECT 52.645 101.035 52.900 101.065 ;
        RECT 53.535 100.895 53.705 101.655 ;
        RECT 53.885 100.725 54.215 101.485 ;
        RECT 54.385 100.895 54.655 101.800 ;
        RECT 54.825 100.725 56.495 101.815 ;
        RECT 57.125 100.725 57.415 101.890 ;
        RECT 58.965 101.815 60.175 102.335 ;
        RECT 60.365 102.035 60.695 102.285 ;
        RECT 60.865 101.875 61.115 102.475 ;
        RECT 61.285 102.455 61.495 103.275 ;
        RECT 61.730 102.535 61.985 103.105 ;
        RECT 62.155 102.875 62.485 103.275 ;
        RECT 62.910 102.740 63.440 103.105 ;
        RECT 63.630 102.935 63.905 103.105 ;
        RECT 63.625 102.765 63.905 102.935 ;
        RECT 62.910 102.705 63.085 102.740 ;
        RECT 62.155 102.535 63.085 102.705 ;
        RECT 57.585 100.725 60.175 101.815 ;
        RECT 60.385 100.725 60.615 101.865 ;
        RECT 60.785 100.895 61.115 101.875 ;
        RECT 61.730 101.865 61.900 102.535 ;
        RECT 62.155 102.365 62.325 102.535 ;
        RECT 62.070 102.035 62.325 102.365 ;
        RECT 62.550 102.035 62.745 102.365 ;
        RECT 61.285 100.725 61.495 101.865 ;
        RECT 61.730 100.895 62.065 101.865 ;
        RECT 62.235 100.725 62.405 101.865 ;
        RECT 62.575 101.065 62.745 102.035 ;
        RECT 62.915 101.405 63.085 102.535 ;
        RECT 63.255 101.745 63.425 102.545 ;
        RECT 63.630 101.945 63.905 102.765 ;
        RECT 64.075 101.745 64.265 103.105 ;
        RECT 64.445 102.740 64.955 103.275 ;
        RECT 65.175 102.465 65.420 103.070 ;
        RECT 65.955 102.725 66.125 103.015 ;
        RECT 66.295 102.895 66.625 103.275 ;
        RECT 65.955 102.555 66.620 102.725 ;
        RECT 64.465 102.295 65.695 102.465 ;
        RECT 63.255 101.575 64.265 101.745 ;
        RECT 64.435 101.730 65.185 101.920 ;
        RECT 62.915 101.235 64.040 101.405 ;
        RECT 64.435 101.065 64.605 101.730 ;
        RECT 65.355 101.485 65.695 102.295 ;
        RECT 65.870 101.735 66.220 102.385 ;
        RECT 66.390 101.565 66.620 102.555 ;
        RECT 62.575 100.895 64.605 101.065 ;
        RECT 64.775 100.725 64.945 101.485 ;
        RECT 65.180 101.075 65.695 101.485 ;
        RECT 65.955 101.395 66.620 101.565 ;
        RECT 65.955 100.895 66.125 101.395 ;
        RECT 66.295 100.725 66.625 101.225 ;
        RECT 66.795 100.895 67.020 103.015 ;
        RECT 67.235 102.895 67.565 103.275 ;
        RECT 67.735 102.725 67.905 103.055 ;
        RECT 68.205 102.895 69.220 103.095 ;
        RECT 67.210 102.535 67.905 102.725 ;
        RECT 67.210 101.565 67.380 102.535 ;
        RECT 67.550 101.735 67.960 102.355 ;
        RECT 68.130 101.785 68.350 102.655 ;
        RECT 68.530 102.345 68.880 102.715 ;
        RECT 69.050 102.165 69.220 102.895 ;
        RECT 69.390 102.835 69.800 103.275 ;
        RECT 70.090 102.635 70.340 103.065 ;
        RECT 70.540 102.815 70.860 103.275 ;
        RECT 71.420 102.885 72.270 103.055 ;
        RECT 69.390 102.295 69.800 102.625 ;
        RECT 70.090 102.295 70.510 102.635 ;
        RECT 68.800 102.125 69.220 102.165 ;
        RECT 68.800 101.955 70.150 102.125 ;
        RECT 67.210 101.395 67.905 101.565 ;
        RECT 68.130 101.405 68.630 101.785 ;
        RECT 67.235 100.725 67.565 101.225 ;
        RECT 67.735 100.895 67.905 101.395 ;
        RECT 68.800 101.110 68.970 101.955 ;
        RECT 69.900 101.795 70.150 101.955 ;
        RECT 69.140 101.525 69.390 101.785 ;
        RECT 70.320 101.525 70.510 102.295 ;
        RECT 69.140 101.275 70.510 101.525 ;
        RECT 70.680 102.465 71.930 102.635 ;
        RECT 70.680 101.705 70.850 102.465 ;
        RECT 71.600 102.345 71.930 102.465 ;
        RECT 71.020 101.885 71.200 102.295 ;
        RECT 72.100 102.125 72.270 102.885 ;
        RECT 72.470 102.795 73.130 103.275 ;
        RECT 73.310 102.680 73.630 103.010 ;
        RECT 72.460 102.355 73.120 102.625 ;
        RECT 72.460 102.295 72.790 102.355 ;
        RECT 72.940 102.125 73.270 102.185 ;
        RECT 71.370 101.955 73.270 102.125 ;
        RECT 70.680 101.395 71.200 101.705 ;
        RECT 71.370 101.445 71.540 101.955 ;
        RECT 73.440 101.785 73.630 102.680 ;
        RECT 71.710 101.615 73.630 101.785 ;
        RECT 73.310 101.595 73.630 101.615 ;
        RECT 73.830 102.365 74.080 103.015 ;
        RECT 74.260 102.815 74.545 103.275 ;
        RECT 74.725 102.565 74.980 103.095 ;
        RECT 73.830 102.035 74.630 102.365 ;
        RECT 71.370 101.275 72.580 101.445 ;
        RECT 68.140 100.940 68.970 101.110 ;
        RECT 69.210 100.725 69.590 101.105 ;
        RECT 69.770 100.985 69.940 101.275 ;
        RECT 71.370 101.195 71.540 101.275 ;
        RECT 70.110 100.725 70.440 101.105 ;
        RECT 70.910 100.945 71.540 101.195 ;
        RECT 71.720 100.725 72.140 101.105 ;
        RECT 72.340 100.985 72.580 101.275 ;
        RECT 72.810 100.725 73.140 101.415 ;
        RECT 73.310 100.985 73.480 101.595 ;
        RECT 73.830 101.445 74.080 102.035 ;
        RECT 74.800 101.705 74.980 102.565 ;
        RECT 75.615 102.625 75.785 103.105 ;
        RECT 75.965 102.795 76.205 103.275 ;
        RECT 76.455 102.625 76.625 103.105 ;
        RECT 76.795 102.795 77.125 103.275 ;
        RECT 77.295 102.625 77.465 103.105 ;
        RECT 75.615 102.455 76.250 102.625 ;
        RECT 76.455 102.455 77.465 102.625 ;
        RECT 77.635 102.475 77.965 103.275 ;
        RECT 78.285 102.525 79.495 103.275 ;
        RECT 79.755 102.725 79.925 103.105 ;
        RECT 80.105 102.895 80.435 103.275 ;
        RECT 79.755 102.555 80.420 102.725 ;
        RECT 80.615 102.600 80.875 103.105 ;
        RECT 76.080 102.285 76.250 102.455 ;
        RECT 76.965 102.425 77.465 102.455 ;
        RECT 75.530 102.045 75.910 102.285 ;
        RECT 76.080 102.115 76.580 102.285 ;
        RECT 76.080 101.875 76.250 102.115 ;
        RECT 76.970 101.915 77.465 102.425 ;
        RECT 78.285 101.985 78.805 102.525 ;
        RECT 73.750 100.935 74.080 101.445 ;
        RECT 74.260 100.725 74.545 101.525 ;
        RECT 74.725 101.235 74.980 101.705 ;
        RECT 75.535 101.705 76.250 101.875 ;
        RECT 76.455 101.745 77.465 101.915 ;
        RECT 74.725 101.065 75.065 101.235 ;
        RECT 74.725 101.035 74.980 101.065 ;
        RECT 75.535 100.895 75.865 101.705 ;
        RECT 76.035 100.725 76.275 101.525 ;
        RECT 76.455 100.895 76.625 101.745 ;
        RECT 76.795 100.725 77.125 101.525 ;
        RECT 77.295 100.895 77.465 101.745 ;
        RECT 77.635 100.725 77.965 101.875 ;
        RECT 78.975 101.815 79.495 102.355 ;
        RECT 79.685 102.005 80.015 102.375 ;
        RECT 80.250 102.300 80.420 102.555 ;
        RECT 80.250 101.970 80.535 102.300 ;
        RECT 80.250 101.825 80.420 101.970 ;
        RECT 78.285 100.725 79.495 101.815 ;
        RECT 79.755 101.655 80.420 101.825 ;
        RECT 80.705 101.800 80.875 102.600 ;
        RECT 81.545 102.455 81.775 103.275 ;
        RECT 81.945 102.475 82.275 103.105 ;
        RECT 81.525 102.035 81.855 102.285 ;
        RECT 82.025 101.875 82.275 102.475 ;
        RECT 82.445 102.455 82.655 103.275 ;
        RECT 82.885 102.550 83.175 103.275 ;
        RECT 83.345 102.525 84.555 103.275 ;
        RECT 84.815 102.725 84.985 103.105 ;
        RECT 85.165 102.895 85.495 103.275 ;
        RECT 84.815 102.555 85.480 102.725 ;
        RECT 85.675 102.600 85.935 103.105 ;
        RECT 83.345 101.985 83.865 102.525 ;
        RECT 79.755 100.895 79.925 101.655 ;
        RECT 80.105 100.725 80.435 101.485 ;
        RECT 80.605 100.895 80.875 101.800 ;
        RECT 81.545 100.725 81.775 101.865 ;
        RECT 81.945 100.895 82.275 101.875 ;
        RECT 82.445 100.725 82.655 101.865 ;
        RECT 82.885 100.725 83.175 101.890 ;
        RECT 84.035 101.815 84.555 102.355 ;
        RECT 84.745 102.005 85.075 102.375 ;
        RECT 85.310 102.300 85.480 102.555 ;
        RECT 85.310 101.970 85.595 102.300 ;
        RECT 85.310 101.825 85.480 101.970 ;
        RECT 83.345 100.725 84.555 101.815 ;
        RECT 84.815 101.655 85.480 101.825 ;
        RECT 85.765 101.800 85.935 102.600 ;
        RECT 86.195 102.725 86.365 103.015 ;
        RECT 86.535 102.895 86.865 103.275 ;
        RECT 86.195 102.555 86.860 102.725 ;
        RECT 84.815 100.895 84.985 101.655 ;
        RECT 85.165 100.725 85.495 101.485 ;
        RECT 85.665 100.895 85.935 101.800 ;
        RECT 86.110 101.735 86.460 102.385 ;
        RECT 86.630 101.565 86.860 102.555 ;
        RECT 86.195 101.395 86.860 101.565 ;
        RECT 86.195 100.895 86.365 101.395 ;
        RECT 86.535 100.725 86.865 101.225 ;
        RECT 87.035 100.895 87.260 103.015 ;
        RECT 87.475 102.895 87.805 103.275 ;
        RECT 87.975 102.725 88.145 103.055 ;
        RECT 88.445 102.895 89.460 103.095 ;
        RECT 87.450 102.535 88.145 102.725 ;
        RECT 87.450 101.565 87.620 102.535 ;
        RECT 87.790 101.735 88.200 102.355 ;
        RECT 88.370 101.785 88.590 102.655 ;
        RECT 88.770 102.345 89.120 102.715 ;
        RECT 89.290 102.165 89.460 102.895 ;
        RECT 89.630 102.835 90.040 103.275 ;
        RECT 90.330 102.635 90.580 103.065 ;
        RECT 90.780 102.815 91.100 103.275 ;
        RECT 91.660 102.885 92.510 103.055 ;
        RECT 89.630 102.295 90.040 102.625 ;
        RECT 90.330 102.295 90.750 102.635 ;
        RECT 89.040 102.125 89.460 102.165 ;
        RECT 89.040 101.955 90.390 102.125 ;
        RECT 87.450 101.395 88.145 101.565 ;
        RECT 88.370 101.405 88.870 101.785 ;
        RECT 87.475 100.725 87.805 101.225 ;
        RECT 87.975 100.895 88.145 101.395 ;
        RECT 89.040 101.110 89.210 101.955 ;
        RECT 90.140 101.795 90.390 101.955 ;
        RECT 89.380 101.525 89.630 101.785 ;
        RECT 90.560 101.525 90.750 102.295 ;
        RECT 89.380 101.275 90.750 101.525 ;
        RECT 90.920 102.465 92.170 102.635 ;
        RECT 90.920 101.705 91.090 102.465 ;
        RECT 91.840 102.345 92.170 102.465 ;
        RECT 91.260 101.885 91.440 102.295 ;
        RECT 92.340 102.125 92.510 102.885 ;
        RECT 92.710 102.795 93.370 103.275 ;
        RECT 93.550 102.680 93.870 103.010 ;
        RECT 92.700 102.355 93.360 102.625 ;
        RECT 92.700 102.295 93.030 102.355 ;
        RECT 93.180 102.125 93.510 102.185 ;
        RECT 91.610 101.955 93.510 102.125 ;
        RECT 90.920 101.395 91.440 101.705 ;
        RECT 91.610 101.445 91.780 101.955 ;
        RECT 93.680 101.785 93.870 102.680 ;
        RECT 91.950 101.615 93.870 101.785 ;
        RECT 93.550 101.595 93.870 101.615 ;
        RECT 94.070 102.365 94.320 103.015 ;
        RECT 94.500 102.815 94.785 103.275 ;
        RECT 94.965 102.565 95.220 103.095 ;
        RECT 96.225 102.765 96.530 103.275 ;
        RECT 94.070 102.035 94.870 102.365 ;
        RECT 91.610 101.275 92.820 101.445 ;
        RECT 88.380 100.940 89.210 101.110 ;
        RECT 89.450 100.725 89.830 101.105 ;
        RECT 90.010 100.985 90.180 101.275 ;
        RECT 91.610 101.195 91.780 101.275 ;
        RECT 90.350 100.725 90.680 101.105 ;
        RECT 91.150 100.945 91.780 101.195 ;
        RECT 91.960 100.725 92.380 101.105 ;
        RECT 92.580 100.985 92.820 101.275 ;
        RECT 93.050 100.725 93.380 101.415 ;
        RECT 93.550 100.985 93.720 101.595 ;
        RECT 94.070 101.445 94.320 102.035 ;
        RECT 95.040 101.705 95.220 102.565 ;
        RECT 96.225 102.035 96.540 102.595 ;
        RECT 96.710 102.285 96.960 103.095 ;
        RECT 97.130 102.750 97.390 103.275 ;
        RECT 97.570 102.285 97.820 103.095 ;
        RECT 97.990 102.715 98.250 103.275 ;
        RECT 98.420 102.625 98.680 103.080 ;
        RECT 98.850 102.795 99.110 103.275 ;
        RECT 99.280 102.625 99.540 103.080 ;
        RECT 99.710 102.795 99.970 103.275 ;
        RECT 100.140 102.625 100.400 103.080 ;
        RECT 100.570 102.795 100.815 103.275 ;
        RECT 100.985 102.625 101.260 103.080 ;
        RECT 101.430 102.795 101.675 103.275 ;
        RECT 101.845 102.625 102.105 103.080 ;
        RECT 102.285 102.795 102.535 103.275 ;
        RECT 102.705 102.625 102.965 103.080 ;
        RECT 103.145 102.795 103.395 103.275 ;
        RECT 103.565 102.625 103.825 103.080 ;
        RECT 104.005 102.795 104.265 103.275 ;
        RECT 104.435 102.625 104.695 103.080 ;
        RECT 104.865 102.795 105.165 103.275 ;
        RECT 98.420 102.455 105.165 102.625 ;
        RECT 96.710 102.035 103.830 102.285 ;
        RECT 93.990 100.935 94.320 101.445 ;
        RECT 94.500 100.725 94.785 101.525 ;
        RECT 94.965 101.235 95.220 101.705 ;
        RECT 94.965 101.065 95.305 101.235 ;
        RECT 94.965 101.035 95.220 101.065 ;
        RECT 96.235 100.725 96.530 101.535 ;
        RECT 96.710 100.895 96.955 102.035 ;
        RECT 97.130 100.725 97.390 101.535 ;
        RECT 97.570 100.900 97.820 102.035 ;
        RECT 104.000 101.865 105.165 102.455 ;
        RECT 98.420 101.640 105.165 101.865 ;
        RECT 105.425 102.600 105.685 103.105 ;
        RECT 105.865 102.895 106.195 103.275 ;
        RECT 106.375 102.725 106.545 103.105 ;
        RECT 105.425 101.800 105.595 102.600 ;
        RECT 105.880 102.555 106.545 102.725 ;
        RECT 105.880 102.300 106.050 102.555 ;
        RECT 106.845 102.455 107.075 103.275 ;
        RECT 107.245 102.475 107.575 103.105 ;
        RECT 105.765 101.970 106.050 102.300 ;
        RECT 106.285 102.005 106.615 102.375 ;
        RECT 106.825 102.035 107.155 102.285 ;
        RECT 105.880 101.825 106.050 101.970 ;
        RECT 107.325 101.875 107.575 102.475 ;
        RECT 107.745 102.455 107.955 103.275 ;
        RECT 108.645 102.550 108.935 103.275 ;
        RECT 109.105 102.505 111.695 103.275 ;
        RECT 112.325 102.525 113.535 103.275 ;
        RECT 109.105 101.985 110.315 102.505 ;
        RECT 98.420 101.625 103.825 101.640 ;
        RECT 97.990 100.730 98.250 101.525 ;
        RECT 98.420 100.900 98.680 101.625 ;
        RECT 98.850 100.730 99.110 101.455 ;
        RECT 99.280 100.900 99.540 101.625 ;
        RECT 99.710 100.730 99.970 101.455 ;
        RECT 100.140 100.900 100.400 101.625 ;
        RECT 100.570 100.730 100.830 101.455 ;
        RECT 101.000 100.900 101.260 101.625 ;
        RECT 101.430 100.730 101.675 101.455 ;
        RECT 101.845 100.900 102.105 101.625 ;
        RECT 102.290 100.730 102.535 101.455 ;
        RECT 102.705 100.900 102.965 101.625 ;
        RECT 103.150 100.730 103.395 101.455 ;
        RECT 103.565 100.900 103.825 101.625 ;
        RECT 104.010 100.730 104.265 101.455 ;
        RECT 104.435 100.900 104.725 101.640 ;
        RECT 97.990 100.725 104.265 100.730 ;
        RECT 104.895 100.725 105.165 101.470 ;
        RECT 105.425 100.895 105.695 101.800 ;
        RECT 105.880 101.655 106.545 101.825 ;
        RECT 105.865 100.725 106.195 101.485 ;
        RECT 106.375 100.895 106.545 101.655 ;
        RECT 106.845 100.725 107.075 101.865 ;
        RECT 107.245 100.895 107.575 101.875 ;
        RECT 107.745 100.725 107.955 101.865 ;
        RECT 108.645 100.725 108.935 101.890 ;
        RECT 110.485 101.815 111.695 102.335 ;
        RECT 109.105 100.725 111.695 101.815 ;
        RECT 112.325 101.815 112.845 102.355 ;
        RECT 113.015 101.985 113.535 102.525 ;
        RECT 112.325 100.725 113.535 101.815 ;
        RECT 5.520 100.555 113.620 100.725 ;
        RECT 5.605 99.465 6.815 100.555 ;
        RECT 7.995 99.885 8.165 100.385 ;
        RECT 8.335 100.055 8.665 100.555 ;
        RECT 7.995 99.715 8.660 99.885 ;
        RECT 5.605 98.755 6.125 99.295 ;
        RECT 6.295 98.925 6.815 99.465 ;
        RECT 7.910 98.895 8.260 99.545 ;
        RECT 5.605 98.005 6.815 98.755 ;
        RECT 8.430 98.725 8.660 99.715 ;
        RECT 7.995 98.555 8.660 98.725 ;
        RECT 7.995 98.265 8.165 98.555 ;
        RECT 8.335 98.005 8.665 98.385 ;
        RECT 8.835 98.265 9.060 100.385 ;
        RECT 9.275 100.055 9.605 100.555 ;
        RECT 9.775 99.885 9.945 100.385 ;
        RECT 10.180 100.170 11.010 100.340 ;
        RECT 11.250 100.175 11.630 100.555 ;
        RECT 9.250 99.715 9.945 99.885 ;
        RECT 9.250 98.745 9.420 99.715 ;
        RECT 9.590 98.925 10.000 99.545 ;
        RECT 10.170 99.495 10.670 99.875 ;
        RECT 9.250 98.555 9.945 98.745 ;
        RECT 10.170 98.625 10.390 99.495 ;
        RECT 10.840 99.325 11.010 100.170 ;
        RECT 11.810 100.005 11.980 100.295 ;
        RECT 12.150 100.175 12.480 100.555 ;
        RECT 12.950 100.085 13.580 100.335 ;
        RECT 13.760 100.175 14.180 100.555 ;
        RECT 13.410 100.005 13.580 100.085 ;
        RECT 14.380 100.005 14.620 100.295 ;
        RECT 11.180 99.755 12.550 100.005 ;
        RECT 11.180 99.495 11.430 99.755 ;
        RECT 11.940 99.325 12.190 99.485 ;
        RECT 10.840 99.155 12.190 99.325 ;
        RECT 10.840 99.115 11.260 99.155 ;
        RECT 10.570 98.565 10.920 98.935 ;
        RECT 9.275 98.005 9.605 98.385 ;
        RECT 9.775 98.225 9.945 98.555 ;
        RECT 11.090 98.385 11.260 99.115 ;
        RECT 12.360 98.985 12.550 99.755 ;
        RECT 11.430 98.655 11.840 98.985 ;
        RECT 12.130 98.645 12.550 98.985 ;
        RECT 12.720 99.575 13.240 99.885 ;
        RECT 13.410 99.835 14.620 100.005 ;
        RECT 14.850 99.865 15.180 100.555 ;
        RECT 12.720 98.815 12.890 99.575 ;
        RECT 13.060 98.985 13.240 99.395 ;
        RECT 13.410 99.325 13.580 99.835 ;
        RECT 15.350 99.685 15.520 100.295 ;
        RECT 15.790 99.835 16.120 100.345 ;
        RECT 15.350 99.665 15.670 99.685 ;
        RECT 13.750 99.495 15.670 99.665 ;
        RECT 13.410 99.155 15.310 99.325 ;
        RECT 13.640 98.815 13.970 98.935 ;
        RECT 12.720 98.645 13.970 98.815 ;
        RECT 10.245 98.185 11.260 98.385 ;
        RECT 11.430 98.005 11.840 98.445 ;
        RECT 12.130 98.215 12.380 98.645 ;
        RECT 12.580 98.005 12.900 98.465 ;
        RECT 14.140 98.395 14.310 99.155 ;
        RECT 14.980 99.095 15.310 99.155 ;
        RECT 14.500 98.925 14.830 98.985 ;
        RECT 14.500 98.655 15.160 98.925 ;
        RECT 15.480 98.600 15.670 99.495 ;
        RECT 13.460 98.225 14.310 98.395 ;
        RECT 14.510 98.005 15.170 98.485 ;
        RECT 15.350 98.270 15.670 98.600 ;
        RECT 15.870 99.245 16.120 99.835 ;
        RECT 16.300 99.755 16.585 100.555 ;
        RECT 16.765 99.575 17.020 100.245 ;
        RECT 15.870 98.915 16.670 99.245 ;
        RECT 16.840 99.195 17.020 99.575 ;
        RECT 18.485 99.390 18.775 100.555 ;
        RECT 18.950 99.415 19.285 100.385 ;
        RECT 19.455 99.415 19.625 100.555 ;
        RECT 19.795 100.215 21.825 100.385 ;
        RECT 16.840 99.025 17.105 99.195 ;
        RECT 15.870 98.265 16.120 98.915 ;
        RECT 16.840 98.715 17.020 99.025 ;
        RECT 18.950 98.745 19.120 99.415 ;
        RECT 19.795 99.245 19.965 100.215 ;
        RECT 19.290 98.915 19.545 99.245 ;
        RECT 19.770 98.915 19.965 99.245 ;
        RECT 20.135 99.875 21.260 100.045 ;
        RECT 19.375 98.745 19.545 98.915 ;
        RECT 20.135 98.745 20.305 99.875 ;
        RECT 16.300 98.005 16.585 98.465 ;
        RECT 16.765 98.185 17.020 98.715 ;
        RECT 18.485 98.005 18.775 98.730 ;
        RECT 18.950 98.175 19.205 98.745 ;
        RECT 19.375 98.575 20.305 98.745 ;
        RECT 20.475 99.535 21.485 99.705 ;
        RECT 20.475 98.735 20.645 99.535 ;
        RECT 20.850 98.855 21.125 99.335 ;
        RECT 20.845 98.685 21.125 98.855 ;
        RECT 20.130 98.540 20.305 98.575 ;
        RECT 19.375 98.005 19.705 98.405 ;
        RECT 20.130 98.175 20.660 98.540 ;
        RECT 20.850 98.175 21.125 98.685 ;
        RECT 21.295 98.175 21.485 99.535 ;
        RECT 21.655 99.550 21.825 100.215 ;
        RECT 21.995 99.795 22.165 100.555 ;
        RECT 22.400 99.795 22.915 100.205 ;
        RECT 21.655 99.360 22.405 99.550 ;
        RECT 22.575 98.985 22.915 99.795 ;
        RECT 23.145 99.415 23.355 100.555 ;
        RECT 21.685 98.815 22.915 98.985 ;
        RECT 23.525 99.405 23.855 100.385 ;
        RECT 24.025 99.415 24.255 100.555 ;
        RECT 25.385 99.480 25.655 100.385 ;
        RECT 25.825 99.795 26.155 100.555 ;
        RECT 26.335 99.625 26.505 100.385 ;
        RECT 21.665 98.005 22.175 98.540 ;
        RECT 22.395 98.210 22.640 98.815 ;
        RECT 23.145 98.005 23.355 98.825 ;
        RECT 23.525 98.805 23.775 99.405 ;
        RECT 23.945 98.995 24.275 99.245 ;
        RECT 23.525 98.175 23.855 98.805 ;
        RECT 24.025 98.005 24.255 98.825 ;
        RECT 25.385 98.680 25.555 99.480 ;
        RECT 25.840 99.455 26.505 99.625 ;
        RECT 25.840 99.310 26.010 99.455 ;
        RECT 25.725 98.980 26.010 99.310 ;
        RECT 26.770 99.415 27.105 100.385 ;
        RECT 27.275 99.415 27.445 100.555 ;
        RECT 27.615 100.215 29.645 100.385 ;
        RECT 25.840 98.725 26.010 98.980 ;
        RECT 26.245 98.905 26.575 99.275 ;
        RECT 26.770 98.745 26.940 99.415 ;
        RECT 27.615 99.245 27.785 100.215 ;
        RECT 27.110 98.915 27.365 99.245 ;
        RECT 27.590 98.915 27.785 99.245 ;
        RECT 27.955 99.875 29.080 100.045 ;
        RECT 27.195 98.745 27.365 98.915 ;
        RECT 27.955 98.745 28.125 99.875 ;
        RECT 25.385 98.175 25.645 98.680 ;
        RECT 25.840 98.555 26.505 98.725 ;
        RECT 25.825 98.005 26.155 98.385 ;
        RECT 26.335 98.175 26.505 98.555 ;
        RECT 26.770 98.175 27.025 98.745 ;
        RECT 27.195 98.575 28.125 98.745 ;
        RECT 28.295 99.535 29.305 99.705 ;
        RECT 28.295 98.735 28.465 99.535 ;
        RECT 28.670 99.195 28.945 99.335 ;
        RECT 28.665 99.025 28.945 99.195 ;
        RECT 27.950 98.540 28.125 98.575 ;
        RECT 27.195 98.005 27.525 98.405 ;
        RECT 27.950 98.175 28.480 98.540 ;
        RECT 28.670 98.175 28.945 99.025 ;
        RECT 29.115 98.175 29.305 99.535 ;
        RECT 29.475 99.550 29.645 100.215 ;
        RECT 29.815 99.795 29.985 100.555 ;
        RECT 30.220 99.795 30.735 100.205 ;
        RECT 29.475 99.360 30.225 99.550 ;
        RECT 30.395 98.985 30.735 99.795 ;
        RECT 31.455 99.625 31.625 100.385 ;
        RECT 31.805 99.795 32.135 100.555 ;
        RECT 31.455 99.455 32.120 99.625 ;
        RECT 32.305 99.480 32.575 100.385 ;
        RECT 32.835 99.885 33.005 100.385 ;
        RECT 33.175 100.055 33.505 100.555 ;
        RECT 32.835 99.715 33.500 99.885 ;
        RECT 31.950 99.310 32.120 99.455 ;
        RECT 29.505 98.815 30.735 98.985 ;
        RECT 31.385 98.905 31.715 99.275 ;
        RECT 31.950 98.980 32.235 99.310 ;
        RECT 29.485 98.005 29.995 98.540 ;
        RECT 30.215 98.210 30.460 98.815 ;
        RECT 31.950 98.725 32.120 98.980 ;
        RECT 31.455 98.555 32.120 98.725 ;
        RECT 32.405 98.680 32.575 99.480 ;
        RECT 32.750 98.895 33.100 99.545 ;
        RECT 33.270 98.725 33.500 99.715 ;
        RECT 31.455 98.175 31.625 98.555 ;
        RECT 31.805 98.005 32.135 98.385 ;
        RECT 32.315 98.175 32.575 98.680 ;
        RECT 32.835 98.555 33.500 98.725 ;
        RECT 32.835 98.265 33.005 98.555 ;
        RECT 33.175 98.005 33.505 98.385 ;
        RECT 33.675 98.265 33.900 100.385 ;
        RECT 34.115 100.055 34.445 100.555 ;
        RECT 34.615 99.885 34.785 100.385 ;
        RECT 35.020 100.170 35.850 100.340 ;
        RECT 36.090 100.175 36.470 100.555 ;
        RECT 34.090 99.715 34.785 99.885 ;
        RECT 34.090 98.745 34.260 99.715 ;
        RECT 34.430 98.925 34.840 99.545 ;
        RECT 35.010 99.495 35.510 99.875 ;
        RECT 34.090 98.555 34.785 98.745 ;
        RECT 35.010 98.625 35.230 99.495 ;
        RECT 35.680 99.325 35.850 100.170 ;
        RECT 36.650 100.005 36.820 100.295 ;
        RECT 36.990 100.175 37.320 100.555 ;
        RECT 37.790 100.085 38.420 100.335 ;
        RECT 38.600 100.175 39.020 100.555 ;
        RECT 38.250 100.005 38.420 100.085 ;
        RECT 39.220 100.005 39.460 100.295 ;
        RECT 36.020 99.755 37.390 100.005 ;
        RECT 36.020 99.495 36.270 99.755 ;
        RECT 36.780 99.325 37.030 99.485 ;
        RECT 35.680 99.155 37.030 99.325 ;
        RECT 35.680 99.115 36.100 99.155 ;
        RECT 35.410 98.565 35.760 98.935 ;
        RECT 34.115 98.005 34.445 98.385 ;
        RECT 34.615 98.225 34.785 98.555 ;
        RECT 35.930 98.385 36.100 99.115 ;
        RECT 37.200 98.985 37.390 99.755 ;
        RECT 36.270 98.655 36.680 98.985 ;
        RECT 36.970 98.645 37.390 98.985 ;
        RECT 37.560 99.575 38.080 99.885 ;
        RECT 38.250 99.835 39.460 100.005 ;
        RECT 39.690 99.865 40.020 100.555 ;
        RECT 37.560 98.815 37.730 99.575 ;
        RECT 37.900 98.985 38.080 99.395 ;
        RECT 38.250 99.325 38.420 99.835 ;
        RECT 40.190 99.685 40.360 100.295 ;
        RECT 40.630 99.835 40.960 100.345 ;
        RECT 40.190 99.665 40.510 99.685 ;
        RECT 38.590 99.495 40.510 99.665 ;
        RECT 38.250 99.155 40.150 99.325 ;
        RECT 38.480 98.815 38.810 98.935 ;
        RECT 37.560 98.645 38.810 98.815 ;
        RECT 35.085 98.185 36.100 98.385 ;
        RECT 36.270 98.005 36.680 98.445 ;
        RECT 36.970 98.215 37.220 98.645 ;
        RECT 37.420 98.005 37.740 98.465 ;
        RECT 38.980 98.395 39.150 99.155 ;
        RECT 39.820 99.095 40.150 99.155 ;
        RECT 39.340 98.925 39.670 98.985 ;
        RECT 39.340 98.655 40.000 98.925 ;
        RECT 40.320 98.600 40.510 99.495 ;
        RECT 38.300 98.225 39.150 98.395 ;
        RECT 39.350 98.005 40.010 98.485 ;
        RECT 40.190 98.270 40.510 98.600 ;
        RECT 40.710 99.245 40.960 99.835 ;
        RECT 41.140 99.755 41.425 100.555 ;
        RECT 41.605 99.575 41.860 100.245 ;
        RECT 40.710 98.915 41.510 99.245 ;
        RECT 40.710 98.265 40.960 98.915 ;
        RECT 41.680 98.855 41.860 99.575 ;
        RECT 42.495 99.625 42.665 100.385 ;
        RECT 42.845 99.795 43.175 100.555 ;
        RECT 42.495 99.455 43.160 99.625 ;
        RECT 43.345 99.480 43.615 100.385 ;
        RECT 42.990 99.310 43.160 99.455 ;
        RECT 42.425 98.905 42.755 99.275 ;
        RECT 42.990 98.980 43.275 99.310 ;
        RECT 41.680 98.715 41.945 98.855 ;
        RECT 42.990 98.725 43.160 98.980 ;
        RECT 41.605 98.685 41.945 98.715 ;
        RECT 41.140 98.005 41.425 98.465 ;
        RECT 41.605 98.185 41.860 98.685 ;
        RECT 42.495 98.555 43.160 98.725 ;
        RECT 43.445 98.680 43.615 99.480 ;
        RECT 44.245 99.390 44.535 100.555 ;
        RECT 45.625 99.480 45.895 100.385 ;
        RECT 46.065 99.795 46.395 100.555 ;
        RECT 46.575 99.625 46.745 100.385 ;
        RECT 42.495 98.175 42.665 98.555 ;
        RECT 42.845 98.005 43.175 98.385 ;
        RECT 43.355 98.175 43.615 98.680 ;
        RECT 44.245 98.005 44.535 98.730 ;
        RECT 45.625 98.680 45.795 99.480 ;
        RECT 46.080 99.455 46.745 99.625 ;
        RECT 47.380 99.575 47.635 100.245 ;
        RECT 47.815 99.755 48.100 100.555 ;
        RECT 48.280 99.835 48.610 100.345 ;
        RECT 46.080 99.310 46.250 99.455 ;
        RECT 45.965 98.980 46.250 99.310 ;
        RECT 46.080 98.725 46.250 98.980 ;
        RECT 46.485 98.905 46.815 99.275 ;
        RECT 45.625 98.175 45.885 98.680 ;
        RECT 46.080 98.555 46.745 98.725 ;
        RECT 46.065 98.005 46.395 98.385 ;
        RECT 46.575 98.175 46.745 98.555 ;
        RECT 47.380 98.715 47.560 99.575 ;
        RECT 48.280 99.245 48.530 99.835 ;
        RECT 48.880 99.685 49.050 100.295 ;
        RECT 49.220 99.865 49.550 100.555 ;
        RECT 49.780 100.005 50.020 100.295 ;
        RECT 50.220 100.175 50.640 100.555 ;
        RECT 50.820 100.085 51.450 100.335 ;
        RECT 51.920 100.175 52.250 100.555 ;
        RECT 50.820 100.005 50.990 100.085 ;
        RECT 52.420 100.005 52.590 100.295 ;
        RECT 52.770 100.175 53.150 100.555 ;
        RECT 53.390 100.170 54.220 100.340 ;
        RECT 49.780 99.835 50.990 100.005 ;
        RECT 47.730 98.915 48.530 99.245 ;
        RECT 47.380 98.515 47.635 98.715 ;
        RECT 47.295 98.345 47.635 98.515 ;
        RECT 47.380 98.185 47.635 98.345 ;
        RECT 47.815 98.005 48.100 98.465 ;
        RECT 48.280 98.265 48.530 98.915 ;
        RECT 48.730 99.665 49.050 99.685 ;
        RECT 48.730 99.495 50.650 99.665 ;
        RECT 48.730 98.600 48.920 99.495 ;
        RECT 50.820 99.325 50.990 99.835 ;
        RECT 51.160 99.575 51.680 99.885 ;
        RECT 49.090 99.155 50.990 99.325 ;
        RECT 49.090 99.095 49.420 99.155 ;
        RECT 49.570 98.925 49.900 98.985 ;
        RECT 49.240 98.655 49.900 98.925 ;
        RECT 48.730 98.270 49.050 98.600 ;
        RECT 49.230 98.005 49.890 98.485 ;
        RECT 50.090 98.395 50.260 99.155 ;
        RECT 51.160 98.985 51.340 99.395 ;
        RECT 50.430 98.815 50.760 98.935 ;
        RECT 51.510 98.815 51.680 99.575 ;
        RECT 50.430 98.645 51.680 98.815 ;
        RECT 51.850 99.755 53.220 100.005 ;
        RECT 51.850 98.985 52.040 99.755 ;
        RECT 52.970 99.495 53.220 99.755 ;
        RECT 52.210 99.325 52.460 99.485 ;
        RECT 53.390 99.325 53.560 100.170 ;
        RECT 54.455 99.885 54.625 100.385 ;
        RECT 54.795 100.055 55.125 100.555 ;
        RECT 53.730 99.495 54.230 99.875 ;
        RECT 54.455 99.715 55.150 99.885 ;
        RECT 52.210 99.155 53.560 99.325 ;
        RECT 53.140 99.115 53.560 99.155 ;
        RECT 51.850 98.645 52.270 98.985 ;
        RECT 52.560 98.655 52.970 98.985 ;
        RECT 50.090 98.225 50.940 98.395 ;
        RECT 51.500 98.005 51.820 98.465 ;
        RECT 52.020 98.215 52.270 98.645 ;
        RECT 52.560 98.005 52.970 98.445 ;
        RECT 53.140 98.385 53.310 99.115 ;
        RECT 53.480 98.565 53.830 98.935 ;
        RECT 54.010 98.625 54.230 99.495 ;
        RECT 54.400 98.925 54.810 99.545 ;
        RECT 54.980 98.745 55.150 99.715 ;
        RECT 54.455 98.555 55.150 98.745 ;
        RECT 53.140 98.185 54.155 98.385 ;
        RECT 54.455 98.225 54.625 98.555 ;
        RECT 54.795 98.005 55.125 98.385 ;
        RECT 55.340 98.265 55.565 100.385 ;
        RECT 55.735 100.055 56.065 100.555 ;
        RECT 56.235 99.885 56.405 100.385 ;
        RECT 55.740 99.715 56.405 99.885 ;
        RECT 56.755 99.885 56.925 100.385 ;
        RECT 57.095 100.055 57.425 100.555 ;
        RECT 56.755 99.715 57.420 99.885 ;
        RECT 55.740 98.725 55.970 99.715 ;
        RECT 56.140 98.895 56.490 99.545 ;
        RECT 56.670 98.895 57.020 99.545 ;
        RECT 57.190 98.725 57.420 99.715 ;
        RECT 55.740 98.555 56.405 98.725 ;
        RECT 55.735 98.005 56.065 98.385 ;
        RECT 56.235 98.265 56.405 98.555 ;
        RECT 56.755 98.555 57.420 98.725 ;
        RECT 56.755 98.265 56.925 98.555 ;
        RECT 57.095 98.005 57.425 98.385 ;
        RECT 57.595 98.265 57.820 100.385 ;
        RECT 58.035 100.055 58.365 100.555 ;
        RECT 58.535 99.885 58.705 100.385 ;
        RECT 58.940 100.170 59.770 100.340 ;
        RECT 60.010 100.175 60.390 100.555 ;
        RECT 58.010 99.715 58.705 99.885 ;
        RECT 58.010 98.745 58.180 99.715 ;
        RECT 58.350 98.925 58.760 99.545 ;
        RECT 58.930 99.495 59.430 99.875 ;
        RECT 58.010 98.555 58.705 98.745 ;
        RECT 58.930 98.625 59.150 99.495 ;
        RECT 59.600 99.325 59.770 100.170 ;
        RECT 60.570 100.005 60.740 100.295 ;
        RECT 60.910 100.175 61.240 100.555 ;
        RECT 61.710 100.085 62.340 100.335 ;
        RECT 62.520 100.175 62.940 100.555 ;
        RECT 62.170 100.005 62.340 100.085 ;
        RECT 63.140 100.005 63.380 100.295 ;
        RECT 59.940 99.755 61.310 100.005 ;
        RECT 59.940 99.495 60.190 99.755 ;
        RECT 60.700 99.325 60.950 99.485 ;
        RECT 59.600 99.155 60.950 99.325 ;
        RECT 59.600 99.115 60.020 99.155 ;
        RECT 59.330 98.565 59.680 98.935 ;
        RECT 58.035 98.005 58.365 98.385 ;
        RECT 58.535 98.225 58.705 98.555 ;
        RECT 59.850 98.385 60.020 99.115 ;
        RECT 61.120 98.985 61.310 99.755 ;
        RECT 60.190 98.655 60.600 98.985 ;
        RECT 60.890 98.645 61.310 98.985 ;
        RECT 61.480 99.575 62.000 99.885 ;
        RECT 62.170 99.835 63.380 100.005 ;
        RECT 63.610 99.865 63.940 100.555 ;
        RECT 61.480 98.815 61.650 99.575 ;
        RECT 61.820 98.985 62.000 99.395 ;
        RECT 62.170 99.325 62.340 99.835 ;
        RECT 64.110 99.685 64.280 100.295 ;
        RECT 64.550 99.835 64.880 100.345 ;
        RECT 64.110 99.665 64.430 99.685 ;
        RECT 62.510 99.495 64.430 99.665 ;
        RECT 62.170 99.155 64.070 99.325 ;
        RECT 62.400 98.815 62.730 98.935 ;
        RECT 61.480 98.645 62.730 98.815 ;
        RECT 59.005 98.185 60.020 98.385 ;
        RECT 60.190 98.005 60.600 98.445 ;
        RECT 60.890 98.215 61.140 98.645 ;
        RECT 61.340 98.005 61.660 98.465 ;
        RECT 62.900 98.395 63.070 99.155 ;
        RECT 63.740 99.095 64.070 99.155 ;
        RECT 63.260 98.925 63.590 98.985 ;
        RECT 63.260 98.655 63.920 98.925 ;
        RECT 64.240 98.600 64.430 99.495 ;
        RECT 62.220 98.225 63.070 98.395 ;
        RECT 63.270 98.005 63.930 98.485 ;
        RECT 64.110 98.270 64.430 98.600 ;
        RECT 64.630 99.245 64.880 99.835 ;
        RECT 65.060 99.755 65.345 100.555 ;
        RECT 65.525 99.575 65.780 100.245 ;
        RECT 64.630 98.915 65.430 99.245 ;
        RECT 64.630 98.265 64.880 98.915 ;
        RECT 65.600 98.715 65.780 99.575 ;
        RECT 66.325 99.465 67.995 100.555 ;
        RECT 65.525 98.515 65.780 98.715 ;
        RECT 66.325 98.775 67.075 99.295 ;
        RECT 67.245 98.945 67.995 99.465 ;
        RECT 68.165 99.480 68.435 100.385 ;
        RECT 68.605 99.795 68.935 100.555 ;
        RECT 69.115 99.625 69.285 100.385 ;
        RECT 65.060 98.005 65.345 98.465 ;
        RECT 65.525 98.345 65.865 98.515 ;
        RECT 65.525 98.185 65.780 98.345 ;
        RECT 66.325 98.005 67.995 98.775 ;
        RECT 68.165 98.680 68.335 99.480 ;
        RECT 68.620 99.455 69.285 99.625 ;
        RECT 68.620 99.310 68.790 99.455 ;
        RECT 70.005 99.390 70.295 100.555 ;
        RECT 70.465 99.465 72.135 100.555 ;
        RECT 68.505 98.980 68.790 99.310 ;
        RECT 68.620 98.725 68.790 98.980 ;
        RECT 69.025 98.905 69.355 99.275 ;
        RECT 70.465 98.775 71.215 99.295 ;
        RECT 71.385 98.945 72.135 99.465 ;
        RECT 72.775 99.535 73.105 100.385 ;
        RECT 73.275 99.705 73.445 100.555 ;
        RECT 73.615 99.535 73.945 100.385 ;
        RECT 74.115 99.705 74.285 100.555 ;
        RECT 74.455 99.535 74.785 100.385 ;
        RECT 74.955 99.755 75.125 100.555 ;
        RECT 75.295 99.535 75.625 100.385 ;
        RECT 75.795 99.755 75.965 100.555 ;
        RECT 76.135 99.535 76.465 100.385 ;
        RECT 76.635 99.755 76.805 100.555 ;
        RECT 76.975 99.535 77.305 100.385 ;
        RECT 77.475 99.755 77.645 100.555 ;
        RECT 77.815 99.535 78.145 100.385 ;
        RECT 78.315 99.755 78.485 100.555 ;
        RECT 78.655 99.535 78.985 100.385 ;
        RECT 79.155 99.755 79.325 100.555 ;
        RECT 79.495 99.535 79.825 100.385 ;
        RECT 79.995 99.755 80.165 100.555 ;
        RECT 80.335 99.535 80.665 100.385 ;
        RECT 80.835 99.755 81.005 100.555 ;
        RECT 81.175 99.535 81.505 100.385 ;
        RECT 81.675 99.755 81.845 100.555 ;
        RECT 82.015 99.535 82.345 100.385 ;
        RECT 82.515 99.755 82.685 100.555 ;
        RECT 82.855 99.535 83.185 100.385 ;
        RECT 83.355 99.755 83.525 100.555 ;
        RECT 83.895 99.885 84.065 100.385 ;
        RECT 84.235 100.055 84.565 100.555 ;
        RECT 83.895 99.715 84.560 99.885 ;
        RECT 72.775 99.365 74.285 99.535 ;
        RECT 74.455 99.365 76.805 99.535 ;
        RECT 76.975 99.365 83.635 99.535 ;
        RECT 74.115 99.195 74.285 99.365 ;
        RECT 76.630 99.195 76.805 99.365 ;
        RECT 72.770 98.995 73.945 99.195 ;
        RECT 74.115 98.995 76.425 99.195 ;
        RECT 76.630 98.995 83.190 99.195 ;
        RECT 74.115 98.825 74.285 98.995 ;
        RECT 76.630 98.825 76.805 98.995 ;
        RECT 83.360 98.825 83.635 99.365 ;
        RECT 83.810 98.895 84.160 99.545 ;
        RECT 68.165 98.175 68.425 98.680 ;
        RECT 68.620 98.555 69.285 98.725 ;
        RECT 68.605 98.005 68.935 98.385 ;
        RECT 69.115 98.175 69.285 98.555 ;
        RECT 70.005 98.005 70.295 98.730 ;
        RECT 70.465 98.005 72.135 98.775 ;
        RECT 72.775 98.655 74.285 98.825 ;
        RECT 74.455 98.655 76.805 98.825 ;
        RECT 76.975 98.655 83.635 98.825 ;
        RECT 84.330 98.725 84.560 99.715 ;
        RECT 72.775 98.180 73.105 98.655 ;
        RECT 73.275 98.005 73.445 98.485 ;
        RECT 73.615 98.180 73.945 98.655 ;
        RECT 74.115 98.005 74.285 98.485 ;
        RECT 74.455 98.180 74.785 98.655 ;
        RECT 74.955 98.005 75.125 98.485 ;
        RECT 75.295 98.180 75.625 98.655 ;
        RECT 75.795 98.005 75.965 98.485 ;
        RECT 76.135 98.180 76.465 98.655 ;
        RECT 76.635 98.005 76.805 98.485 ;
        RECT 76.975 98.180 77.305 98.655 ;
        RECT 76.975 98.175 77.225 98.180 ;
        RECT 77.475 98.005 77.645 98.485 ;
        RECT 77.815 98.180 78.145 98.655 ;
        RECT 77.895 98.175 78.065 98.180 ;
        RECT 78.315 98.005 78.485 98.485 ;
        RECT 78.655 98.180 78.985 98.655 ;
        RECT 78.735 98.175 78.905 98.180 ;
        RECT 79.155 98.005 79.325 98.485 ;
        RECT 79.495 98.180 79.825 98.655 ;
        RECT 79.995 98.005 80.165 98.485 ;
        RECT 80.335 98.180 80.665 98.655 ;
        RECT 80.835 98.005 81.005 98.485 ;
        RECT 81.175 98.180 81.505 98.655 ;
        RECT 81.675 98.005 81.845 98.485 ;
        RECT 82.015 98.180 82.345 98.655 ;
        RECT 82.515 98.005 82.685 98.485 ;
        RECT 82.855 98.180 83.185 98.655 ;
        RECT 83.895 98.555 84.560 98.725 ;
        RECT 83.355 98.005 83.525 98.485 ;
        RECT 83.895 98.265 84.065 98.555 ;
        RECT 84.235 98.005 84.565 98.385 ;
        RECT 84.735 98.265 84.960 100.385 ;
        RECT 85.175 100.055 85.505 100.555 ;
        RECT 85.675 99.885 85.845 100.385 ;
        RECT 86.080 100.170 86.910 100.340 ;
        RECT 87.150 100.175 87.530 100.555 ;
        RECT 85.150 99.715 85.845 99.885 ;
        RECT 85.150 98.745 85.320 99.715 ;
        RECT 85.490 98.925 85.900 99.545 ;
        RECT 86.070 99.495 86.570 99.875 ;
        RECT 85.150 98.555 85.845 98.745 ;
        RECT 86.070 98.625 86.290 99.495 ;
        RECT 86.740 99.325 86.910 100.170 ;
        RECT 87.710 100.005 87.880 100.295 ;
        RECT 88.050 100.175 88.380 100.555 ;
        RECT 88.850 100.085 89.480 100.335 ;
        RECT 89.660 100.175 90.080 100.555 ;
        RECT 89.310 100.005 89.480 100.085 ;
        RECT 90.280 100.005 90.520 100.295 ;
        RECT 87.080 99.755 88.450 100.005 ;
        RECT 87.080 99.495 87.330 99.755 ;
        RECT 87.840 99.325 88.090 99.485 ;
        RECT 86.740 99.155 88.090 99.325 ;
        RECT 86.740 99.115 87.160 99.155 ;
        RECT 86.470 98.565 86.820 98.935 ;
        RECT 85.175 98.005 85.505 98.385 ;
        RECT 85.675 98.225 85.845 98.555 ;
        RECT 86.990 98.385 87.160 99.115 ;
        RECT 88.260 98.985 88.450 99.755 ;
        RECT 87.330 98.655 87.740 98.985 ;
        RECT 88.030 98.645 88.450 98.985 ;
        RECT 88.620 99.575 89.140 99.885 ;
        RECT 89.310 99.835 90.520 100.005 ;
        RECT 90.750 99.865 91.080 100.555 ;
        RECT 88.620 98.815 88.790 99.575 ;
        RECT 88.960 98.985 89.140 99.395 ;
        RECT 89.310 99.325 89.480 99.835 ;
        RECT 91.250 99.685 91.420 100.295 ;
        RECT 91.690 99.835 92.020 100.345 ;
        RECT 91.250 99.665 91.570 99.685 ;
        RECT 89.650 99.495 91.570 99.665 ;
        RECT 89.310 99.155 91.210 99.325 ;
        RECT 89.540 98.815 89.870 98.935 ;
        RECT 88.620 98.645 89.870 98.815 ;
        RECT 86.145 98.185 87.160 98.385 ;
        RECT 87.330 98.005 87.740 98.445 ;
        RECT 88.030 98.215 88.280 98.645 ;
        RECT 88.480 98.005 88.800 98.465 ;
        RECT 90.040 98.395 90.210 99.155 ;
        RECT 90.880 99.095 91.210 99.155 ;
        RECT 90.400 98.925 90.730 98.985 ;
        RECT 90.400 98.655 91.060 98.925 ;
        RECT 91.380 98.600 91.570 99.495 ;
        RECT 89.360 98.225 90.210 98.395 ;
        RECT 90.410 98.005 91.070 98.485 ;
        RECT 91.250 98.270 91.570 98.600 ;
        RECT 91.770 99.245 92.020 99.835 ;
        RECT 92.200 99.755 92.485 100.555 ;
        RECT 92.665 99.575 92.920 100.245 ;
        RECT 91.770 98.915 92.570 99.245 ;
        RECT 91.770 98.265 92.020 98.915 ;
        RECT 92.740 98.715 92.920 99.575 ;
        RECT 92.665 98.515 92.920 98.715 ;
        RECT 93.925 99.480 94.195 100.385 ;
        RECT 94.365 99.795 94.695 100.555 ;
        RECT 94.875 99.625 95.045 100.385 ;
        RECT 93.925 98.680 94.095 99.480 ;
        RECT 94.380 99.455 95.045 99.625 ;
        RECT 94.380 99.310 94.550 99.455 ;
        RECT 95.765 99.390 96.055 100.555 ;
        RECT 96.230 99.415 96.565 100.385 ;
        RECT 96.735 99.415 96.905 100.555 ;
        RECT 97.075 100.215 99.105 100.385 ;
        RECT 94.265 98.980 94.550 99.310 ;
        RECT 94.380 98.725 94.550 98.980 ;
        RECT 94.785 98.905 95.115 99.275 ;
        RECT 96.230 98.745 96.400 99.415 ;
        RECT 97.075 99.245 97.245 100.215 ;
        RECT 96.570 98.915 96.825 99.245 ;
        RECT 97.050 98.915 97.245 99.245 ;
        RECT 97.415 99.875 98.540 100.045 ;
        RECT 96.655 98.745 96.825 98.915 ;
        RECT 97.415 98.745 97.585 99.875 ;
        RECT 92.200 98.005 92.485 98.465 ;
        RECT 92.665 98.345 93.005 98.515 ;
        RECT 92.665 98.185 92.920 98.345 ;
        RECT 93.925 98.175 94.185 98.680 ;
        RECT 94.380 98.555 95.045 98.725 ;
        RECT 94.365 98.005 94.695 98.385 ;
        RECT 94.875 98.175 95.045 98.555 ;
        RECT 95.765 98.005 96.055 98.730 ;
        RECT 96.230 98.175 96.485 98.745 ;
        RECT 96.655 98.575 97.585 98.745 ;
        RECT 97.755 99.535 98.765 99.705 ;
        RECT 97.755 98.735 97.925 99.535 ;
        RECT 97.410 98.540 97.585 98.575 ;
        RECT 96.655 98.005 96.985 98.405 ;
        RECT 97.410 98.175 97.940 98.540 ;
        RECT 98.130 98.515 98.405 99.335 ;
        RECT 98.125 98.345 98.405 98.515 ;
        RECT 98.130 98.175 98.405 98.345 ;
        RECT 98.575 98.175 98.765 99.535 ;
        RECT 98.935 99.550 99.105 100.215 ;
        RECT 99.275 99.795 99.445 100.555 ;
        RECT 99.680 99.795 100.195 100.205 ;
        RECT 98.935 99.360 99.685 99.550 ;
        RECT 99.855 98.985 100.195 99.795 ;
        RECT 100.365 99.585 100.625 100.555 ;
        RECT 98.965 98.815 100.195 98.985 ;
        RECT 98.945 98.005 99.455 98.540 ;
        RECT 99.675 98.210 99.920 98.815 ;
        RECT 100.365 98.295 100.605 99.245 ;
        RECT 100.795 99.210 101.125 100.385 ;
        RECT 101.295 99.585 101.575 100.555 ;
        RECT 102.755 99.885 102.925 100.385 ;
        RECT 103.095 100.055 103.425 100.555 ;
        RECT 102.755 99.715 103.420 99.885 ;
        RECT 100.795 98.680 101.575 99.210 ;
        RECT 102.670 98.895 103.020 99.545 ;
        RECT 103.190 98.725 103.420 99.715 ;
        RECT 100.795 98.175 101.120 98.680 ;
        RECT 102.755 98.555 103.420 98.725 ;
        RECT 101.290 98.005 101.575 98.510 ;
        RECT 102.755 98.265 102.925 98.555 ;
        RECT 103.095 98.005 103.425 98.385 ;
        RECT 103.595 98.265 103.820 100.385 ;
        RECT 104.035 100.055 104.365 100.555 ;
        RECT 104.535 99.885 104.705 100.385 ;
        RECT 104.940 100.170 105.770 100.340 ;
        RECT 106.010 100.175 106.390 100.555 ;
        RECT 104.010 99.715 104.705 99.885 ;
        RECT 104.010 98.745 104.180 99.715 ;
        RECT 104.350 98.925 104.760 99.545 ;
        RECT 104.930 99.495 105.430 99.875 ;
        RECT 104.010 98.555 104.705 98.745 ;
        RECT 104.930 98.625 105.150 99.495 ;
        RECT 105.600 99.325 105.770 100.170 ;
        RECT 106.570 100.005 106.740 100.295 ;
        RECT 106.910 100.175 107.240 100.555 ;
        RECT 107.710 100.085 108.340 100.335 ;
        RECT 108.520 100.175 108.940 100.555 ;
        RECT 108.170 100.005 108.340 100.085 ;
        RECT 109.140 100.005 109.380 100.295 ;
        RECT 105.940 99.755 107.310 100.005 ;
        RECT 105.940 99.495 106.190 99.755 ;
        RECT 106.700 99.325 106.950 99.485 ;
        RECT 105.600 99.155 106.950 99.325 ;
        RECT 105.600 99.115 106.020 99.155 ;
        RECT 105.330 98.565 105.680 98.935 ;
        RECT 104.035 98.005 104.365 98.385 ;
        RECT 104.535 98.225 104.705 98.555 ;
        RECT 105.850 98.385 106.020 99.115 ;
        RECT 107.120 98.985 107.310 99.755 ;
        RECT 106.190 98.655 106.600 98.985 ;
        RECT 106.890 98.645 107.310 98.985 ;
        RECT 107.480 99.575 108.000 99.885 ;
        RECT 108.170 99.835 109.380 100.005 ;
        RECT 109.610 99.865 109.940 100.555 ;
        RECT 107.480 98.815 107.650 99.575 ;
        RECT 107.820 98.985 108.000 99.395 ;
        RECT 108.170 99.325 108.340 99.835 ;
        RECT 110.110 99.685 110.280 100.295 ;
        RECT 110.550 99.835 110.880 100.345 ;
        RECT 110.110 99.665 110.430 99.685 ;
        RECT 108.510 99.495 110.430 99.665 ;
        RECT 108.170 99.155 110.070 99.325 ;
        RECT 108.400 98.815 108.730 98.935 ;
        RECT 107.480 98.645 108.730 98.815 ;
        RECT 105.005 98.185 106.020 98.385 ;
        RECT 106.190 98.005 106.600 98.445 ;
        RECT 106.890 98.215 107.140 98.645 ;
        RECT 107.340 98.005 107.660 98.465 ;
        RECT 108.900 98.395 109.070 99.155 ;
        RECT 109.740 99.095 110.070 99.155 ;
        RECT 109.260 98.925 109.590 98.985 ;
        RECT 109.260 98.655 109.920 98.925 ;
        RECT 110.240 98.600 110.430 99.495 ;
        RECT 108.220 98.225 109.070 98.395 ;
        RECT 109.270 98.005 109.930 98.485 ;
        RECT 110.110 98.270 110.430 98.600 ;
        RECT 110.630 99.245 110.880 99.835 ;
        RECT 111.060 99.755 111.345 100.555 ;
        RECT 111.525 99.575 111.780 100.245 ;
        RECT 110.630 98.915 111.430 99.245 ;
        RECT 110.630 98.265 110.880 98.915 ;
        RECT 111.600 98.715 111.780 99.575 ;
        RECT 112.325 99.465 113.535 100.555 ;
        RECT 112.325 98.925 112.845 99.465 ;
        RECT 113.015 98.755 113.535 99.295 ;
        RECT 111.525 98.515 111.780 98.715 ;
        RECT 111.060 98.005 111.345 98.465 ;
        RECT 111.525 98.345 111.865 98.515 ;
        RECT 111.525 98.185 111.780 98.345 ;
        RECT 112.325 98.005 113.535 98.755 ;
        RECT 5.520 97.835 113.620 98.005 ;
        RECT 5.605 97.085 6.815 97.835 ;
        RECT 5.605 96.545 6.125 97.085 ;
        RECT 6.985 97.065 10.495 97.835 ;
        RECT 11.125 97.160 11.385 97.665 ;
        RECT 11.565 97.455 11.895 97.835 ;
        RECT 12.075 97.285 12.245 97.665 ;
        RECT 6.295 96.375 6.815 96.915 ;
        RECT 6.985 96.545 8.635 97.065 ;
        RECT 8.805 96.375 10.495 96.895 ;
        RECT 5.605 95.285 6.815 96.375 ;
        RECT 6.985 95.285 10.495 96.375 ;
        RECT 11.125 96.360 11.295 97.160 ;
        RECT 11.580 97.115 12.245 97.285 ;
        RECT 11.580 96.860 11.750 97.115 ;
        RECT 13.025 97.015 13.235 97.835 ;
        RECT 13.405 97.035 13.735 97.665 ;
        RECT 11.465 96.530 11.750 96.860 ;
        RECT 11.985 96.565 12.315 96.935 ;
        RECT 11.580 96.385 11.750 96.530 ;
        RECT 13.405 96.435 13.655 97.035 ;
        RECT 13.905 97.015 14.135 97.835 ;
        RECT 14.345 97.065 16.935 97.835 ;
        RECT 17.565 97.160 17.825 97.665 ;
        RECT 18.005 97.455 18.335 97.835 ;
        RECT 18.515 97.285 18.685 97.665 ;
        RECT 13.825 96.595 14.155 96.845 ;
        RECT 14.345 96.545 15.555 97.065 ;
        RECT 11.125 95.455 11.395 96.360 ;
        RECT 11.580 96.215 12.245 96.385 ;
        RECT 11.565 95.285 11.895 96.045 ;
        RECT 12.075 95.455 12.245 96.215 ;
        RECT 13.025 95.285 13.235 96.425 ;
        RECT 13.405 95.455 13.735 96.435 ;
        RECT 13.905 95.285 14.135 96.425 ;
        RECT 15.725 96.375 16.935 96.895 ;
        RECT 14.345 95.285 16.935 96.375 ;
        RECT 17.565 96.360 17.735 97.160 ;
        RECT 18.020 97.115 18.685 97.285 ;
        RECT 18.020 96.860 18.190 97.115 ;
        RECT 17.905 96.530 18.190 96.860 ;
        RECT 18.425 96.565 18.755 96.935 ;
        RECT 18.945 96.595 19.185 97.545 ;
        RECT 19.375 97.160 19.700 97.665 ;
        RECT 19.870 97.330 20.155 97.835 ;
        RECT 20.325 97.325 20.630 97.835 ;
        RECT 19.375 96.630 20.155 97.160 ;
        RECT 18.020 96.385 18.190 96.530 ;
        RECT 17.565 95.455 17.835 96.360 ;
        RECT 18.020 96.215 18.685 96.385 ;
        RECT 18.005 95.285 18.335 96.045 ;
        RECT 18.515 95.455 18.685 96.215 ;
        RECT 18.945 95.285 19.205 96.255 ;
        RECT 19.375 95.455 19.705 96.630 ;
        RECT 20.325 96.595 20.640 97.155 ;
        RECT 20.810 96.845 21.060 97.655 ;
        RECT 21.230 97.310 21.490 97.835 ;
        RECT 21.670 96.845 21.920 97.655 ;
        RECT 22.090 97.275 22.350 97.835 ;
        RECT 22.520 97.185 22.780 97.640 ;
        RECT 22.950 97.355 23.210 97.835 ;
        RECT 23.380 97.185 23.640 97.640 ;
        RECT 23.810 97.355 24.070 97.835 ;
        RECT 24.240 97.185 24.500 97.640 ;
        RECT 24.670 97.355 24.915 97.835 ;
        RECT 25.085 97.185 25.360 97.640 ;
        RECT 25.530 97.355 25.775 97.835 ;
        RECT 25.945 97.185 26.205 97.640 ;
        RECT 26.385 97.355 26.635 97.835 ;
        RECT 26.805 97.185 27.065 97.640 ;
        RECT 27.245 97.355 27.495 97.835 ;
        RECT 27.665 97.185 27.925 97.640 ;
        RECT 28.105 97.355 28.365 97.835 ;
        RECT 28.535 97.185 28.795 97.640 ;
        RECT 28.965 97.355 29.265 97.835 ;
        RECT 22.520 97.015 29.265 97.185 ;
        RECT 29.585 97.015 29.795 97.835 ;
        RECT 29.965 97.035 30.295 97.665 ;
        RECT 20.810 96.595 27.930 96.845 ;
        RECT 19.875 95.285 20.155 96.255 ;
        RECT 20.335 95.285 20.630 96.095 ;
        RECT 20.810 95.455 21.055 96.595 ;
        RECT 21.230 95.285 21.490 96.095 ;
        RECT 21.670 95.460 21.920 96.595 ;
        RECT 28.100 96.425 29.265 97.015 ;
        RECT 29.965 96.435 30.215 97.035 ;
        RECT 30.465 97.015 30.695 97.835 ;
        RECT 31.365 97.110 31.655 97.835 ;
        RECT 31.825 97.085 33.035 97.835 ;
        RECT 33.210 97.095 33.465 97.665 ;
        RECT 33.635 97.435 33.965 97.835 ;
        RECT 34.390 97.300 34.920 97.665 ;
        RECT 35.110 97.495 35.385 97.665 ;
        RECT 35.105 97.325 35.385 97.495 ;
        RECT 34.390 97.265 34.565 97.300 ;
        RECT 33.635 97.095 34.565 97.265 ;
        RECT 30.385 96.595 30.715 96.845 ;
        RECT 31.825 96.545 32.345 97.085 ;
        RECT 22.520 96.200 29.265 96.425 ;
        RECT 22.520 96.185 27.925 96.200 ;
        RECT 22.090 95.290 22.350 96.085 ;
        RECT 22.520 95.460 22.780 96.185 ;
        RECT 22.950 95.290 23.210 96.015 ;
        RECT 23.380 95.460 23.640 96.185 ;
        RECT 23.810 95.290 24.070 96.015 ;
        RECT 24.240 95.460 24.500 96.185 ;
        RECT 24.670 95.290 24.930 96.015 ;
        RECT 25.100 95.460 25.360 96.185 ;
        RECT 25.530 95.290 25.775 96.015 ;
        RECT 25.945 95.460 26.205 96.185 ;
        RECT 26.390 95.290 26.635 96.015 ;
        RECT 26.805 95.460 27.065 96.185 ;
        RECT 27.250 95.290 27.495 96.015 ;
        RECT 27.665 95.460 27.925 96.185 ;
        RECT 28.110 95.290 28.365 96.015 ;
        RECT 28.535 95.460 28.825 96.200 ;
        RECT 22.090 95.285 28.365 95.290 ;
        RECT 28.995 95.285 29.265 96.030 ;
        RECT 29.585 95.285 29.795 96.425 ;
        RECT 29.965 95.455 30.295 96.435 ;
        RECT 30.465 95.285 30.695 96.425 ;
        RECT 31.365 95.285 31.655 96.450 ;
        RECT 32.515 96.375 33.035 96.915 ;
        RECT 31.825 95.285 33.035 96.375 ;
        RECT 33.210 96.425 33.380 97.095 ;
        RECT 33.635 96.925 33.805 97.095 ;
        RECT 33.550 96.595 33.805 96.925 ;
        RECT 34.030 96.595 34.225 96.925 ;
        RECT 33.210 95.455 33.545 96.425 ;
        RECT 33.715 95.285 33.885 96.425 ;
        RECT 34.055 95.625 34.225 96.595 ;
        RECT 34.395 95.965 34.565 97.095 ;
        RECT 34.735 96.305 34.905 97.105 ;
        RECT 35.110 96.505 35.385 97.325 ;
        RECT 35.555 96.305 35.745 97.665 ;
        RECT 35.925 97.300 36.435 97.835 ;
        RECT 36.655 97.025 36.900 97.630 ;
        RECT 37.720 97.125 37.975 97.655 ;
        RECT 38.155 97.375 38.440 97.835 ;
        RECT 35.945 96.855 37.175 97.025 ;
        RECT 34.735 96.135 35.745 96.305 ;
        RECT 35.915 96.290 36.665 96.480 ;
        RECT 34.395 95.795 35.520 95.965 ;
        RECT 35.915 95.625 36.085 96.290 ;
        RECT 36.835 96.045 37.175 96.855 ;
        RECT 37.720 96.815 37.900 97.125 ;
        RECT 38.620 96.925 38.870 97.575 ;
        RECT 37.635 96.645 37.900 96.815 ;
        RECT 34.055 95.455 36.085 95.625 ;
        RECT 36.255 95.285 36.425 96.045 ;
        RECT 36.660 95.635 37.175 96.045 ;
        RECT 37.720 96.265 37.900 96.645 ;
        RECT 38.070 96.595 38.870 96.925 ;
        RECT 37.720 95.595 37.975 96.265 ;
        RECT 38.155 95.285 38.440 96.085 ;
        RECT 38.620 96.005 38.870 96.595 ;
        RECT 39.070 97.240 39.390 97.570 ;
        RECT 39.570 97.355 40.230 97.835 ;
        RECT 40.430 97.445 41.280 97.615 ;
        RECT 39.070 96.345 39.260 97.240 ;
        RECT 39.580 96.915 40.240 97.185 ;
        RECT 39.910 96.855 40.240 96.915 ;
        RECT 39.430 96.685 39.760 96.745 ;
        RECT 40.430 96.685 40.600 97.445 ;
        RECT 41.840 97.375 42.160 97.835 ;
        RECT 42.360 97.195 42.610 97.625 ;
        RECT 42.900 97.395 43.310 97.835 ;
        RECT 43.480 97.455 44.495 97.655 ;
        RECT 40.770 97.025 42.020 97.195 ;
        RECT 40.770 96.905 41.100 97.025 ;
        RECT 39.430 96.515 41.330 96.685 ;
        RECT 39.070 96.175 40.990 96.345 ;
        RECT 39.070 96.155 39.390 96.175 ;
        RECT 38.620 95.495 38.950 96.005 ;
        RECT 39.220 95.545 39.390 96.155 ;
        RECT 41.160 96.005 41.330 96.515 ;
        RECT 41.500 96.445 41.680 96.855 ;
        RECT 41.850 96.265 42.020 97.025 ;
        RECT 39.560 95.285 39.890 95.975 ;
        RECT 40.120 95.835 41.330 96.005 ;
        RECT 41.500 95.955 42.020 96.265 ;
        RECT 42.190 96.855 42.610 97.195 ;
        RECT 42.900 96.855 43.310 97.185 ;
        RECT 42.190 96.085 42.380 96.855 ;
        RECT 43.480 96.725 43.650 97.455 ;
        RECT 44.795 97.285 44.965 97.615 ;
        RECT 45.135 97.455 45.465 97.835 ;
        RECT 43.820 96.905 44.170 97.275 ;
        RECT 43.480 96.685 43.900 96.725 ;
        RECT 42.550 96.515 43.900 96.685 ;
        RECT 42.550 96.355 42.800 96.515 ;
        RECT 43.310 96.085 43.560 96.345 ;
        RECT 42.190 95.835 43.560 96.085 ;
        RECT 40.120 95.545 40.360 95.835 ;
        RECT 41.160 95.755 41.330 95.835 ;
        RECT 40.560 95.285 40.980 95.665 ;
        RECT 41.160 95.505 41.790 95.755 ;
        RECT 42.260 95.285 42.590 95.665 ;
        RECT 42.760 95.545 42.930 95.835 ;
        RECT 43.730 95.670 43.900 96.515 ;
        RECT 44.350 96.345 44.570 97.215 ;
        RECT 44.795 97.095 45.490 97.285 ;
        RECT 44.070 95.965 44.570 96.345 ;
        RECT 44.740 96.295 45.150 96.915 ;
        RECT 45.320 96.125 45.490 97.095 ;
        RECT 44.795 95.955 45.490 96.125 ;
        RECT 43.110 95.285 43.490 95.665 ;
        RECT 43.730 95.500 44.560 95.670 ;
        RECT 44.795 95.455 44.965 95.955 ;
        RECT 45.135 95.285 45.465 95.785 ;
        RECT 45.680 95.455 45.905 97.575 ;
        RECT 46.075 97.455 46.405 97.835 ;
        RECT 46.575 97.285 46.745 97.575 ;
        RECT 47.005 97.325 47.310 97.835 ;
        RECT 46.080 97.115 46.745 97.285 ;
        RECT 46.080 96.125 46.310 97.115 ;
        RECT 46.480 96.295 46.830 96.945 ;
        RECT 47.005 96.595 47.320 97.155 ;
        RECT 47.490 96.845 47.740 97.655 ;
        RECT 47.910 97.310 48.170 97.835 ;
        RECT 48.350 96.845 48.600 97.655 ;
        RECT 48.770 97.275 49.030 97.835 ;
        RECT 49.200 97.185 49.460 97.640 ;
        RECT 49.630 97.355 49.890 97.835 ;
        RECT 50.060 97.185 50.320 97.640 ;
        RECT 50.490 97.355 50.750 97.835 ;
        RECT 50.920 97.185 51.180 97.640 ;
        RECT 51.350 97.355 51.595 97.835 ;
        RECT 51.765 97.185 52.040 97.640 ;
        RECT 52.210 97.355 52.455 97.835 ;
        RECT 52.625 97.185 52.885 97.640 ;
        RECT 53.065 97.355 53.315 97.835 ;
        RECT 53.485 97.185 53.745 97.640 ;
        RECT 53.925 97.355 54.175 97.835 ;
        RECT 54.345 97.185 54.605 97.640 ;
        RECT 54.785 97.355 55.045 97.835 ;
        RECT 55.215 97.185 55.475 97.640 ;
        RECT 55.645 97.355 55.945 97.835 ;
        RECT 49.200 97.015 55.945 97.185 ;
        RECT 57.125 97.110 57.415 97.835 ;
        RECT 57.645 97.015 57.855 97.835 ;
        RECT 58.025 97.035 58.355 97.665 ;
        RECT 47.490 96.595 54.610 96.845 ;
        RECT 46.080 95.955 46.745 96.125 ;
        RECT 46.075 95.285 46.405 95.785 ;
        RECT 46.575 95.455 46.745 95.955 ;
        RECT 47.015 95.285 47.310 96.095 ;
        RECT 47.490 95.455 47.735 96.595 ;
        RECT 47.910 95.285 48.170 96.095 ;
        RECT 48.350 95.460 48.600 96.595 ;
        RECT 54.780 96.425 55.945 97.015 ;
        RECT 49.200 96.200 55.945 96.425 ;
        RECT 49.200 96.185 54.605 96.200 ;
        RECT 48.770 95.290 49.030 96.085 ;
        RECT 49.200 95.460 49.460 96.185 ;
        RECT 49.630 95.290 49.890 96.015 ;
        RECT 50.060 95.460 50.320 96.185 ;
        RECT 50.490 95.290 50.750 96.015 ;
        RECT 50.920 95.460 51.180 96.185 ;
        RECT 51.350 95.290 51.610 96.015 ;
        RECT 51.780 95.460 52.040 96.185 ;
        RECT 52.210 95.290 52.455 96.015 ;
        RECT 52.625 95.460 52.885 96.185 ;
        RECT 53.070 95.290 53.315 96.015 ;
        RECT 53.485 95.460 53.745 96.185 ;
        RECT 53.930 95.290 54.175 96.015 ;
        RECT 54.345 95.460 54.605 96.185 ;
        RECT 54.790 95.290 55.045 96.015 ;
        RECT 55.215 95.460 55.505 96.200 ;
        RECT 48.770 95.285 55.045 95.290 ;
        RECT 55.675 95.285 55.945 96.030 ;
        RECT 57.125 95.285 57.415 96.450 ;
        RECT 58.025 96.435 58.275 97.035 ;
        RECT 58.525 97.015 58.755 97.835 ;
        RECT 59.885 97.160 60.145 97.665 ;
        RECT 60.325 97.455 60.655 97.835 ;
        RECT 60.835 97.285 61.005 97.665 ;
        RECT 58.445 96.595 58.775 96.845 ;
        RECT 57.645 95.285 57.855 96.425 ;
        RECT 58.025 95.455 58.355 96.435 ;
        RECT 58.525 95.285 58.755 96.425 ;
        RECT 59.885 96.360 60.055 97.160 ;
        RECT 60.340 97.115 61.005 97.285 ;
        RECT 60.340 96.860 60.510 97.115 ;
        RECT 61.265 97.065 64.775 97.835 ;
        RECT 65.495 97.285 65.665 97.575 ;
        RECT 65.835 97.455 66.165 97.835 ;
        RECT 65.495 97.115 66.160 97.285 ;
        RECT 60.225 96.530 60.510 96.860 ;
        RECT 60.745 96.565 61.075 96.935 ;
        RECT 61.265 96.545 62.915 97.065 ;
        RECT 60.340 96.385 60.510 96.530 ;
        RECT 59.885 95.455 60.155 96.360 ;
        RECT 60.340 96.215 61.005 96.385 ;
        RECT 63.085 96.375 64.775 96.895 ;
        RECT 60.325 95.285 60.655 96.045 ;
        RECT 60.835 95.455 61.005 96.215 ;
        RECT 61.265 95.285 64.775 96.375 ;
        RECT 65.410 96.295 65.760 96.945 ;
        RECT 65.930 96.125 66.160 97.115 ;
        RECT 65.495 95.955 66.160 96.125 ;
        RECT 65.495 95.455 65.665 95.955 ;
        RECT 65.835 95.285 66.165 95.785 ;
        RECT 66.335 95.455 66.560 97.575 ;
        RECT 66.775 97.455 67.105 97.835 ;
        RECT 67.275 97.285 67.445 97.615 ;
        RECT 67.745 97.455 68.760 97.655 ;
        RECT 66.750 97.095 67.445 97.285 ;
        RECT 66.750 96.125 66.920 97.095 ;
        RECT 67.090 96.295 67.500 96.915 ;
        RECT 67.670 96.345 67.890 97.215 ;
        RECT 68.070 96.905 68.420 97.275 ;
        RECT 68.590 96.725 68.760 97.455 ;
        RECT 68.930 97.395 69.340 97.835 ;
        RECT 69.630 97.195 69.880 97.625 ;
        RECT 70.080 97.375 70.400 97.835 ;
        RECT 70.960 97.445 71.810 97.615 ;
        RECT 68.930 96.855 69.340 97.185 ;
        RECT 69.630 96.855 70.050 97.195 ;
        RECT 68.340 96.685 68.760 96.725 ;
        RECT 68.340 96.515 69.690 96.685 ;
        RECT 66.750 95.955 67.445 96.125 ;
        RECT 67.670 95.965 68.170 96.345 ;
        RECT 66.775 95.285 67.105 95.785 ;
        RECT 67.275 95.455 67.445 95.955 ;
        RECT 68.340 95.670 68.510 96.515 ;
        RECT 69.440 96.355 69.690 96.515 ;
        RECT 68.680 96.085 68.930 96.345 ;
        RECT 69.860 96.085 70.050 96.855 ;
        RECT 68.680 95.835 70.050 96.085 ;
        RECT 70.220 97.025 71.470 97.195 ;
        RECT 70.220 96.265 70.390 97.025 ;
        RECT 71.140 96.905 71.470 97.025 ;
        RECT 70.560 96.445 70.740 96.855 ;
        RECT 71.640 96.685 71.810 97.445 ;
        RECT 72.010 97.355 72.670 97.835 ;
        RECT 72.850 97.240 73.170 97.570 ;
        RECT 72.000 96.915 72.660 97.185 ;
        RECT 72.000 96.855 72.330 96.915 ;
        RECT 72.480 96.685 72.810 96.745 ;
        RECT 70.910 96.515 72.810 96.685 ;
        RECT 70.220 95.955 70.740 96.265 ;
        RECT 70.910 96.005 71.080 96.515 ;
        RECT 72.980 96.345 73.170 97.240 ;
        RECT 71.250 96.175 73.170 96.345 ;
        RECT 72.850 96.155 73.170 96.175 ;
        RECT 73.370 96.925 73.620 97.575 ;
        RECT 73.800 97.375 74.085 97.835 ;
        RECT 74.265 97.125 74.520 97.655 ;
        RECT 73.370 96.595 74.170 96.925 ;
        RECT 70.910 95.835 72.120 96.005 ;
        RECT 67.680 95.500 68.510 95.670 ;
        RECT 68.750 95.285 69.130 95.665 ;
        RECT 69.310 95.545 69.480 95.835 ;
        RECT 70.910 95.755 71.080 95.835 ;
        RECT 69.650 95.285 69.980 95.665 ;
        RECT 70.450 95.505 71.080 95.755 ;
        RECT 71.260 95.285 71.680 95.665 ;
        RECT 71.880 95.545 72.120 95.835 ;
        RECT 72.350 95.285 72.680 95.975 ;
        RECT 72.850 95.545 73.020 96.155 ;
        RECT 73.370 96.005 73.620 96.595 ;
        RECT 74.340 96.475 74.520 97.125 ;
        RECT 75.270 97.055 75.770 97.665 ;
        RECT 75.065 96.595 75.415 96.845 ;
        RECT 74.340 96.305 74.605 96.475 ;
        RECT 75.600 96.425 75.770 97.055 ;
        RECT 76.400 97.185 76.730 97.665 ;
        RECT 76.900 97.375 77.125 97.835 ;
        RECT 77.295 97.185 77.625 97.665 ;
        RECT 76.400 97.015 77.625 97.185 ;
        RECT 77.815 97.035 78.065 97.835 ;
        RECT 78.235 97.035 78.575 97.665 ;
        RECT 78.345 96.985 78.575 97.035 ;
        RECT 78.945 97.205 79.275 97.565 ;
        RECT 79.895 97.375 80.145 97.835 ;
        RECT 80.315 97.375 80.875 97.665 ;
        RECT 78.945 97.015 80.335 97.205 ;
        RECT 75.940 96.645 76.270 96.845 ;
        RECT 76.440 96.645 76.770 96.845 ;
        RECT 76.940 96.645 77.360 96.845 ;
        RECT 77.535 96.675 78.230 96.845 ;
        RECT 77.535 96.425 77.705 96.675 ;
        RECT 78.400 96.425 78.575 96.985 ;
        RECT 80.165 96.925 80.335 97.015 ;
        RECT 74.340 96.265 74.520 96.305 ;
        RECT 73.290 95.495 73.620 96.005 ;
        RECT 73.800 95.285 74.085 96.085 ;
        RECT 74.265 95.595 74.520 96.265 ;
        RECT 75.270 96.255 77.705 96.425 ;
        RECT 75.270 95.455 75.600 96.255 ;
        RECT 75.770 95.285 76.100 96.085 ;
        RECT 76.400 95.455 76.730 96.255 ;
        RECT 77.375 95.285 77.625 96.085 ;
        RECT 77.895 95.285 78.065 96.425 ;
        RECT 78.235 95.455 78.575 96.425 ;
        RECT 78.760 96.595 79.435 96.845 ;
        RECT 79.655 96.595 79.995 96.845 ;
        RECT 80.165 96.595 80.455 96.925 ;
        RECT 78.760 96.235 79.025 96.595 ;
        RECT 80.165 96.345 80.335 96.595 ;
        RECT 79.395 96.175 80.335 96.345 ;
        RECT 78.945 95.285 79.225 95.955 ;
        RECT 79.395 95.625 79.695 96.175 ;
        RECT 80.625 96.005 80.875 97.375 ;
        RECT 81.045 97.065 82.715 97.835 ;
        RECT 82.885 97.110 83.175 97.835 ;
        RECT 83.350 97.095 83.605 97.665 ;
        RECT 83.775 97.435 84.105 97.835 ;
        RECT 84.530 97.300 85.060 97.665 ;
        RECT 84.530 97.265 84.705 97.300 ;
        RECT 83.775 97.095 84.705 97.265 ;
        RECT 81.045 96.545 81.795 97.065 ;
        RECT 81.965 96.375 82.715 96.895 ;
        RECT 79.895 95.285 80.225 96.005 ;
        RECT 80.415 95.455 80.875 96.005 ;
        RECT 81.045 95.285 82.715 96.375 ;
        RECT 82.885 95.285 83.175 96.450 ;
        RECT 83.350 96.425 83.520 97.095 ;
        RECT 83.775 96.925 83.945 97.095 ;
        RECT 83.690 96.595 83.945 96.925 ;
        RECT 84.170 96.595 84.365 96.925 ;
        RECT 83.350 95.455 83.685 96.425 ;
        RECT 83.855 95.285 84.025 96.425 ;
        RECT 84.195 95.625 84.365 96.595 ;
        RECT 84.535 95.965 84.705 97.095 ;
        RECT 84.875 96.305 85.045 97.105 ;
        RECT 85.250 96.815 85.525 97.665 ;
        RECT 85.245 96.645 85.525 96.815 ;
        RECT 85.250 96.505 85.525 96.645 ;
        RECT 85.695 96.305 85.885 97.665 ;
        RECT 86.065 97.300 86.575 97.835 ;
        RECT 86.795 97.025 87.040 97.630 ;
        RECT 87.490 97.095 87.745 97.665 ;
        RECT 87.915 97.435 88.245 97.835 ;
        RECT 88.670 97.300 89.200 97.665 ;
        RECT 88.670 97.265 88.845 97.300 ;
        RECT 87.915 97.095 88.845 97.265 ;
        RECT 86.085 96.855 87.315 97.025 ;
        RECT 84.875 96.135 85.885 96.305 ;
        RECT 86.055 96.290 86.805 96.480 ;
        RECT 84.535 95.795 85.660 95.965 ;
        RECT 86.055 95.625 86.225 96.290 ;
        RECT 86.975 96.045 87.315 96.855 ;
        RECT 84.195 95.455 86.225 95.625 ;
        RECT 86.395 95.285 86.565 96.045 ;
        RECT 86.800 95.635 87.315 96.045 ;
        RECT 87.490 96.425 87.660 97.095 ;
        RECT 87.915 96.925 88.085 97.095 ;
        RECT 87.830 96.595 88.085 96.925 ;
        RECT 88.310 96.595 88.505 96.925 ;
        RECT 87.490 95.455 87.825 96.425 ;
        RECT 87.995 95.285 88.165 96.425 ;
        RECT 88.335 95.625 88.505 96.595 ;
        RECT 88.675 95.965 88.845 97.095 ;
        RECT 89.015 96.305 89.185 97.105 ;
        RECT 89.390 96.815 89.665 97.665 ;
        RECT 89.385 96.645 89.665 96.815 ;
        RECT 89.390 96.505 89.665 96.645 ;
        RECT 89.835 96.305 90.025 97.665 ;
        RECT 90.205 97.300 90.715 97.835 ;
        RECT 90.935 97.025 91.180 97.630 ;
        RECT 91.715 97.285 91.885 97.575 ;
        RECT 92.055 97.455 92.385 97.835 ;
        RECT 91.715 97.115 92.380 97.285 ;
        RECT 90.225 96.855 91.455 97.025 ;
        RECT 89.015 96.135 90.025 96.305 ;
        RECT 90.195 96.290 90.945 96.480 ;
        RECT 88.675 95.795 89.800 95.965 ;
        RECT 90.195 95.625 90.365 96.290 ;
        RECT 91.115 96.045 91.455 96.855 ;
        RECT 91.630 96.295 91.980 96.945 ;
        RECT 92.150 96.125 92.380 97.115 ;
        RECT 88.335 95.455 90.365 95.625 ;
        RECT 90.535 95.285 90.705 96.045 ;
        RECT 90.940 95.635 91.455 96.045 ;
        RECT 91.715 95.955 92.380 96.125 ;
        RECT 91.715 95.455 91.885 95.955 ;
        RECT 92.055 95.285 92.385 95.785 ;
        RECT 92.555 95.455 92.780 97.575 ;
        RECT 92.995 97.455 93.325 97.835 ;
        RECT 93.495 97.285 93.665 97.615 ;
        RECT 93.965 97.455 94.980 97.655 ;
        RECT 92.970 97.095 93.665 97.285 ;
        RECT 92.970 96.125 93.140 97.095 ;
        RECT 93.310 96.295 93.720 96.915 ;
        RECT 93.890 96.345 94.110 97.215 ;
        RECT 94.290 96.905 94.640 97.275 ;
        RECT 94.810 96.725 94.980 97.455 ;
        RECT 95.150 97.395 95.560 97.835 ;
        RECT 95.850 97.195 96.100 97.625 ;
        RECT 96.300 97.375 96.620 97.835 ;
        RECT 97.180 97.445 98.030 97.615 ;
        RECT 95.150 96.855 95.560 97.185 ;
        RECT 95.850 96.855 96.270 97.195 ;
        RECT 94.560 96.685 94.980 96.725 ;
        RECT 94.560 96.515 95.910 96.685 ;
        RECT 92.970 95.955 93.665 96.125 ;
        RECT 93.890 95.965 94.390 96.345 ;
        RECT 92.995 95.285 93.325 95.785 ;
        RECT 93.495 95.455 93.665 95.955 ;
        RECT 94.560 95.670 94.730 96.515 ;
        RECT 95.660 96.355 95.910 96.515 ;
        RECT 94.900 96.085 95.150 96.345 ;
        RECT 96.080 96.085 96.270 96.855 ;
        RECT 94.900 95.835 96.270 96.085 ;
        RECT 96.440 97.025 97.690 97.195 ;
        RECT 96.440 96.265 96.610 97.025 ;
        RECT 97.360 96.905 97.690 97.025 ;
        RECT 96.780 96.445 96.960 96.855 ;
        RECT 97.860 96.685 98.030 97.445 ;
        RECT 98.230 97.355 98.890 97.835 ;
        RECT 99.070 97.240 99.390 97.570 ;
        RECT 98.220 96.915 98.880 97.185 ;
        RECT 98.220 96.855 98.550 96.915 ;
        RECT 98.700 96.685 99.030 96.745 ;
        RECT 97.130 96.515 99.030 96.685 ;
        RECT 96.440 95.955 96.960 96.265 ;
        RECT 97.130 96.005 97.300 96.515 ;
        RECT 99.200 96.345 99.390 97.240 ;
        RECT 97.470 96.175 99.390 96.345 ;
        RECT 99.070 96.155 99.390 96.175 ;
        RECT 99.590 96.925 99.840 97.575 ;
        RECT 100.020 97.375 100.305 97.835 ;
        RECT 100.485 97.495 100.740 97.655 ;
        RECT 100.485 97.325 100.825 97.495 ;
        RECT 100.485 97.125 100.740 97.325 ;
        RECT 99.590 96.595 100.390 96.925 ;
        RECT 97.130 95.835 98.340 96.005 ;
        RECT 93.900 95.500 94.730 95.670 ;
        RECT 94.970 95.285 95.350 95.665 ;
        RECT 95.530 95.545 95.700 95.835 ;
        RECT 97.130 95.755 97.300 95.835 ;
        RECT 95.870 95.285 96.200 95.665 ;
        RECT 96.670 95.505 97.300 95.755 ;
        RECT 97.480 95.285 97.900 95.665 ;
        RECT 98.100 95.545 98.340 95.835 ;
        RECT 98.570 95.285 98.900 95.975 ;
        RECT 99.070 95.545 99.240 96.155 ;
        RECT 99.590 96.005 99.840 96.595 ;
        RECT 100.560 96.265 100.740 97.125 ;
        RECT 101.345 97.015 101.555 97.835 ;
        RECT 101.725 97.035 102.055 97.665 ;
        RECT 101.725 96.435 101.975 97.035 ;
        RECT 102.225 97.015 102.455 97.835 ;
        RECT 103.860 97.025 104.105 97.630 ;
        RECT 104.325 97.300 104.835 97.835 ;
        RECT 103.585 96.855 104.815 97.025 ;
        RECT 102.145 96.595 102.475 96.845 ;
        RECT 99.510 95.495 99.840 96.005 ;
        RECT 100.020 95.285 100.305 96.085 ;
        RECT 100.485 95.595 100.740 96.265 ;
        RECT 101.345 95.285 101.555 96.425 ;
        RECT 101.725 95.455 102.055 96.435 ;
        RECT 102.225 95.285 102.455 96.425 ;
        RECT 103.585 96.045 103.925 96.855 ;
        RECT 104.095 96.290 104.845 96.480 ;
        RECT 103.585 95.635 104.100 96.045 ;
        RECT 104.335 95.285 104.505 96.045 ;
        RECT 104.675 95.625 104.845 96.290 ;
        RECT 105.015 96.305 105.205 97.665 ;
        RECT 105.375 96.815 105.650 97.665 ;
        RECT 105.840 97.300 106.370 97.665 ;
        RECT 106.795 97.435 107.125 97.835 ;
        RECT 106.195 97.265 106.370 97.300 ;
        RECT 105.375 96.645 105.655 96.815 ;
        RECT 105.375 96.505 105.650 96.645 ;
        RECT 105.855 96.305 106.025 97.105 ;
        RECT 105.015 96.135 106.025 96.305 ;
        RECT 106.195 97.095 107.125 97.265 ;
        RECT 107.295 97.095 107.550 97.665 ;
        RECT 108.645 97.110 108.935 97.835 ;
        RECT 106.195 95.965 106.365 97.095 ;
        RECT 106.955 96.925 107.125 97.095 ;
        RECT 105.240 95.795 106.365 95.965 ;
        RECT 106.535 96.595 106.730 96.925 ;
        RECT 106.955 96.595 107.210 96.925 ;
        RECT 106.535 95.625 106.705 96.595 ;
        RECT 107.380 96.425 107.550 97.095 ;
        RECT 109.105 97.065 111.695 97.835 ;
        RECT 112.325 97.085 113.535 97.835 ;
        RECT 109.105 96.545 110.315 97.065 ;
        RECT 104.675 95.455 106.705 95.625 ;
        RECT 106.875 95.285 107.045 96.425 ;
        RECT 107.215 95.455 107.550 96.425 ;
        RECT 108.645 95.285 108.935 96.450 ;
        RECT 110.485 96.375 111.695 96.895 ;
        RECT 109.105 95.285 111.695 96.375 ;
        RECT 112.325 96.375 112.845 96.915 ;
        RECT 113.015 96.545 113.535 97.085 ;
        RECT 112.325 95.285 113.535 96.375 ;
        RECT 5.520 95.115 113.620 95.285 ;
        RECT 5.605 94.025 6.815 95.115 ;
        RECT 6.985 94.025 10.495 95.115 ;
        RECT 5.605 93.315 6.125 93.855 ;
        RECT 6.295 93.485 6.815 94.025 ;
        RECT 6.985 93.335 8.635 93.855 ;
        RECT 8.805 93.505 10.495 94.025 ;
        RECT 11.125 94.040 11.395 94.945 ;
        RECT 11.565 94.355 11.895 95.115 ;
        RECT 12.075 94.185 12.245 94.945 ;
        RECT 5.605 92.565 6.815 93.315 ;
        RECT 6.985 92.565 10.495 93.335 ;
        RECT 11.125 93.240 11.295 94.040 ;
        RECT 11.580 94.015 12.245 94.185 ;
        RECT 11.580 93.870 11.750 94.015 ;
        RECT 13.025 93.975 13.235 95.115 ;
        RECT 11.465 93.540 11.750 93.870 ;
        RECT 13.405 93.965 13.735 94.945 ;
        RECT 13.905 93.975 14.135 95.115 ;
        RECT 14.350 93.975 14.685 94.945 ;
        RECT 14.855 93.975 15.025 95.115 ;
        RECT 15.195 94.775 17.225 94.945 ;
        RECT 11.580 93.285 11.750 93.540 ;
        RECT 11.985 93.465 12.315 93.835 ;
        RECT 11.125 92.735 11.385 93.240 ;
        RECT 11.580 93.115 12.245 93.285 ;
        RECT 11.565 92.565 11.895 92.945 ;
        RECT 12.075 92.735 12.245 93.115 ;
        RECT 13.025 92.565 13.235 93.385 ;
        RECT 13.405 93.365 13.655 93.965 ;
        RECT 13.825 93.555 14.155 93.805 ;
        RECT 13.405 92.735 13.735 93.365 ;
        RECT 13.905 92.565 14.135 93.385 ;
        RECT 14.350 93.305 14.520 93.975 ;
        RECT 15.195 93.805 15.365 94.775 ;
        RECT 14.690 93.475 14.945 93.805 ;
        RECT 15.170 93.475 15.365 93.805 ;
        RECT 15.535 94.435 16.660 94.605 ;
        RECT 14.775 93.305 14.945 93.475 ;
        RECT 15.535 93.305 15.705 94.435 ;
        RECT 14.350 92.735 14.605 93.305 ;
        RECT 14.775 93.135 15.705 93.305 ;
        RECT 15.875 94.095 16.885 94.265 ;
        RECT 15.875 93.295 16.045 94.095 ;
        RECT 16.250 93.755 16.525 93.895 ;
        RECT 16.245 93.585 16.525 93.755 ;
        RECT 15.530 93.100 15.705 93.135 ;
        RECT 14.775 92.565 15.105 92.965 ;
        RECT 15.530 92.735 16.060 93.100 ;
        RECT 16.250 92.735 16.525 93.585 ;
        RECT 16.695 92.735 16.885 94.095 ;
        RECT 17.055 94.110 17.225 94.775 ;
        RECT 17.395 94.355 17.565 95.115 ;
        RECT 17.800 94.355 18.315 94.765 ;
        RECT 17.055 93.920 17.805 94.110 ;
        RECT 17.975 93.545 18.315 94.355 ;
        RECT 18.485 93.950 18.775 95.115 ;
        RECT 18.945 94.025 21.535 95.115 ;
        RECT 22.255 94.445 22.425 94.945 ;
        RECT 22.595 94.615 22.925 95.115 ;
        RECT 22.255 94.275 22.920 94.445 ;
        RECT 17.085 93.375 18.315 93.545 ;
        RECT 17.065 92.565 17.575 93.100 ;
        RECT 17.795 92.770 18.040 93.375 ;
        RECT 18.945 93.335 20.155 93.855 ;
        RECT 20.325 93.505 21.535 94.025 ;
        RECT 22.170 93.455 22.520 94.105 ;
        RECT 18.485 92.565 18.775 93.290 ;
        RECT 18.945 92.565 21.535 93.335 ;
        RECT 22.690 93.285 22.920 94.275 ;
        RECT 22.255 93.115 22.920 93.285 ;
        RECT 22.255 92.825 22.425 93.115 ;
        RECT 22.595 92.565 22.925 92.945 ;
        RECT 23.095 92.825 23.320 94.945 ;
        RECT 23.535 94.615 23.865 95.115 ;
        RECT 24.035 94.445 24.205 94.945 ;
        RECT 24.440 94.730 25.270 94.900 ;
        RECT 25.510 94.735 25.890 95.115 ;
        RECT 23.510 94.275 24.205 94.445 ;
        RECT 23.510 93.305 23.680 94.275 ;
        RECT 23.850 93.485 24.260 94.105 ;
        RECT 24.430 94.055 24.930 94.435 ;
        RECT 23.510 93.115 24.205 93.305 ;
        RECT 24.430 93.185 24.650 94.055 ;
        RECT 25.100 93.885 25.270 94.730 ;
        RECT 26.070 94.565 26.240 94.855 ;
        RECT 26.410 94.735 26.740 95.115 ;
        RECT 27.210 94.645 27.840 94.895 ;
        RECT 28.020 94.735 28.440 95.115 ;
        RECT 27.670 94.565 27.840 94.645 ;
        RECT 28.640 94.565 28.880 94.855 ;
        RECT 25.440 94.315 26.810 94.565 ;
        RECT 25.440 94.055 25.690 94.315 ;
        RECT 26.200 93.885 26.450 94.045 ;
        RECT 25.100 93.715 26.450 93.885 ;
        RECT 25.100 93.675 25.520 93.715 ;
        RECT 24.830 93.125 25.180 93.495 ;
        RECT 23.535 92.565 23.865 92.945 ;
        RECT 24.035 92.785 24.205 93.115 ;
        RECT 25.350 92.945 25.520 93.675 ;
        RECT 26.620 93.545 26.810 94.315 ;
        RECT 25.690 93.215 26.100 93.545 ;
        RECT 26.390 93.205 26.810 93.545 ;
        RECT 26.980 94.135 27.500 94.445 ;
        RECT 27.670 94.395 28.880 94.565 ;
        RECT 29.110 94.425 29.440 95.115 ;
        RECT 26.980 93.375 27.150 94.135 ;
        RECT 27.320 93.545 27.500 93.955 ;
        RECT 27.670 93.885 27.840 94.395 ;
        RECT 29.610 94.245 29.780 94.855 ;
        RECT 30.050 94.395 30.380 94.905 ;
        RECT 29.610 94.225 29.930 94.245 ;
        RECT 28.010 94.055 29.930 94.225 ;
        RECT 27.670 93.715 29.570 93.885 ;
        RECT 27.900 93.375 28.230 93.495 ;
        RECT 26.980 93.205 28.230 93.375 ;
        RECT 24.505 92.745 25.520 92.945 ;
        RECT 25.690 92.565 26.100 93.005 ;
        RECT 26.390 92.775 26.640 93.205 ;
        RECT 26.840 92.565 27.160 93.025 ;
        RECT 28.400 92.955 28.570 93.715 ;
        RECT 29.240 93.655 29.570 93.715 ;
        RECT 28.760 93.485 29.090 93.545 ;
        RECT 28.760 93.215 29.420 93.485 ;
        RECT 29.740 93.160 29.930 94.055 ;
        RECT 27.720 92.785 28.570 92.955 ;
        RECT 28.770 92.565 29.430 93.045 ;
        RECT 29.610 92.830 29.930 93.160 ;
        RECT 30.130 93.805 30.380 94.395 ;
        RECT 30.560 94.315 30.845 95.115 ;
        RECT 31.025 94.135 31.280 94.805 ;
        RECT 31.825 94.680 37.170 95.115 ;
        RECT 30.130 93.475 30.930 93.805 ;
        RECT 30.130 92.825 30.380 93.475 ;
        RECT 31.100 93.275 31.280 94.135 ;
        RECT 31.025 93.075 31.280 93.275 ;
        RECT 33.410 93.110 33.750 93.940 ;
        RECT 35.230 93.430 35.580 94.680 ;
        RECT 37.345 94.025 40.855 95.115 ;
        RECT 37.345 93.335 38.995 93.855 ;
        RECT 39.165 93.505 40.855 94.025 ;
        RECT 41.545 93.975 41.755 95.115 ;
        RECT 41.925 93.965 42.255 94.945 ;
        RECT 42.425 93.975 42.655 95.115 ;
        RECT 42.865 94.025 44.075 95.115 ;
        RECT 30.560 92.565 30.845 93.025 ;
        RECT 31.025 92.905 31.365 93.075 ;
        RECT 31.025 92.745 31.280 92.905 ;
        RECT 31.825 92.565 37.170 93.110 ;
        RECT 37.345 92.565 40.855 93.335 ;
        RECT 41.545 92.565 41.755 93.385 ;
        RECT 41.925 93.365 42.175 93.965 ;
        RECT 42.345 93.555 42.675 93.805 ;
        RECT 41.925 92.735 42.255 93.365 ;
        RECT 42.425 92.565 42.655 93.385 ;
        RECT 42.865 93.315 43.385 93.855 ;
        RECT 43.555 93.485 44.075 94.025 ;
        RECT 44.245 93.950 44.535 95.115 ;
        RECT 44.710 93.975 45.045 94.945 ;
        RECT 45.215 93.975 45.385 95.115 ;
        RECT 45.555 94.775 47.585 94.945 ;
        RECT 42.865 92.565 44.075 93.315 ;
        RECT 44.710 93.305 44.880 93.975 ;
        RECT 45.555 93.805 45.725 94.775 ;
        RECT 45.050 93.475 45.305 93.805 ;
        RECT 45.530 93.475 45.725 93.805 ;
        RECT 45.895 94.435 47.020 94.605 ;
        RECT 45.135 93.305 45.305 93.475 ;
        RECT 45.895 93.305 46.065 94.435 ;
        RECT 44.245 92.565 44.535 93.290 ;
        RECT 44.710 92.735 44.965 93.305 ;
        RECT 45.135 93.135 46.065 93.305 ;
        RECT 46.235 94.095 47.245 94.265 ;
        RECT 46.235 93.295 46.405 94.095 ;
        RECT 45.890 93.100 46.065 93.135 ;
        RECT 45.135 92.565 45.465 92.965 ;
        RECT 45.890 92.735 46.420 93.100 ;
        RECT 46.610 93.075 46.885 93.895 ;
        RECT 46.605 92.905 46.885 93.075 ;
        RECT 46.610 92.735 46.885 92.905 ;
        RECT 47.055 92.735 47.245 94.095 ;
        RECT 47.415 94.110 47.585 94.775 ;
        RECT 47.755 94.355 47.925 95.115 ;
        RECT 48.160 94.355 48.675 94.765 ;
        RECT 47.415 93.920 48.165 94.110 ;
        RECT 48.335 93.545 48.675 94.355 ;
        RECT 48.905 93.975 49.115 95.115 ;
        RECT 47.445 93.375 48.675 93.545 ;
        RECT 49.285 93.965 49.615 94.945 ;
        RECT 49.785 93.975 50.015 95.115 ;
        RECT 50.225 94.355 50.740 94.765 ;
        RECT 50.975 94.355 51.145 95.115 ;
        RECT 51.315 94.775 53.345 94.945 ;
        RECT 47.425 92.565 47.935 93.100 ;
        RECT 48.155 92.770 48.400 93.375 ;
        RECT 48.905 92.565 49.115 93.385 ;
        RECT 49.285 93.365 49.535 93.965 ;
        RECT 49.705 93.555 50.035 93.805 ;
        RECT 50.225 93.545 50.565 94.355 ;
        RECT 51.315 94.110 51.485 94.775 ;
        RECT 51.880 94.435 53.005 94.605 ;
        RECT 50.735 93.920 51.485 94.110 ;
        RECT 51.655 94.095 52.665 94.265 ;
        RECT 49.285 92.735 49.615 93.365 ;
        RECT 49.785 92.565 50.015 93.385 ;
        RECT 50.225 93.375 51.455 93.545 ;
        RECT 50.500 92.770 50.745 93.375 ;
        RECT 50.965 92.565 51.475 93.100 ;
        RECT 51.655 92.735 51.845 94.095 ;
        RECT 52.015 93.415 52.290 93.895 ;
        RECT 52.015 93.245 52.295 93.415 ;
        RECT 52.495 93.295 52.665 94.095 ;
        RECT 52.835 93.305 53.005 94.435 ;
        RECT 53.175 93.805 53.345 94.775 ;
        RECT 53.515 93.975 53.685 95.115 ;
        RECT 53.855 93.975 54.190 94.945 ;
        RECT 53.175 93.475 53.370 93.805 ;
        RECT 53.595 93.475 53.850 93.805 ;
        RECT 53.595 93.305 53.765 93.475 ;
        RECT 54.020 93.305 54.190 93.975 ;
        RECT 52.015 92.735 52.290 93.245 ;
        RECT 52.835 93.135 53.765 93.305 ;
        RECT 52.835 93.100 53.010 93.135 ;
        RECT 52.480 92.735 53.010 93.100 ;
        RECT 53.435 92.565 53.765 92.965 ;
        RECT 53.935 92.735 54.190 93.305 ;
        RECT 54.365 94.395 54.825 94.945 ;
        RECT 55.015 94.395 55.345 95.115 ;
        RECT 54.365 93.025 54.615 94.395 ;
        RECT 55.545 94.225 55.845 94.775 ;
        RECT 56.015 94.445 56.295 95.115 ;
        RECT 56.665 94.680 62.010 95.115 ;
        RECT 62.185 94.680 67.530 95.115 ;
        RECT 54.905 94.055 55.845 94.225 ;
        RECT 54.905 93.805 55.075 94.055 ;
        RECT 56.215 93.805 56.480 94.165 ;
        RECT 54.785 93.475 55.075 93.805 ;
        RECT 55.245 93.555 55.585 93.805 ;
        RECT 55.805 93.555 56.480 93.805 ;
        RECT 54.905 93.385 55.075 93.475 ;
        RECT 54.905 93.195 56.295 93.385 ;
        RECT 54.365 92.735 54.925 93.025 ;
        RECT 55.095 92.565 55.345 93.025 ;
        RECT 55.965 92.835 56.295 93.195 ;
        RECT 58.250 93.110 58.590 93.940 ;
        RECT 60.070 93.430 60.420 94.680 ;
        RECT 63.770 93.110 64.110 93.940 ;
        RECT 65.590 93.430 65.940 94.680 ;
        RECT 67.705 94.040 67.975 94.945 ;
        RECT 68.145 94.355 68.475 95.115 ;
        RECT 68.655 94.185 68.825 94.945 ;
        RECT 67.705 93.240 67.875 94.040 ;
        RECT 68.160 94.015 68.825 94.185 ;
        RECT 68.160 93.870 68.330 94.015 ;
        RECT 70.005 93.950 70.295 95.115 ;
        RECT 70.465 94.025 72.135 95.115 ;
        RECT 72.775 94.305 73.070 95.115 ;
        RECT 68.045 93.540 68.330 93.870 ;
        RECT 68.160 93.285 68.330 93.540 ;
        RECT 68.565 93.465 68.895 93.835 ;
        RECT 70.465 93.335 71.215 93.855 ;
        RECT 71.385 93.505 72.135 94.025 ;
        RECT 73.250 93.805 73.495 94.945 ;
        RECT 73.670 94.305 73.930 95.115 ;
        RECT 74.530 95.110 80.805 95.115 ;
        RECT 74.110 93.805 74.360 94.940 ;
        RECT 74.530 94.315 74.790 95.110 ;
        RECT 74.960 94.215 75.220 94.940 ;
        RECT 75.390 94.385 75.650 95.110 ;
        RECT 75.820 94.215 76.080 94.940 ;
        RECT 76.250 94.385 76.510 95.110 ;
        RECT 76.680 94.215 76.940 94.940 ;
        RECT 77.110 94.385 77.370 95.110 ;
        RECT 77.540 94.215 77.800 94.940 ;
        RECT 77.970 94.385 78.215 95.110 ;
        RECT 78.385 94.215 78.645 94.940 ;
        RECT 78.830 94.385 79.075 95.110 ;
        RECT 79.245 94.215 79.505 94.940 ;
        RECT 79.690 94.385 79.935 95.110 ;
        RECT 80.105 94.215 80.365 94.940 ;
        RECT 80.550 94.385 80.805 95.110 ;
        RECT 74.960 94.200 80.365 94.215 ;
        RECT 80.975 94.200 81.265 94.940 ;
        RECT 81.435 94.370 81.705 95.115 ;
        RECT 81.965 94.395 82.425 94.945 ;
        RECT 82.615 94.395 82.945 95.115 ;
        RECT 74.960 93.975 81.705 94.200 ;
        RECT 56.665 92.565 62.010 93.110 ;
        RECT 62.185 92.565 67.530 93.110 ;
        RECT 67.705 92.735 67.965 93.240 ;
        RECT 68.160 93.115 68.825 93.285 ;
        RECT 68.145 92.565 68.475 92.945 ;
        RECT 68.655 92.735 68.825 93.115 ;
        RECT 70.005 92.565 70.295 93.290 ;
        RECT 70.465 92.565 72.135 93.335 ;
        RECT 72.765 93.245 73.080 93.805 ;
        RECT 73.250 93.555 80.370 93.805 ;
        RECT 72.765 92.565 73.070 93.075 ;
        RECT 73.250 92.745 73.500 93.555 ;
        RECT 73.670 92.565 73.930 93.090 ;
        RECT 74.110 92.745 74.360 93.555 ;
        RECT 80.540 93.385 81.705 93.975 ;
        RECT 74.960 93.215 81.705 93.385 ;
        RECT 74.530 92.565 74.790 93.125 ;
        RECT 74.960 92.760 75.220 93.215 ;
        RECT 75.390 92.565 75.650 93.045 ;
        RECT 75.820 92.760 76.080 93.215 ;
        RECT 76.250 92.565 76.510 93.045 ;
        RECT 76.680 92.760 76.940 93.215 ;
        RECT 77.110 92.565 77.355 93.045 ;
        RECT 77.525 92.760 77.800 93.215 ;
        RECT 77.970 92.565 78.215 93.045 ;
        RECT 78.385 92.760 78.645 93.215 ;
        RECT 78.825 92.565 79.075 93.045 ;
        RECT 79.245 92.760 79.505 93.215 ;
        RECT 79.685 92.565 79.935 93.045 ;
        RECT 80.105 92.760 80.365 93.215 ;
        RECT 80.545 92.565 80.805 93.045 ;
        RECT 80.975 92.760 81.235 93.215 ;
        RECT 81.405 92.565 81.705 93.045 ;
        RECT 81.965 93.025 82.215 94.395 ;
        RECT 83.145 94.225 83.445 94.775 ;
        RECT 83.615 94.445 83.895 95.115 ;
        RECT 82.505 94.055 83.445 94.225 ;
        RECT 84.265 94.395 84.725 94.945 ;
        RECT 84.915 94.395 85.245 95.115 ;
        RECT 82.505 93.805 82.675 94.055 ;
        RECT 83.815 93.805 84.080 94.165 ;
        RECT 82.385 93.475 82.675 93.805 ;
        RECT 82.845 93.555 83.185 93.805 ;
        RECT 83.405 93.555 84.080 93.805 ;
        RECT 82.505 93.385 82.675 93.475 ;
        RECT 82.505 93.195 83.895 93.385 ;
        RECT 81.965 92.735 82.525 93.025 ;
        RECT 82.695 92.565 82.945 93.025 ;
        RECT 83.565 92.835 83.895 93.195 ;
        RECT 84.265 93.025 84.515 94.395 ;
        RECT 85.445 94.225 85.745 94.775 ;
        RECT 85.915 94.445 86.195 95.115 ;
        RECT 84.805 94.055 85.745 94.225 ;
        RECT 86.565 94.395 87.025 94.945 ;
        RECT 87.215 94.395 87.545 95.115 ;
        RECT 84.805 93.805 84.975 94.055 ;
        RECT 86.115 93.805 86.380 94.165 ;
        RECT 84.685 93.475 84.975 93.805 ;
        RECT 85.145 93.555 85.485 93.805 ;
        RECT 85.705 93.555 86.380 93.805 ;
        RECT 84.805 93.385 84.975 93.475 ;
        RECT 84.805 93.195 86.195 93.385 ;
        RECT 84.265 92.735 84.825 93.025 ;
        RECT 84.995 92.565 85.245 93.025 ;
        RECT 85.865 92.835 86.195 93.195 ;
        RECT 86.565 93.025 86.815 94.395 ;
        RECT 87.745 94.225 88.045 94.775 ;
        RECT 88.215 94.445 88.495 95.115 ;
        RECT 87.105 94.055 88.045 94.225 ;
        RECT 87.105 93.805 87.275 94.055 ;
        RECT 88.415 93.805 88.680 94.165 ;
        RECT 88.865 94.025 90.075 95.115 ;
        RECT 86.985 93.475 87.275 93.805 ;
        RECT 87.445 93.555 87.785 93.805 ;
        RECT 88.005 93.555 88.680 93.805 ;
        RECT 87.105 93.385 87.275 93.475 ;
        RECT 87.105 93.195 88.495 93.385 ;
        RECT 86.565 92.735 87.125 93.025 ;
        RECT 87.295 92.565 87.545 93.025 ;
        RECT 88.165 92.835 88.495 93.195 ;
        RECT 88.865 93.315 89.385 93.855 ;
        RECT 89.555 93.485 90.075 94.025 ;
        RECT 90.245 94.040 90.515 94.945 ;
        RECT 90.685 94.355 91.015 95.115 ;
        RECT 91.195 94.185 91.365 94.945 ;
        RECT 88.865 92.565 90.075 93.315 ;
        RECT 90.245 93.240 90.415 94.040 ;
        RECT 90.700 94.015 91.365 94.185 ;
        RECT 91.625 94.025 95.135 95.115 ;
        RECT 90.700 93.870 90.870 94.015 ;
        RECT 90.585 93.540 90.870 93.870 ;
        RECT 90.700 93.285 90.870 93.540 ;
        RECT 91.105 93.465 91.435 93.835 ;
        RECT 91.625 93.335 93.275 93.855 ;
        RECT 93.445 93.505 95.135 94.025 ;
        RECT 95.765 93.950 96.055 95.115 ;
        RECT 96.225 94.025 98.815 95.115 ;
        RECT 96.225 93.335 97.435 93.855 ;
        RECT 97.605 93.505 98.815 94.025 ;
        RECT 99.535 94.185 99.705 94.945 ;
        RECT 99.885 94.355 100.215 95.115 ;
        RECT 99.535 94.015 100.200 94.185 ;
        RECT 100.385 94.040 100.655 94.945 ;
        RECT 100.915 94.445 101.085 94.945 ;
        RECT 101.255 94.615 101.585 95.115 ;
        RECT 100.915 94.275 101.580 94.445 ;
        RECT 100.030 93.870 100.200 94.015 ;
        RECT 99.465 93.465 99.795 93.835 ;
        RECT 100.030 93.540 100.315 93.870 ;
        RECT 90.245 92.735 90.505 93.240 ;
        RECT 90.700 93.115 91.365 93.285 ;
        RECT 90.685 92.565 91.015 92.945 ;
        RECT 91.195 92.735 91.365 93.115 ;
        RECT 91.625 92.565 95.135 93.335 ;
        RECT 95.765 92.565 96.055 93.290 ;
        RECT 96.225 92.565 98.815 93.335 ;
        RECT 100.030 93.285 100.200 93.540 ;
        RECT 99.535 93.115 100.200 93.285 ;
        RECT 100.485 93.240 100.655 94.040 ;
        RECT 100.830 93.455 101.180 94.105 ;
        RECT 101.350 93.285 101.580 94.275 ;
        RECT 99.535 92.735 99.705 93.115 ;
        RECT 99.885 92.565 100.215 92.945 ;
        RECT 100.395 92.735 100.655 93.240 ;
        RECT 100.915 93.115 101.580 93.285 ;
        RECT 100.915 92.825 101.085 93.115 ;
        RECT 101.255 92.565 101.585 92.945 ;
        RECT 101.755 92.825 101.980 94.945 ;
        RECT 102.195 94.615 102.525 95.115 ;
        RECT 102.695 94.445 102.865 94.945 ;
        RECT 103.100 94.730 103.930 94.900 ;
        RECT 104.170 94.735 104.550 95.115 ;
        RECT 102.170 94.275 102.865 94.445 ;
        RECT 102.170 93.305 102.340 94.275 ;
        RECT 102.510 93.485 102.920 94.105 ;
        RECT 103.090 94.055 103.590 94.435 ;
        RECT 102.170 93.115 102.865 93.305 ;
        RECT 103.090 93.185 103.310 94.055 ;
        RECT 103.760 93.885 103.930 94.730 ;
        RECT 104.730 94.565 104.900 94.855 ;
        RECT 105.070 94.735 105.400 95.115 ;
        RECT 105.870 94.645 106.500 94.895 ;
        RECT 106.680 94.735 107.100 95.115 ;
        RECT 106.330 94.565 106.500 94.645 ;
        RECT 107.300 94.565 107.540 94.855 ;
        RECT 104.100 94.315 105.470 94.565 ;
        RECT 104.100 94.055 104.350 94.315 ;
        RECT 104.860 93.885 105.110 94.045 ;
        RECT 103.760 93.715 105.110 93.885 ;
        RECT 103.760 93.675 104.180 93.715 ;
        RECT 103.490 93.125 103.840 93.495 ;
        RECT 102.195 92.565 102.525 92.945 ;
        RECT 102.695 92.785 102.865 93.115 ;
        RECT 104.010 92.945 104.180 93.675 ;
        RECT 105.280 93.545 105.470 94.315 ;
        RECT 104.350 93.215 104.760 93.545 ;
        RECT 105.050 93.205 105.470 93.545 ;
        RECT 105.640 94.135 106.160 94.445 ;
        RECT 106.330 94.395 107.540 94.565 ;
        RECT 107.770 94.425 108.100 95.115 ;
        RECT 105.640 93.375 105.810 94.135 ;
        RECT 105.980 93.545 106.160 93.955 ;
        RECT 106.330 93.885 106.500 94.395 ;
        RECT 108.270 94.245 108.440 94.855 ;
        RECT 108.710 94.395 109.040 94.905 ;
        RECT 108.270 94.225 108.590 94.245 ;
        RECT 106.670 94.055 108.590 94.225 ;
        RECT 106.330 93.715 108.230 93.885 ;
        RECT 106.560 93.375 106.890 93.495 ;
        RECT 105.640 93.205 106.890 93.375 ;
        RECT 103.165 92.745 104.180 92.945 ;
        RECT 104.350 92.565 104.760 93.005 ;
        RECT 105.050 92.775 105.300 93.205 ;
        RECT 105.500 92.565 105.820 93.025 ;
        RECT 107.060 92.955 107.230 93.715 ;
        RECT 107.900 93.655 108.230 93.715 ;
        RECT 107.420 93.485 107.750 93.545 ;
        RECT 107.420 93.215 108.080 93.485 ;
        RECT 108.400 93.160 108.590 94.055 ;
        RECT 106.380 92.785 107.230 92.955 ;
        RECT 107.430 92.565 108.090 93.045 ;
        RECT 108.270 92.830 108.590 93.160 ;
        RECT 108.790 93.805 109.040 94.395 ;
        RECT 109.220 94.315 109.505 95.115 ;
        RECT 109.685 94.135 109.940 94.805 ;
        RECT 109.760 94.095 109.940 94.135 ;
        RECT 109.760 93.925 110.025 94.095 ;
        RECT 110.525 93.975 110.755 95.115 ;
        RECT 110.925 93.965 111.255 94.945 ;
        RECT 111.425 93.975 111.635 95.115 ;
        RECT 112.325 94.025 113.535 95.115 ;
        RECT 108.790 93.475 109.590 93.805 ;
        RECT 108.790 92.825 109.040 93.475 ;
        RECT 109.760 93.275 109.940 93.925 ;
        RECT 110.505 93.555 110.835 93.805 ;
        RECT 109.220 92.565 109.505 93.025 ;
        RECT 109.685 92.745 109.940 93.275 ;
        RECT 110.525 92.565 110.755 93.385 ;
        RECT 111.005 93.365 111.255 93.965 ;
        RECT 112.325 93.485 112.845 94.025 ;
        RECT 110.925 92.735 111.255 93.365 ;
        RECT 111.425 92.565 111.635 93.385 ;
        RECT 113.015 93.315 113.535 93.855 ;
        RECT 112.325 92.565 113.535 93.315 ;
        RECT 5.520 92.395 113.620 92.565 ;
        RECT 5.605 91.645 6.815 92.395 ;
        RECT 7.995 91.845 8.165 92.135 ;
        RECT 8.335 92.015 8.665 92.395 ;
        RECT 7.995 91.675 8.660 91.845 ;
        RECT 5.605 91.105 6.125 91.645 ;
        RECT 6.295 90.935 6.815 91.475 ;
        RECT 5.605 89.845 6.815 90.935 ;
        RECT 7.910 90.855 8.260 91.505 ;
        RECT 8.430 90.685 8.660 91.675 ;
        RECT 7.995 90.515 8.660 90.685 ;
        RECT 7.995 90.015 8.165 90.515 ;
        RECT 8.335 89.845 8.665 90.345 ;
        RECT 8.835 90.015 9.060 92.135 ;
        RECT 9.275 92.015 9.605 92.395 ;
        RECT 9.775 91.845 9.945 92.175 ;
        RECT 10.245 92.015 11.260 92.215 ;
        RECT 9.250 91.655 9.945 91.845 ;
        RECT 9.250 90.685 9.420 91.655 ;
        RECT 9.590 90.855 10.000 91.475 ;
        RECT 10.170 90.905 10.390 91.775 ;
        RECT 10.570 91.465 10.920 91.835 ;
        RECT 11.090 91.285 11.260 92.015 ;
        RECT 11.430 91.955 11.840 92.395 ;
        RECT 12.130 91.755 12.380 92.185 ;
        RECT 12.580 91.935 12.900 92.395 ;
        RECT 13.460 92.005 14.310 92.175 ;
        RECT 11.430 91.415 11.840 91.745 ;
        RECT 12.130 91.415 12.550 91.755 ;
        RECT 10.840 91.245 11.260 91.285 ;
        RECT 10.840 91.075 12.190 91.245 ;
        RECT 9.250 90.515 9.945 90.685 ;
        RECT 10.170 90.525 10.670 90.905 ;
        RECT 9.275 89.845 9.605 90.345 ;
        RECT 9.775 90.015 9.945 90.515 ;
        RECT 10.840 90.230 11.010 91.075 ;
        RECT 11.940 90.915 12.190 91.075 ;
        RECT 11.180 90.645 11.430 90.905 ;
        RECT 12.360 90.645 12.550 91.415 ;
        RECT 11.180 90.395 12.550 90.645 ;
        RECT 12.720 91.585 13.970 91.755 ;
        RECT 12.720 90.825 12.890 91.585 ;
        RECT 13.640 91.465 13.970 91.585 ;
        RECT 13.060 91.005 13.240 91.415 ;
        RECT 14.140 91.245 14.310 92.005 ;
        RECT 14.510 91.915 15.170 92.395 ;
        RECT 15.350 91.800 15.670 92.130 ;
        RECT 14.500 91.475 15.160 91.745 ;
        RECT 14.500 91.415 14.830 91.475 ;
        RECT 14.980 91.245 15.310 91.305 ;
        RECT 13.410 91.075 15.310 91.245 ;
        RECT 12.720 90.515 13.240 90.825 ;
        RECT 13.410 90.565 13.580 91.075 ;
        RECT 15.480 90.905 15.670 91.800 ;
        RECT 13.750 90.735 15.670 90.905 ;
        RECT 15.350 90.715 15.670 90.735 ;
        RECT 15.870 91.485 16.120 92.135 ;
        RECT 16.300 91.935 16.585 92.395 ;
        RECT 16.765 91.685 17.020 92.215 ;
        RECT 15.870 91.155 16.670 91.485 ;
        RECT 13.410 90.395 14.620 90.565 ;
        RECT 10.180 90.060 11.010 90.230 ;
        RECT 11.250 89.845 11.630 90.225 ;
        RECT 11.810 90.105 11.980 90.395 ;
        RECT 13.410 90.315 13.580 90.395 ;
        RECT 12.150 89.845 12.480 90.225 ;
        RECT 12.950 90.065 13.580 90.315 ;
        RECT 13.760 89.845 14.180 90.225 ;
        RECT 14.380 90.105 14.620 90.395 ;
        RECT 14.850 89.845 15.180 90.535 ;
        RECT 15.350 90.105 15.520 90.715 ;
        RECT 15.870 90.565 16.120 91.155 ;
        RECT 16.840 90.825 17.020 91.685 ;
        RECT 16.765 90.695 17.020 90.825 ;
        RECT 17.570 91.655 17.825 92.225 ;
        RECT 17.995 91.995 18.325 92.395 ;
        RECT 18.750 91.860 19.280 92.225 ;
        RECT 18.750 91.825 18.925 91.860 ;
        RECT 17.995 91.655 18.925 91.825 ;
        RECT 17.570 90.985 17.740 91.655 ;
        RECT 17.995 91.485 18.165 91.655 ;
        RECT 17.910 91.155 18.165 91.485 ;
        RECT 18.390 91.155 18.585 91.485 ;
        RECT 15.790 90.055 16.120 90.565 ;
        RECT 16.300 89.845 16.585 90.645 ;
        RECT 16.765 90.525 17.105 90.695 ;
        RECT 16.765 90.155 17.020 90.525 ;
        RECT 17.570 90.015 17.905 90.985 ;
        RECT 18.075 89.845 18.245 90.985 ;
        RECT 18.415 90.185 18.585 91.155 ;
        RECT 18.755 90.525 18.925 91.655 ;
        RECT 19.095 90.865 19.265 91.665 ;
        RECT 19.470 91.375 19.745 92.225 ;
        RECT 19.465 91.205 19.745 91.375 ;
        RECT 19.470 91.065 19.745 91.205 ;
        RECT 19.915 90.865 20.105 92.225 ;
        RECT 20.285 91.860 20.795 92.395 ;
        RECT 21.015 91.585 21.260 92.190 ;
        RECT 21.705 91.625 24.295 92.395 ;
        RECT 24.665 91.765 24.995 92.125 ;
        RECT 25.615 91.935 25.865 92.395 ;
        RECT 26.035 91.935 26.595 92.225 ;
        RECT 20.305 91.415 21.535 91.585 ;
        RECT 19.095 90.695 20.105 90.865 ;
        RECT 20.275 90.850 21.025 91.040 ;
        RECT 18.755 90.355 19.880 90.525 ;
        RECT 20.275 90.185 20.445 90.850 ;
        RECT 21.195 90.605 21.535 91.415 ;
        RECT 21.705 91.105 22.915 91.625 ;
        RECT 24.665 91.575 26.055 91.765 ;
        RECT 25.885 91.485 26.055 91.575 ;
        RECT 23.085 90.935 24.295 91.455 ;
        RECT 18.415 90.015 20.445 90.185 ;
        RECT 20.615 89.845 20.785 90.605 ;
        RECT 21.020 90.195 21.535 90.605 ;
        RECT 21.705 89.845 24.295 90.935 ;
        RECT 24.480 91.155 25.155 91.405 ;
        RECT 25.375 91.155 25.715 91.405 ;
        RECT 25.885 91.155 26.175 91.485 ;
        RECT 24.480 90.795 24.745 91.155 ;
        RECT 25.885 90.905 26.055 91.155 ;
        RECT 25.115 90.735 26.055 90.905 ;
        RECT 24.665 89.845 24.945 90.515 ;
        RECT 25.115 90.185 25.415 90.735 ;
        RECT 26.345 90.565 26.595 91.935 ;
        RECT 25.615 89.845 25.945 90.565 ;
        RECT 26.135 90.015 26.595 90.565 ;
        RECT 27.230 91.655 27.485 92.225 ;
        RECT 27.655 91.995 27.985 92.395 ;
        RECT 28.410 91.860 28.940 92.225 ;
        RECT 29.130 92.055 29.405 92.225 ;
        RECT 29.125 91.885 29.405 92.055 ;
        RECT 28.410 91.825 28.585 91.860 ;
        RECT 27.655 91.655 28.585 91.825 ;
        RECT 27.230 90.985 27.400 91.655 ;
        RECT 27.655 91.485 27.825 91.655 ;
        RECT 27.570 91.155 27.825 91.485 ;
        RECT 28.050 91.155 28.245 91.485 ;
        RECT 27.230 90.015 27.565 90.985 ;
        RECT 27.735 89.845 27.905 90.985 ;
        RECT 28.075 90.185 28.245 91.155 ;
        RECT 28.415 90.525 28.585 91.655 ;
        RECT 28.755 90.865 28.925 91.665 ;
        RECT 29.130 91.065 29.405 91.885 ;
        RECT 29.575 90.865 29.765 92.225 ;
        RECT 29.945 91.860 30.455 92.395 ;
        RECT 30.675 91.585 30.920 92.190 ;
        RECT 31.365 91.670 31.655 92.395 ;
        RECT 31.825 91.935 32.385 92.225 ;
        RECT 32.555 91.935 32.805 92.395 ;
        RECT 29.965 91.415 31.195 91.585 ;
        RECT 28.755 90.695 29.765 90.865 ;
        RECT 29.935 90.850 30.685 91.040 ;
        RECT 28.415 90.355 29.540 90.525 ;
        RECT 29.935 90.185 30.105 90.850 ;
        RECT 30.855 90.605 31.195 91.415 ;
        RECT 28.075 90.015 30.105 90.185 ;
        RECT 30.275 89.845 30.445 90.605 ;
        RECT 30.680 90.195 31.195 90.605 ;
        RECT 31.365 89.845 31.655 91.010 ;
        RECT 31.825 90.565 32.075 91.935 ;
        RECT 33.425 91.765 33.755 92.125 ;
        RECT 34.125 91.850 39.470 92.395 ;
        RECT 39.645 91.850 44.990 92.395 ;
        RECT 32.365 91.575 33.755 91.765 ;
        RECT 32.365 91.485 32.535 91.575 ;
        RECT 32.245 91.155 32.535 91.485 ;
        RECT 32.705 91.155 33.045 91.405 ;
        RECT 33.265 91.155 33.940 91.405 ;
        RECT 32.365 90.905 32.535 91.155 ;
        RECT 32.365 90.735 33.305 90.905 ;
        RECT 33.675 90.795 33.940 91.155 ;
        RECT 35.710 91.020 36.050 91.850 ;
        RECT 31.825 90.015 32.285 90.565 ;
        RECT 32.475 89.845 32.805 90.565 ;
        RECT 33.005 90.185 33.305 90.735 ;
        RECT 33.475 89.845 33.755 90.515 ;
        RECT 37.530 90.280 37.880 91.530 ;
        RECT 41.230 91.020 41.570 91.850 ;
        RECT 45.165 91.625 47.755 92.395 ;
        RECT 48.585 91.765 48.915 92.125 ;
        RECT 49.535 91.935 49.785 92.395 ;
        RECT 49.955 91.935 50.515 92.225 ;
        RECT 43.050 90.280 43.400 91.530 ;
        RECT 45.165 91.105 46.375 91.625 ;
        RECT 48.585 91.575 49.975 91.765 ;
        RECT 49.805 91.485 49.975 91.575 ;
        RECT 46.545 90.935 47.755 91.455 ;
        RECT 34.125 89.845 39.470 90.280 ;
        RECT 39.645 89.845 44.990 90.280 ;
        RECT 45.165 89.845 47.755 90.935 ;
        RECT 48.400 91.155 49.075 91.405 ;
        RECT 49.295 91.155 49.635 91.405 ;
        RECT 49.805 91.155 50.095 91.485 ;
        RECT 48.400 90.795 48.665 91.155 ;
        RECT 49.805 90.905 49.975 91.155 ;
        RECT 49.035 90.735 49.975 90.905 ;
        RECT 48.585 89.845 48.865 90.515 ;
        RECT 49.035 90.185 49.335 90.735 ;
        RECT 50.265 90.565 50.515 91.935 ;
        RECT 50.885 91.765 51.215 92.125 ;
        RECT 51.835 91.935 52.085 92.395 ;
        RECT 52.255 91.935 52.815 92.225 ;
        RECT 50.885 91.575 52.275 91.765 ;
        RECT 52.105 91.485 52.275 91.575 ;
        RECT 50.700 91.155 51.375 91.405 ;
        RECT 51.595 91.155 51.935 91.405 ;
        RECT 52.105 91.155 52.395 91.485 ;
        RECT 50.700 90.795 50.965 91.155 ;
        RECT 52.105 90.905 52.275 91.155 ;
        RECT 49.535 89.845 49.865 90.565 ;
        RECT 50.055 90.015 50.515 90.565 ;
        RECT 51.335 90.735 52.275 90.905 ;
        RECT 50.885 89.845 51.165 90.515 ;
        RECT 51.335 90.185 51.635 90.735 ;
        RECT 52.565 90.565 52.815 91.935 ;
        RECT 53.185 91.765 53.515 92.125 ;
        RECT 54.135 91.935 54.385 92.395 ;
        RECT 54.555 91.935 55.115 92.225 ;
        RECT 53.185 91.575 54.575 91.765 ;
        RECT 54.405 91.485 54.575 91.575 ;
        RECT 53.000 91.155 53.675 91.405 ;
        RECT 53.895 91.155 54.235 91.405 ;
        RECT 54.405 91.155 54.695 91.485 ;
        RECT 53.000 90.795 53.265 91.155 ;
        RECT 54.405 90.905 54.575 91.155 ;
        RECT 51.835 89.845 52.165 90.565 ;
        RECT 52.355 90.015 52.815 90.565 ;
        RECT 53.635 90.735 54.575 90.905 ;
        RECT 53.185 89.845 53.465 90.515 ;
        RECT 53.635 90.185 53.935 90.735 ;
        RECT 54.865 90.565 55.115 91.935 ;
        RECT 55.285 91.625 56.955 92.395 ;
        RECT 57.125 91.670 57.415 92.395 ;
        RECT 57.645 91.915 57.925 92.395 ;
        RECT 58.095 91.745 58.355 92.135 ;
        RECT 58.530 91.915 58.785 92.395 ;
        RECT 58.955 91.745 59.250 92.135 ;
        RECT 59.430 91.915 59.705 92.395 ;
        RECT 59.875 91.895 60.175 92.225 ;
        RECT 55.285 91.105 56.035 91.625 ;
        RECT 57.600 91.575 59.250 91.745 ;
        RECT 56.205 90.935 56.955 91.455 ;
        RECT 57.600 91.065 58.005 91.575 ;
        RECT 58.175 91.235 59.315 91.405 ;
        RECT 54.135 89.845 54.465 90.565 ;
        RECT 54.655 90.015 55.115 90.565 ;
        RECT 55.285 89.845 56.955 90.935 ;
        RECT 57.125 89.845 57.415 91.010 ;
        RECT 57.600 90.895 58.355 91.065 ;
        RECT 57.640 89.845 57.925 90.715 ;
        RECT 58.095 90.645 58.355 90.895 ;
        RECT 59.145 90.985 59.315 91.235 ;
        RECT 59.485 91.155 59.835 91.725 ;
        RECT 60.005 90.985 60.175 91.895 ;
        RECT 59.145 90.815 60.175 90.985 ;
        RECT 58.095 90.475 59.215 90.645 ;
        RECT 58.095 90.015 58.355 90.475 ;
        RECT 58.530 89.845 58.785 90.305 ;
        RECT 58.955 90.015 59.215 90.475 ;
        RECT 59.385 89.845 59.695 90.645 ;
        RECT 59.865 90.015 60.175 90.815 ;
        RECT 60.345 91.935 60.905 92.225 ;
        RECT 61.075 91.935 61.325 92.395 ;
        RECT 60.345 90.565 60.595 91.935 ;
        RECT 61.945 91.765 62.275 92.125 ;
        RECT 60.885 91.575 62.275 91.765 ;
        RECT 62.705 91.575 62.915 92.395 ;
        RECT 63.085 91.595 63.415 92.225 ;
        RECT 60.885 91.485 61.055 91.575 ;
        RECT 60.765 91.155 61.055 91.485 ;
        RECT 61.225 91.155 61.565 91.405 ;
        RECT 61.785 91.155 62.460 91.405 ;
        RECT 60.885 90.905 61.055 91.155 ;
        RECT 60.885 90.735 61.825 90.905 ;
        RECT 62.195 90.795 62.460 91.155 ;
        RECT 63.085 90.995 63.335 91.595 ;
        RECT 63.585 91.575 63.815 92.395 ;
        RECT 64.025 91.625 67.535 92.395 ;
        RECT 67.705 91.645 68.915 92.395 ;
        RECT 63.505 91.155 63.835 91.405 ;
        RECT 64.025 91.105 65.675 91.625 ;
        RECT 60.345 90.015 60.805 90.565 ;
        RECT 60.995 89.845 61.325 90.565 ;
        RECT 61.525 90.185 61.825 90.735 ;
        RECT 61.995 89.845 62.275 90.515 ;
        RECT 62.705 89.845 62.915 90.985 ;
        RECT 63.085 90.015 63.415 90.995 ;
        RECT 63.585 89.845 63.815 90.985 ;
        RECT 65.845 90.935 67.535 91.455 ;
        RECT 67.705 91.105 68.225 91.645 ;
        RECT 69.125 91.575 69.355 92.395 ;
        RECT 69.525 91.595 69.855 92.225 ;
        RECT 68.395 90.935 68.915 91.475 ;
        RECT 69.105 91.155 69.435 91.405 ;
        RECT 69.605 90.995 69.855 91.595 ;
        RECT 70.025 91.575 70.235 92.395 ;
        RECT 70.470 91.655 70.725 92.225 ;
        RECT 70.895 91.995 71.225 92.395 ;
        RECT 71.650 91.860 72.180 92.225 ;
        RECT 71.650 91.825 71.825 91.860 ;
        RECT 70.895 91.655 71.825 91.825 ;
        RECT 64.025 89.845 67.535 90.935 ;
        RECT 67.705 89.845 68.915 90.935 ;
        RECT 69.125 89.845 69.355 90.985 ;
        RECT 69.525 90.015 69.855 90.995 ;
        RECT 70.470 90.985 70.640 91.655 ;
        RECT 70.895 91.485 71.065 91.655 ;
        RECT 70.810 91.155 71.065 91.485 ;
        RECT 71.290 91.155 71.485 91.485 ;
        RECT 70.025 89.845 70.235 90.985 ;
        RECT 70.470 90.015 70.805 90.985 ;
        RECT 70.975 89.845 71.145 90.985 ;
        RECT 71.315 90.185 71.485 91.155 ;
        RECT 71.655 90.525 71.825 91.655 ;
        RECT 71.995 90.865 72.165 91.665 ;
        RECT 72.370 91.375 72.645 92.225 ;
        RECT 72.365 91.205 72.645 91.375 ;
        RECT 72.370 91.065 72.645 91.205 ;
        RECT 72.815 90.865 73.005 92.225 ;
        RECT 73.185 91.860 73.695 92.395 ;
        RECT 73.915 91.585 74.160 92.190 ;
        RECT 75.730 91.615 76.230 92.225 ;
        RECT 73.205 91.415 74.435 91.585 ;
        RECT 71.995 90.695 73.005 90.865 ;
        RECT 73.175 90.850 73.925 91.040 ;
        RECT 71.655 90.355 72.780 90.525 ;
        RECT 73.175 90.185 73.345 90.850 ;
        RECT 74.095 90.605 74.435 91.415 ;
        RECT 75.525 91.155 75.875 91.405 ;
        RECT 76.060 90.985 76.230 91.615 ;
        RECT 76.860 91.745 77.190 92.225 ;
        RECT 77.360 91.935 77.585 92.395 ;
        RECT 77.755 91.745 78.085 92.225 ;
        RECT 76.860 91.575 78.085 91.745 ;
        RECT 78.275 91.595 78.525 92.395 ;
        RECT 78.695 91.595 79.035 92.225 ;
        RECT 79.215 91.895 79.545 92.395 ;
        RECT 79.745 91.825 79.915 92.175 ;
        RECT 80.115 91.995 80.445 92.395 ;
        RECT 80.615 91.825 80.785 92.175 ;
        RECT 80.955 91.995 81.335 92.395 ;
        RECT 76.400 91.205 76.730 91.405 ;
        RECT 76.900 91.205 77.230 91.405 ;
        RECT 77.400 91.205 77.820 91.405 ;
        RECT 77.995 91.235 78.690 91.405 ;
        RECT 77.995 90.985 78.165 91.235 ;
        RECT 78.860 90.985 79.035 91.595 ;
        RECT 79.210 91.155 79.560 91.725 ;
        RECT 79.745 91.655 81.355 91.825 ;
        RECT 81.525 91.720 81.795 92.065 ;
        RECT 81.185 91.485 81.355 91.655 ;
        RECT 71.315 90.015 73.345 90.185 ;
        RECT 73.515 89.845 73.685 90.605 ;
        RECT 73.920 90.195 74.435 90.605 ;
        RECT 75.730 90.815 78.165 90.985 ;
        RECT 75.730 90.015 76.060 90.815 ;
        RECT 76.230 89.845 76.560 90.645 ;
        RECT 76.860 90.015 77.190 90.815 ;
        RECT 77.835 89.845 78.085 90.645 ;
        RECT 78.355 89.845 78.525 90.985 ;
        RECT 78.695 90.015 79.035 90.985 ;
        RECT 79.210 90.695 79.530 90.985 ;
        RECT 79.730 90.865 80.440 91.485 ;
        RECT 80.610 91.155 81.015 91.485 ;
        RECT 81.185 91.155 81.455 91.485 ;
        RECT 81.185 90.985 81.355 91.155 ;
        RECT 81.625 90.985 81.795 91.720 ;
        RECT 82.885 91.670 83.175 92.395 ;
        RECT 83.345 91.895 83.645 92.225 ;
        RECT 83.815 91.915 84.090 92.395 ;
        RECT 80.630 90.815 81.355 90.985 ;
        RECT 80.630 90.695 80.800 90.815 ;
        RECT 79.210 90.525 80.800 90.695 ;
        RECT 79.210 90.065 80.865 90.355 ;
        RECT 81.035 89.845 81.315 90.645 ;
        RECT 81.525 90.015 81.795 90.985 ;
        RECT 82.885 89.845 83.175 91.010 ;
        RECT 83.345 90.985 83.515 91.895 ;
        RECT 84.270 91.745 84.565 92.135 ;
        RECT 84.735 91.915 84.990 92.395 ;
        RECT 85.165 91.745 85.425 92.135 ;
        RECT 85.595 91.915 85.875 92.395 ;
        RECT 86.105 91.935 86.665 92.225 ;
        RECT 86.835 91.935 87.085 92.395 ;
        RECT 83.685 91.155 84.035 91.725 ;
        RECT 84.270 91.575 85.920 91.745 ;
        RECT 84.205 91.235 85.345 91.405 ;
        RECT 84.205 90.985 84.375 91.235 ;
        RECT 85.515 91.065 85.920 91.575 ;
        RECT 83.345 90.815 84.375 90.985 ;
        RECT 85.165 90.895 85.920 91.065 ;
        RECT 83.345 90.015 83.655 90.815 ;
        RECT 85.165 90.645 85.425 90.895 ;
        RECT 83.825 89.845 84.135 90.645 ;
        RECT 84.305 90.475 85.425 90.645 ;
        RECT 84.305 90.015 84.565 90.475 ;
        RECT 84.735 89.845 84.990 90.305 ;
        RECT 85.165 90.015 85.425 90.475 ;
        RECT 85.595 89.845 85.880 90.715 ;
        RECT 86.105 90.565 86.355 91.935 ;
        RECT 87.705 91.765 88.035 92.125 ;
        RECT 86.645 91.575 88.035 91.765 ;
        RECT 88.495 91.845 88.665 92.135 ;
        RECT 88.835 92.015 89.165 92.395 ;
        RECT 88.495 91.675 89.160 91.845 ;
        RECT 86.645 91.485 86.815 91.575 ;
        RECT 86.525 91.155 86.815 91.485 ;
        RECT 86.985 91.155 87.325 91.405 ;
        RECT 87.545 91.155 88.220 91.405 ;
        RECT 86.645 90.905 86.815 91.155 ;
        RECT 86.645 90.735 87.585 90.905 ;
        RECT 87.955 90.795 88.220 91.155 ;
        RECT 88.410 90.855 88.760 91.505 ;
        RECT 86.105 90.015 86.565 90.565 ;
        RECT 86.755 89.845 87.085 90.565 ;
        RECT 87.285 90.185 87.585 90.735 ;
        RECT 88.930 90.685 89.160 91.675 ;
        RECT 88.495 90.515 89.160 90.685 ;
        RECT 87.755 89.845 88.035 90.515 ;
        RECT 88.495 90.015 88.665 90.515 ;
        RECT 88.835 89.845 89.165 90.345 ;
        RECT 89.335 90.015 89.560 92.135 ;
        RECT 89.775 92.015 90.105 92.395 ;
        RECT 90.275 91.845 90.445 92.175 ;
        RECT 90.745 92.015 91.760 92.215 ;
        RECT 89.750 91.655 90.445 91.845 ;
        RECT 89.750 90.685 89.920 91.655 ;
        RECT 90.090 90.855 90.500 91.475 ;
        RECT 90.670 90.905 90.890 91.775 ;
        RECT 91.070 91.465 91.420 91.835 ;
        RECT 91.590 91.285 91.760 92.015 ;
        RECT 91.930 91.955 92.340 92.395 ;
        RECT 92.630 91.755 92.880 92.185 ;
        RECT 93.080 91.935 93.400 92.395 ;
        RECT 93.960 92.005 94.810 92.175 ;
        RECT 91.930 91.415 92.340 91.745 ;
        RECT 92.630 91.415 93.050 91.755 ;
        RECT 91.340 91.245 91.760 91.285 ;
        RECT 91.340 91.075 92.690 91.245 ;
        RECT 89.750 90.515 90.445 90.685 ;
        RECT 90.670 90.525 91.170 90.905 ;
        RECT 89.775 89.845 90.105 90.345 ;
        RECT 90.275 90.015 90.445 90.515 ;
        RECT 91.340 90.230 91.510 91.075 ;
        RECT 92.440 90.915 92.690 91.075 ;
        RECT 91.680 90.645 91.930 90.905 ;
        RECT 92.860 90.645 93.050 91.415 ;
        RECT 91.680 90.395 93.050 90.645 ;
        RECT 93.220 91.585 94.470 91.755 ;
        RECT 93.220 90.825 93.390 91.585 ;
        RECT 94.140 91.465 94.470 91.585 ;
        RECT 93.560 91.005 93.740 91.415 ;
        RECT 94.640 91.245 94.810 92.005 ;
        RECT 95.010 91.915 95.670 92.395 ;
        RECT 95.850 91.800 96.170 92.130 ;
        RECT 95.000 91.475 95.660 91.745 ;
        RECT 95.000 91.415 95.330 91.475 ;
        RECT 95.480 91.245 95.810 91.305 ;
        RECT 93.910 91.075 95.810 91.245 ;
        RECT 93.220 90.515 93.740 90.825 ;
        RECT 93.910 90.565 94.080 91.075 ;
        RECT 95.980 90.905 96.170 91.800 ;
        RECT 94.250 90.735 96.170 90.905 ;
        RECT 95.850 90.715 96.170 90.735 ;
        RECT 96.370 91.485 96.620 92.135 ;
        RECT 96.800 91.935 97.085 92.395 ;
        RECT 97.265 91.685 97.520 92.215 ;
        RECT 96.370 91.155 97.170 91.485 ;
        RECT 93.910 90.395 95.120 90.565 ;
        RECT 90.680 90.060 91.510 90.230 ;
        RECT 91.750 89.845 92.130 90.225 ;
        RECT 92.310 90.105 92.480 90.395 ;
        RECT 93.910 90.315 94.080 90.395 ;
        RECT 92.650 89.845 92.980 90.225 ;
        RECT 93.450 90.065 94.080 90.315 ;
        RECT 94.260 89.845 94.680 90.225 ;
        RECT 94.880 90.105 95.120 90.395 ;
        RECT 95.350 89.845 95.680 90.535 ;
        RECT 95.850 90.105 96.020 90.715 ;
        RECT 96.370 90.565 96.620 91.155 ;
        RECT 97.340 90.825 97.520 91.685 ;
        RECT 99.075 91.845 99.245 92.135 ;
        RECT 99.415 92.015 99.745 92.395 ;
        RECT 99.075 91.675 99.740 91.845 ;
        RECT 98.990 90.855 99.340 91.505 ;
        RECT 96.290 90.055 96.620 90.565 ;
        RECT 96.800 89.845 97.085 90.645 ;
        RECT 97.265 90.355 97.520 90.825 ;
        RECT 99.510 90.685 99.740 91.675 ;
        RECT 99.075 90.515 99.740 90.685 ;
        RECT 97.265 90.185 97.605 90.355 ;
        RECT 97.265 90.155 97.520 90.185 ;
        RECT 99.075 90.015 99.245 90.515 ;
        RECT 99.415 89.845 99.745 90.345 ;
        RECT 99.915 90.015 100.140 92.135 ;
        RECT 100.355 92.015 100.685 92.395 ;
        RECT 100.855 91.845 101.025 92.175 ;
        RECT 101.325 92.015 102.340 92.215 ;
        RECT 100.330 91.655 101.025 91.845 ;
        RECT 100.330 90.685 100.500 91.655 ;
        RECT 100.670 90.855 101.080 91.475 ;
        RECT 101.250 90.905 101.470 91.775 ;
        RECT 101.650 91.465 102.000 91.835 ;
        RECT 102.170 91.285 102.340 92.015 ;
        RECT 102.510 91.955 102.920 92.395 ;
        RECT 103.210 91.755 103.460 92.185 ;
        RECT 103.660 91.935 103.980 92.395 ;
        RECT 104.540 92.005 105.390 92.175 ;
        RECT 102.510 91.415 102.920 91.745 ;
        RECT 103.210 91.415 103.630 91.755 ;
        RECT 101.920 91.245 102.340 91.285 ;
        RECT 101.920 91.075 103.270 91.245 ;
        RECT 100.330 90.515 101.025 90.685 ;
        RECT 101.250 90.525 101.750 90.905 ;
        RECT 100.355 89.845 100.685 90.345 ;
        RECT 100.855 90.015 101.025 90.515 ;
        RECT 101.920 90.230 102.090 91.075 ;
        RECT 103.020 90.915 103.270 91.075 ;
        RECT 102.260 90.645 102.510 90.905 ;
        RECT 103.440 90.645 103.630 91.415 ;
        RECT 102.260 90.395 103.630 90.645 ;
        RECT 103.800 91.585 105.050 91.755 ;
        RECT 103.800 90.825 103.970 91.585 ;
        RECT 104.720 91.465 105.050 91.585 ;
        RECT 104.140 91.005 104.320 91.415 ;
        RECT 105.220 91.245 105.390 92.005 ;
        RECT 105.590 91.915 106.250 92.395 ;
        RECT 106.430 91.800 106.750 92.130 ;
        RECT 105.580 91.475 106.240 91.745 ;
        RECT 105.580 91.415 105.910 91.475 ;
        RECT 106.060 91.245 106.390 91.305 ;
        RECT 104.490 91.075 106.390 91.245 ;
        RECT 103.800 90.515 104.320 90.825 ;
        RECT 104.490 90.565 104.660 91.075 ;
        RECT 106.560 90.905 106.750 91.800 ;
        RECT 104.830 90.735 106.750 90.905 ;
        RECT 106.430 90.715 106.750 90.735 ;
        RECT 106.950 91.485 107.200 92.135 ;
        RECT 107.380 91.935 107.665 92.395 ;
        RECT 107.845 91.685 108.100 92.215 ;
        RECT 106.950 91.155 107.750 91.485 ;
        RECT 104.490 90.395 105.700 90.565 ;
        RECT 101.260 90.060 102.090 90.230 ;
        RECT 102.330 89.845 102.710 90.225 ;
        RECT 102.890 90.105 103.060 90.395 ;
        RECT 104.490 90.315 104.660 90.395 ;
        RECT 103.230 89.845 103.560 90.225 ;
        RECT 104.030 90.065 104.660 90.315 ;
        RECT 104.840 89.845 105.260 90.225 ;
        RECT 105.460 90.105 105.700 90.395 ;
        RECT 105.930 89.845 106.260 90.535 ;
        RECT 106.430 90.105 106.600 90.715 ;
        RECT 106.950 90.565 107.200 91.155 ;
        RECT 107.920 90.825 108.100 91.685 ;
        RECT 108.645 91.670 108.935 92.395 ;
        RECT 109.105 91.720 109.365 92.225 ;
        RECT 109.545 92.015 109.875 92.395 ;
        RECT 110.055 91.845 110.225 92.225 ;
        RECT 106.870 90.055 107.200 90.565 ;
        RECT 107.380 89.845 107.665 90.645 ;
        RECT 107.845 90.355 108.100 90.825 ;
        RECT 107.845 90.185 108.185 90.355 ;
        RECT 107.845 90.155 108.100 90.185 ;
        RECT 108.645 89.845 108.935 91.010 ;
        RECT 109.105 90.920 109.275 91.720 ;
        RECT 109.560 91.675 110.225 91.845 ;
        RECT 109.560 91.420 109.730 91.675 ;
        RECT 110.525 91.575 110.755 92.395 ;
        RECT 110.925 91.595 111.255 92.225 ;
        RECT 109.445 91.090 109.730 91.420 ;
        RECT 109.965 91.125 110.295 91.495 ;
        RECT 110.505 91.155 110.835 91.405 ;
        RECT 109.560 90.945 109.730 91.090 ;
        RECT 111.005 90.995 111.255 91.595 ;
        RECT 111.425 91.575 111.635 92.395 ;
        RECT 112.325 91.645 113.535 92.395 ;
        RECT 109.105 90.015 109.375 90.920 ;
        RECT 109.560 90.775 110.225 90.945 ;
        RECT 109.545 89.845 109.875 90.605 ;
        RECT 110.055 90.015 110.225 90.775 ;
        RECT 110.525 89.845 110.755 90.985 ;
        RECT 110.925 90.015 111.255 90.995 ;
        RECT 111.425 89.845 111.635 90.985 ;
        RECT 112.325 90.935 112.845 91.475 ;
        RECT 113.015 91.105 113.535 91.645 ;
        RECT 112.325 89.845 113.535 90.935 ;
        RECT 5.520 89.675 113.620 89.845 ;
        RECT 5.605 88.585 6.815 89.675 ;
        RECT 6.985 88.585 8.655 89.675 ;
        RECT 8.915 89.005 9.085 89.505 ;
        RECT 9.255 89.175 9.585 89.675 ;
        RECT 8.915 88.835 9.580 89.005 ;
        RECT 5.605 87.875 6.125 88.415 ;
        RECT 6.295 88.045 6.815 88.585 ;
        RECT 6.985 87.895 7.735 88.415 ;
        RECT 7.905 88.065 8.655 88.585 ;
        RECT 8.830 88.015 9.180 88.665 ;
        RECT 5.605 87.125 6.815 87.875 ;
        RECT 6.985 87.125 8.655 87.895 ;
        RECT 9.350 87.845 9.580 88.835 ;
        RECT 8.915 87.675 9.580 87.845 ;
        RECT 8.915 87.385 9.085 87.675 ;
        RECT 9.255 87.125 9.585 87.505 ;
        RECT 9.755 87.385 9.980 89.505 ;
        RECT 10.195 89.175 10.525 89.675 ;
        RECT 10.695 89.005 10.865 89.505 ;
        RECT 11.100 89.290 11.930 89.460 ;
        RECT 12.170 89.295 12.550 89.675 ;
        RECT 10.170 88.835 10.865 89.005 ;
        RECT 10.170 87.865 10.340 88.835 ;
        RECT 10.510 88.045 10.920 88.665 ;
        RECT 11.090 88.615 11.590 88.995 ;
        RECT 10.170 87.675 10.865 87.865 ;
        RECT 11.090 87.745 11.310 88.615 ;
        RECT 11.760 88.445 11.930 89.290 ;
        RECT 12.730 89.125 12.900 89.415 ;
        RECT 13.070 89.295 13.400 89.675 ;
        RECT 13.870 89.205 14.500 89.455 ;
        RECT 14.680 89.295 15.100 89.675 ;
        RECT 14.330 89.125 14.500 89.205 ;
        RECT 15.300 89.125 15.540 89.415 ;
        RECT 12.100 88.875 13.470 89.125 ;
        RECT 12.100 88.615 12.350 88.875 ;
        RECT 12.860 88.445 13.110 88.605 ;
        RECT 11.760 88.275 13.110 88.445 ;
        RECT 11.760 88.235 12.180 88.275 ;
        RECT 11.490 87.685 11.840 88.055 ;
        RECT 10.195 87.125 10.525 87.505 ;
        RECT 10.695 87.345 10.865 87.675 ;
        RECT 12.010 87.505 12.180 88.235 ;
        RECT 13.280 88.105 13.470 88.875 ;
        RECT 12.350 87.775 12.760 88.105 ;
        RECT 13.050 87.765 13.470 88.105 ;
        RECT 13.640 88.695 14.160 89.005 ;
        RECT 14.330 88.955 15.540 89.125 ;
        RECT 15.770 88.985 16.100 89.675 ;
        RECT 13.640 87.935 13.810 88.695 ;
        RECT 13.980 88.105 14.160 88.515 ;
        RECT 14.330 88.445 14.500 88.955 ;
        RECT 16.270 88.805 16.440 89.415 ;
        RECT 16.710 88.955 17.040 89.465 ;
        RECT 16.270 88.785 16.590 88.805 ;
        RECT 14.670 88.615 16.590 88.785 ;
        RECT 14.330 88.275 16.230 88.445 ;
        RECT 14.560 87.935 14.890 88.055 ;
        RECT 13.640 87.765 14.890 87.935 ;
        RECT 11.165 87.305 12.180 87.505 ;
        RECT 12.350 87.125 12.760 87.565 ;
        RECT 13.050 87.335 13.300 87.765 ;
        RECT 13.500 87.125 13.820 87.585 ;
        RECT 15.060 87.515 15.230 88.275 ;
        RECT 15.900 88.215 16.230 88.275 ;
        RECT 15.420 88.045 15.750 88.105 ;
        RECT 15.420 87.775 16.080 88.045 ;
        RECT 16.400 87.720 16.590 88.615 ;
        RECT 14.380 87.345 15.230 87.515 ;
        RECT 15.430 87.125 16.090 87.605 ;
        RECT 16.270 87.390 16.590 87.720 ;
        RECT 16.790 88.365 17.040 88.955 ;
        RECT 17.220 88.875 17.505 89.675 ;
        RECT 17.685 88.995 17.940 89.365 ;
        RECT 17.685 88.825 18.025 88.995 ;
        RECT 17.685 88.695 17.940 88.825 ;
        RECT 16.790 88.035 17.590 88.365 ;
        RECT 16.790 87.385 17.040 88.035 ;
        RECT 17.760 87.835 17.940 88.695 ;
        RECT 18.485 88.510 18.775 89.675 ;
        RECT 18.950 88.535 19.285 89.505 ;
        RECT 19.455 88.535 19.625 89.675 ;
        RECT 19.795 89.335 21.825 89.505 ;
        RECT 18.950 87.865 19.120 88.535 ;
        RECT 19.795 88.365 19.965 89.335 ;
        RECT 19.290 88.035 19.545 88.365 ;
        RECT 19.770 88.035 19.965 88.365 ;
        RECT 20.135 88.995 21.260 89.165 ;
        RECT 19.375 87.865 19.545 88.035 ;
        RECT 20.135 87.865 20.305 88.995 ;
        RECT 17.220 87.125 17.505 87.585 ;
        RECT 17.685 87.305 17.940 87.835 ;
        RECT 18.485 87.125 18.775 87.850 ;
        RECT 18.950 87.295 19.205 87.865 ;
        RECT 19.375 87.695 20.305 87.865 ;
        RECT 20.475 88.655 21.485 88.825 ;
        RECT 20.475 87.855 20.645 88.655 ;
        RECT 20.850 88.315 21.125 88.455 ;
        RECT 20.845 88.145 21.125 88.315 ;
        RECT 20.130 87.660 20.305 87.695 ;
        RECT 19.375 87.125 19.705 87.525 ;
        RECT 20.130 87.295 20.660 87.660 ;
        RECT 20.850 87.295 21.125 88.145 ;
        RECT 21.295 87.295 21.485 88.655 ;
        RECT 21.655 88.670 21.825 89.335 ;
        RECT 21.995 88.915 22.165 89.675 ;
        RECT 22.400 88.915 22.915 89.325 ;
        RECT 21.655 88.480 22.405 88.670 ;
        RECT 22.575 88.105 22.915 88.915 ;
        RECT 21.685 87.935 22.915 88.105 ;
        RECT 23.085 88.955 23.545 89.505 ;
        RECT 23.735 88.955 24.065 89.675 ;
        RECT 21.665 87.125 22.175 87.660 ;
        RECT 22.395 87.330 22.640 87.935 ;
        RECT 23.085 87.585 23.335 88.955 ;
        RECT 24.265 88.785 24.565 89.335 ;
        RECT 24.735 89.005 25.015 89.675 ;
        RECT 23.625 88.615 24.565 88.785 ;
        RECT 23.625 88.365 23.795 88.615 ;
        RECT 24.935 88.365 25.200 88.725 ;
        RECT 25.385 88.585 26.595 89.675 ;
        RECT 26.965 89.005 27.245 89.675 ;
        RECT 27.415 88.785 27.715 89.335 ;
        RECT 27.915 88.955 28.245 89.675 ;
        RECT 28.435 88.955 28.895 89.505 ;
        RECT 29.065 89.240 34.410 89.675 ;
        RECT 23.505 88.035 23.795 88.365 ;
        RECT 23.965 88.115 24.305 88.365 ;
        RECT 24.525 88.115 25.200 88.365 ;
        RECT 23.625 87.945 23.795 88.035 ;
        RECT 23.625 87.755 25.015 87.945 ;
        RECT 23.085 87.295 23.645 87.585 ;
        RECT 23.815 87.125 24.065 87.585 ;
        RECT 24.685 87.395 25.015 87.755 ;
        RECT 25.385 87.875 25.905 88.415 ;
        RECT 26.075 88.045 26.595 88.585 ;
        RECT 26.780 88.365 27.045 88.725 ;
        RECT 27.415 88.615 28.355 88.785 ;
        RECT 28.185 88.365 28.355 88.615 ;
        RECT 26.780 88.115 27.455 88.365 ;
        RECT 27.675 88.115 28.015 88.365 ;
        RECT 28.185 88.035 28.475 88.365 ;
        RECT 28.185 87.945 28.355 88.035 ;
        RECT 25.385 87.125 26.595 87.875 ;
        RECT 26.965 87.755 28.355 87.945 ;
        RECT 26.965 87.395 27.295 87.755 ;
        RECT 28.645 87.585 28.895 88.955 ;
        RECT 30.650 87.670 30.990 88.500 ;
        RECT 32.470 87.990 32.820 89.240 ;
        RECT 34.585 88.585 38.095 89.675 ;
        RECT 38.265 88.585 39.475 89.675 ;
        RECT 34.585 87.895 36.235 88.415 ;
        RECT 36.405 88.065 38.095 88.585 ;
        RECT 27.915 87.125 28.165 87.585 ;
        RECT 28.335 87.295 28.895 87.585 ;
        RECT 29.065 87.125 34.410 87.670 ;
        RECT 34.585 87.125 38.095 87.895 ;
        RECT 38.265 87.875 38.785 88.415 ;
        RECT 38.955 88.045 39.475 88.585 ;
        RECT 39.645 88.600 39.915 89.505 ;
        RECT 40.085 88.915 40.415 89.675 ;
        RECT 40.595 88.745 40.765 89.505 ;
        RECT 38.265 87.125 39.475 87.875 ;
        RECT 39.645 87.800 39.815 88.600 ;
        RECT 40.100 88.575 40.765 88.745 ;
        RECT 41.025 88.585 43.615 89.675 ;
        RECT 40.100 88.430 40.270 88.575 ;
        RECT 39.985 88.100 40.270 88.430 ;
        RECT 40.100 87.845 40.270 88.100 ;
        RECT 40.505 88.025 40.835 88.395 ;
        RECT 41.025 87.895 42.235 88.415 ;
        RECT 42.405 88.065 43.615 88.585 ;
        RECT 44.245 88.510 44.535 89.675 ;
        RECT 44.705 88.585 48.215 89.675 ;
        RECT 44.705 87.895 46.355 88.415 ;
        RECT 46.525 88.065 48.215 88.585 ;
        RECT 49.305 88.535 49.575 89.505 ;
        RECT 49.785 88.875 50.065 89.675 ;
        RECT 50.235 89.165 51.890 89.455 ;
        RECT 50.300 88.825 51.890 88.995 ;
        RECT 50.300 88.705 50.470 88.825 ;
        RECT 49.745 88.535 50.470 88.705 ;
        RECT 39.645 87.295 39.905 87.800 ;
        RECT 40.100 87.675 40.765 87.845 ;
        RECT 40.085 87.125 40.415 87.505 ;
        RECT 40.595 87.295 40.765 87.675 ;
        RECT 41.025 87.125 43.615 87.895 ;
        RECT 44.245 87.125 44.535 87.850 ;
        RECT 44.705 87.125 48.215 87.895 ;
        RECT 49.305 87.800 49.475 88.535 ;
        RECT 49.745 88.365 49.915 88.535 ;
        RECT 49.645 88.035 49.915 88.365 ;
        RECT 50.085 88.035 50.490 88.365 ;
        RECT 50.660 88.035 51.370 88.655 ;
        RECT 51.570 88.535 51.890 88.825 ;
        RECT 52.065 88.585 54.655 89.675 ;
        RECT 54.915 89.005 55.085 89.505 ;
        RECT 55.255 89.175 55.585 89.675 ;
        RECT 54.915 88.835 55.580 89.005 ;
        RECT 49.745 87.865 49.915 88.035 ;
        RECT 49.305 87.455 49.575 87.800 ;
        RECT 49.745 87.695 51.355 87.865 ;
        RECT 51.540 87.795 51.890 88.365 ;
        RECT 52.065 87.895 53.275 88.415 ;
        RECT 53.445 88.065 54.655 88.585 ;
        RECT 54.830 88.015 55.180 88.665 ;
        RECT 49.765 87.125 50.145 87.525 ;
        RECT 50.315 87.345 50.485 87.695 ;
        RECT 50.655 87.125 50.985 87.525 ;
        RECT 51.185 87.345 51.355 87.695 ;
        RECT 51.555 87.125 51.885 87.625 ;
        RECT 52.065 87.125 54.655 87.895 ;
        RECT 55.350 87.845 55.580 88.835 ;
        RECT 54.915 87.675 55.580 87.845 ;
        RECT 54.915 87.385 55.085 87.675 ;
        RECT 55.255 87.125 55.585 87.505 ;
        RECT 55.755 87.385 55.980 89.505 ;
        RECT 56.195 89.175 56.525 89.675 ;
        RECT 56.695 89.005 56.865 89.505 ;
        RECT 57.100 89.290 57.930 89.460 ;
        RECT 58.170 89.295 58.550 89.675 ;
        RECT 56.170 88.835 56.865 89.005 ;
        RECT 56.170 87.865 56.340 88.835 ;
        RECT 56.510 88.045 56.920 88.665 ;
        RECT 57.090 88.615 57.590 88.995 ;
        RECT 56.170 87.675 56.865 87.865 ;
        RECT 57.090 87.745 57.310 88.615 ;
        RECT 57.760 88.445 57.930 89.290 ;
        RECT 58.730 89.125 58.900 89.415 ;
        RECT 59.070 89.295 59.400 89.675 ;
        RECT 59.870 89.205 60.500 89.455 ;
        RECT 60.680 89.295 61.100 89.675 ;
        RECT 60.330 89.125 60.500 89.205 ;
        RECT 61.300 89.125 61.540 89.415 ;
        RECT 58.100 88.875 59.470 89.125 ;
        RECT 58.100 88.615 58.350 88.875 ;
        RECT 58.860 88.445 59.110 88.605 ;
        RECT 57.760 88.275 59.110 88.445 ;
        RECT 57.760 88.235 58.180 88.275 ;
        RECT 57.490 87.685 57.840 88.055 ;
        RECT 56.195 87.125 56.525 87.505 ;
        RECT 56.695 87.345 56.865 87.675 ;
        RECT 58.010 87.505 58.180 88.235 ;
        RECT 59.280 88.105 59.470 88.875 ;
        RECT 58.350 87.775 58.760 88.105 ;
        RECT 59.050 87.765 59.470 88.105 ;
        RECT 59.640 88.695 60.160 89.005 ;
        RECT 60.330 88.955 61.540 89.125 ;
        RECT 61.770 88.985 62.100 89.675 ;
        RECT 59.640 87.935 59.810 88.695 ;
        RECT 59.980 88.105 60.160 88.515 ;
        RECT 60.330 88.445 60.500 88.955 ;
        RECT 62.270 88.805 62.440 89.415 ;
        RECT 62.710 88.955 63.040 89.465 ;
        RECT 62.270 88.785 62.590 88.805 ;
        RECT 60.670 88.615 62.590 88.785 ;
        RECT 60.330 88.275 62.230 88.445 ;
        RECT 60.560 87.935 60.890 88.055 ;
        RECT 59.640 87.765 60.890 87.935 ;
        RECT 57.165 87.305 58.180 87.505 ;
        RECT 58.350 87.125 58.760 87.565 ;
        RECT 59.050 87.335 59.300 87.765 ;
        RECT 59.500 87.125 59.820 87.585 ;
        RECT 61.060 87.515 61.230 88.275 ;
        RECT 61.900 88.215 62.230 88.275 ;
        RECT 61.420 88.045 61.750 88.105 ;
        RECT 61.420 87.775 62.080 88.045 ;
        RECT 62.400 87.720 62.590 88.615 ;
        RECT 60.380 87.345 61.230 87.515 ;
        RECT 61.430 87.125 62.090 87.605 ;
        RECT 62.270 87.390 62.590 87.720 ;
        RECT 62.790 88.365 63.040 88.955 ;
        RECT 63.220 88.875 63.505 89.675 ;
        RECT 63.685 88.695 63.940 89.365 ;
        RECT 62.790 88.035 63.590 88.365 ;
        RECT 62.790 87.385 63.040 88.035 ;
        RECT 63.760 87.835 63.940 88.695 ;
        RECT 63.685 87.635 63.940 87.835 ;
        RECT 64.485 88.705 64.755 89.475 ;
        RECT 64.925 88.895 65.255 89.675 ;
        RECT 65.460 89.070 65.645 89.475 ;
        RECT 65.815 89.250 66.150 89.675 ;
        RECT 65.460 88.895 66.125 89.070 ;
        RECT 64.485 88.535 65.615 88.705 ;
        RECT 63.220 87.125 63.505 87.585 ;
        RECT 63.685 87.465 64.025 87.635 ;
        RECT 64.485 87.625 64.655 88.535 ;
        RECT 64.825 87.785 65.185 88.365 ;
        RECT 65.365 88.035 65.615 88.535 ;
        RECT 65.785 87.865 66.125 88.895 ;
        RECT 65.440 87.695 66.125 87.865 ;
        RECT 67.245 88.600 67.515 89.505 ;
        RECT 67.685 88.915 68.015 89.675 ;
        RECT 68.195 88.745 68.365 89.505 ;
        RECT 67.245 87.800 67.415 88.600 ;
        RECT 67.700 88.575 68.365 88.745 ;
        RECT 68.625 88.585 69.835 89.675 ;
        RECT 67.700 88.430 67.870 88.575 ;
        RECT 67.585 88.100 67.870 88.430 ;
        RECT 67.700 87.845 67.870 88.100 ;
        RECT 68.105 88.025 68.435 88.395 ;
        RECT 68.625 87.875 69.145 88.415 ;
        RECT 69.315 88.045 69.835 88.585 ;
        RECT 70.005 88.510 70.295 89.675 ;
        RECT 70.465 88.585 73.975 89.675 ;
        RECT 70.465 87.895 72.115 88.415 ;
        RECT 72.285 88.065 73.975 88.585 ;
        RECT 74.350 88.705 74.680 89.505 ;
        RECT 74.850 88.875 75.180 89.675 ;
        RECT 75.480 88.705 75.810 89.505 ;
        RECT 76.455 88.875 76.705 89.675 ;
        RECT 74.350 88.535 76.785 88.705 ;
        RECT 76.975 88.535 77.145 89.675 ;
        RECT 77.315 88.535 77.655 89.505 ;
        RECT 78.290 89.165 79.945 89.455 ;
        RECT 78.290 88.825 79.880 88.995 ;
        RECT 80.115 88.875 80.395 89.675 ;
        RECT 78.290 88.535 78.610 88.825 ;
        RECT 79.710 88.705 79.880 88.825 ;
        RECT 74.145 88.115 74.495 88.365 ;
        RECT 74.680 87.905 74.850 88.535 ;
        RECT 75.020 88.115 75.350 88.315 ;
        RECT 75.520 88.115 75.850 88.315 ;
        RECT 76.020 88.115 76.440 88.315 ;
        RECT 76.615 88.285 76.785 88.535 ;
        RECT 76.615 88.115 77.310 88.285 ;
        RECT 63.685 87.305 63.940 87.465 ;
        RECT 64.485 87.295 64.745 87.625 ;
        RECT 64.955 87.125 65.230 87.605 ;
        RECT 65.440 87.295 65.645 87.695 ;
        RECT 65.815 87.125 66.150 87.525 ;
        RECT 67.245 87.295 67.505 87.800 ;
        RECT 67.700 87.675 68.365 87.845 ;
        RECT 67.685 87.125 68.015 87.505 ;
        RECT 68.195 87.295 68.365 87.675 ;
        RECT 68.625 87.125 69.835 87.875 ;
        RECT 70.005 87.125 70.295 87.850 ;
        RECT 70.465 87.125 73.975 87.895 ;
        RECT 74.350 87.295 74.850 87.905 ;
        RECT 75.480 87.775 76.705 87.945 ;
        RECT 77.480 87.925 77.655 88.535 ;
        RECT 78.805 88.485 79.520 88.655 ;
        RECT 79.710 88.535 80.435 88.705 ;
        RECT 80.605 88.535 80.875 89.505 ;
        RECT 81.050 89.165 82.705 89.455 ;
        RECT 81.050 88.825 82.640 88.995 ;
        RECT 82.875 88.875 83.155 89.675 ;
        RECT 81.050 88.535 81.370 88.825 ;
        RECT 82.470 88.705 82.640 88.825 ;
        RECT 75.480 87.295 75.810 87.775 ;
        RECT 75.980 87.125 76.205 87.585 ;
        RECT 76.375 87.295 76.705 87.775 ;
        RECT 76.895 87.125 77.145 87.925 ;
        RECT 77.315 87.295 77.655 87.925 ;
        RECT 78.290 87.795 78.640 88.365 ;
        RECT 78.810 88.035 79.520 88.485 ;
        RECT 80.265 88.365 80.435 88.535 ;
        RECT 79.690 88.035 80.095 88.365 ;
        RECT 80.265 88.035 80.535 88.365 ;
        RECT 80.265 87.865 80.435 88.035 ;
        RECT 78.825 87.695 80.435 87.865 ;
        RECT 80.705 87.800 80.875 88.535 ;
        RECT 81.565 88.485 82.280 88.655 ;
        RECT 82.470 88.535 83.195 88.705 ;
        RECT 83.365 88.535 83.635 89.505 ;
        RECT 83.805 88.585 85.015 89.675 ;
        RECT 85.190 89.165 86.845 89.455 ;
        RECT 78.295 87.125 78.625 87.625 ;
        RECT 78.825 87.345 78.995 87.695 ;
        RECT 79.195 87.125 79.525 87.525 ;
        RECT 79.695 87.345 79.865 87.695 ;
        RECT 80.035 87.125 80.415 87.525 ;
        RECT 80.605 87.455 80.875 87.800 ;
        RECT 81.050 87.795 81.400 88.365 ;
        RECT 81.570 88.035 82.280 88.485 ;
        RECT 83.025 88.365 83.195 88.535 ;
        RECT 82.450 88.035 82.855 88.365 ;
        RECT 83.025 88.035 83.295 88.365 ;
        RECT 83.025 87.865 83.195 88.035 ;
        RECT 81.585 87.695 83.195 87.865 ;
        RECT 83.465 87.800 83.635 88.535 ;
        RECT 81.055 87.125 81.385 87.625 ;
        RECT 81.585 87.345 81.755 87.695 ;
        RECT 81.955 87.125 82.285 87.525 ;
        RECT 82.455 87.345 82.625 87.695 ;
        RECT 82.795 87.125 83.175 87.525 ;
        RECT 83.365 87.455 83.635 87.800 ;
        RECT 83.805 87.875 84.325 88.415 ;
        RECT 84.495 88.045 85.015 88.585 ;
        RECT 85.190 88.825 86.780 88.995 ;
        RECT 87.015 88.875 87.295 89.675 ;
        RECT 85.190 88.535 85.510 88.825 ;
        RECT 86.610 88.705 86.780 88.825 ;
        RECT 83.805 87.125 85.015 87.875 ;
        RECT 85.190 87.795 85.540 88.365 ;
        RECT 85.710 88.035 86.420 88.655 ;
        RECT 86.610 88.535 87.335 88.705 ;
        RECT 87.505 88.535 87.775 89.505 ;
        RECT 87.165 88.365 87.335 88.535 ;
        RECT 86.590 88.035 86.995 88.365 ;
        RECT 87.165 88.035 87.435 88.365 ;
        RECT 87.165 87.865 87.335 88.035 ;
        RECT 85.725 87.695 87.335 87.865 ;
        RECT 87.605 87.800 87.775 88.535 ;
        RECT 85.195 87.125 85.525 87.625 ;
        RECT 85.725 87.345 85.895 87.695 ;
        RECT 86.095 87.125 86.425 87.525 ;
        RECT 86.595 87.345 86.765 87.695 ;
        RECT 86.935 87.125 87.315 87.525 ;
        RECT 87.505 87.455 87.775 87.800 ;
        RECT 87.945 88.955 88.405 89.505 ;
        RECT 88.595 88.955 88.925 89.675 ;
        RECT 87.945 87.585 88.195 88.955 ;
        RECT 89.125 88.785 89.425 89.335 ;
        RECT 89.595 89.005 89.875 89.675 ;
        RECT 88.485 88.615 89.425 88.785 ;
        RECT 88.485 88.365 88.655 88.615 ;
        RECT 89.795 88.365 90.060 88.725 ;
        RECT 88.365 88.035 88.655 88.365 ;
        RECT 88.825 88.115 89.165 88.365 ;
        RECT 89.385 88.115 90.060 88.365 ;
        RECT 90.710 88.535 91.045 89.505 ;
        RECT 91.215 88.535 91.385 89.675 ;
        RECT 91.555 89.335 93.585 89.505 ;
        RECT 88.485 87.945 88.655 88.035 ;
        RECT 88.485 87.755 89.875 87.945 ;
        RECT 87.945 87.295 88.505 87.585 ;
        RECT 88.675 87.125 88.925 87.585 ;
        RECT 89.545 87.395 89.875 87.755 ;
        RECT 90.710 87.865 90.880 88.535 ;
        RECT 91.555 88.365 91.725 89.335 ;
        RECT 91.050 88.035 91.305 88.365 ;
        RECT 91.530 88.035 91.725 88.365 ;
        RECT 91.895 88.995 93.020 89.165 ;
        RECT 91.135 87.865 91.305 88.035 ;
        RECT 91.895 87.865 92.065 88.995 ;
        RECT 90.710 87.295 90.965 87.865 ;
        RECT 91.135 87.695 92.065 87.865 ;
        RECT 92.235 88.655 93.245 88.825 ;
        RECT 92.235 87.855 92.405 88.655 ;
        RECT 92.610 88.315 92.885 88.455 ;
        RECT 92.605 88.145 92.885 88.315 ;
        RECT 91.890 87.660 92.065 87.695 ;
        RECT 91.135 87.125 91.465 87.525 ;
        RECT 91.890 87.295 92.420 87.660 ;
        RECT 92.610 87.295 92.885 88.145 ;
        RECT 93.055 87.295 93.245 88.655 ;
        RECT 93.415 88.670 93.585 89.335 ;
        RECT 93.755 88.915 93.925 89.675 ;
        RECT 94.160 88.915 94.675 89.325 ;
        RECT 93.415 88.480 94.165 88.670 ;
        RECT 94.335 88.105 94.675 88.915 ;
        RECT 95.765 88.510 96.055 89.675 ;
        RECT 96.285 88.535 96.495 89.675 ;
        RECT 96.665 88.525 96.995 89.505 ;
        RECT 97.165 88.535 97.395 89.675 ;
        RECT 97.605 88.585 101.115 89.675 ;
        RECT 93.445 87.935 94.675 88.105 ;
        RECT 93.425 87.125 93.935 87.660 ;
        RECT 94.155 87.330 94.400 87.935 ;
        RECT 95.765 87.125 96.055 87.850 ;
        RECT 96.285 87.125 96.495 87.945 ;
        RECT 96.665 87.925 96.915 88.525 ;
        RECT 97.085 88.115 97.415 88.365 ;
        RECT 96.665 87.295 96.995 87.925 ;
        RECT 97.165 87.125 97.395 87.945 ;
        RECT 97.605 87.895 99.255 88.415 ;
        RECT 99.425 88.065 101.115 88.585 ;
        RECT 102.205 88.915 102.720 89.325 ;
        RECT 102.955 88.915 103.125 89.675 ;
        RECT 103.295 89.335 105.325 89.505 ;
        RECT 102.205 88.105 102.545 88.915 ;
        RECT 103.295 88.670 103.465 89.335 ;
        RECT 103.860 88.995 104.985 89.165 ;
        RECT 102.715 88.480 103.465 88.670 ;
        RECT 103.635 88.655 104.645 88.825 ;
        RECT 102.205 87.935 103.435 88.105 ;
        RECT 97.605 87.125 101.115 87.895 ;
        RECT 102.480 87.330 102.725 87.935 ;
        RECT 102.945 87.125 103.455 87.660 ;
        RECT 103.635 87.295 103.825 88.655 ;
        RECT 103.995 87.975 104.270 88.455 ;
        RECT 103.995 87.805 104.275 87.975 ;
        RECT 104.475 87.855 104.645 88.655 ;
        RECT 104.815 87.865 104.985 88.995 ;
        RECT 105.155 88.365 105.325 89.335 ;
        RECT 105.495 88.535 105.665 89.675 ;
        RECT 105.835 88.535 106.170 89.505 ;
        RECT 105.155 88.035 105.350 88.365 ;
        RECT 105.575 88.035 105.830 88.365 ;
        RECT 105.575 87.865 105.745 88.035 ;
        RECT 106.000 87.865 106.170 88.535 ;
        RECT 103.995 87.295 104.270 87.805 ;
        RECT 104.815 87.695 105.745 87.865 ;
        RECT 104.815 87.660 104.990 87.695 ;
        RECT 104.460 87.295 104.990 87.660 ;
        RECT 105.415 87.125 105.745 87.525 ;
        RECT 105.915 87.295 106.170 87.865 ;
        RECT 106.350 88.535 106.685 89.505 ;
        RECT 106.855 88.535 107.025 89.675 ;
        RECT 107.195 89.335 109.225 89.505 ;
        RECT 106.350 87.865 106.520 88.535 ;
        RECT 107.195 88.365 107.365 89.335 ;
        RECT 106.690 88.035 106.945 88.365 ;
        RECT 107.170 88.035 107.365 88.365 ;
        RECT 107.535 88.995 108.660 89.165 ;
        RECT 106.775 87.865 106.945 88.035 ;
        RECT 107.535 87.865 107.705 88.995 ;
        RECT 106.350 87.295 106.605 87.865 ;
        RECT 106.775 87.695 107.705 87.865 ;
        RECT 107.875 88.655 108.885 88.825 ;
        RECT 107.875 87.855 108.045 88.655 ;
        RECT 108.250 88.315 108.525 88.455 ;
        RECT 108.245 88.145 108.525 88.315 ;
        RECT 107.530 87.660 107.705 87.695 ;
        RECT 106.775 87.125 107.105 87.525 ;
        RECT 107.530 87.295 108.060 87.660 ;
        RECT 108.250 87.295 108.525 88.145 ;
        RECT 108.695 87.295 108.885 88.655 ;
        RECT 109.055 88.670 109.225 89.335 ;
        RECT 109.395 88.915 109.565 89.675 ;
        RECT 109.800 88.915 110.315 89.325 ;
        RECT 109.055 88.480 109.805 88.670 ;
        RECT 109.975 88.105 110.315 88.915 ;
        RECT 110.485 88.585 112.155 89.675 ;
        RECT 109.085 87.935 110.315 88.105 ;
        RECT 109.065 87.125 109.575 87.660 ;
        RECT 109.795 87.330 110.040 87.935 ;
        RECT 110.485 87.895 111.235 88.415 ;
        RECT 111.405 88.065 112.155 88.585 ;
        RECT 112.325 88.585 113.535 89.675 ;
        RECT 112.325 88.045 112.845 88.585 ;
        RECT 110.485 87.125 112.155 87.895 ;
        RECT 113.015 87.875 113.535 88.415 ;
        RECT 112.325 87.125 113.535 87.875 ;
        RECT 5.520 86.955 113.620 87.125 ;
        RECT 5.605 86.205 6.815 86.955 ;
        RECT 6.985 86.410 12.330 86.955 ;
        RECT 5.605 85.665 6.125 86.205 ;
        RECT 6.295 85.495 6.815 86.035 ;
        RECT 8.570 85.580 8.910 86.410 ;
        RECT 12.505 86.205 13.715 86.955 ;
        RECT 5.605 84.405 6.815 85.495 ;
        RECT 10.390 84.840 10.740 86.090 ;
        RECT 12.505 85.665 13.025 86.205 ;
        RECT 13.945 86.135 14.155 86.955 ;
        RECT 14.325 86.155 14.655 86.785 ;
        RECT 13.195 85.495 13.715 86.035 ;
        RECT 14.325 85.555 14.575 86.155 ;
        RECT 14.825 86.135 15.055 86.955 ;
        RECT 15.265 86.280 15.525 86.785 ;
        RECT 15.705 86.575 16.035 86.955 ;
        RECT 16.215 86.405 16.385 86.785 ;
        RECT 14.745 85.715 15.075 85.965 ;
        RECT 6.985 84.405 12.330 84.840 ;
        RECT 12.505 84.405 13.715 85.495 ;
        RECT 13.945 84.405 14.155 85.545 ;
        RECT 14.325 84.575 14.655 85.555 ;
        RECT 14.825 84.405 15.055 85.545 ;
        RECT 15.265 85.480 15.435 86.280 ;
        RECT 15.720 86.235 16.385 86.405 ;
        RECT 15.720 85.980 15.890 86.235 ;
        RECT 16.645 86.185 20.155 86.955 ;
        RECT 20.785 86.495 21.345 86.785 ;
        RECT 21.515 86.495 21.765 86.955 ;
        RECT 15.605 85.650 15.890 85.980 ;
        RECT 16.125 85.685 16.455 86.055 ;
        RECT 16.645 85.665 18.295 86.185 ;
        RECT 15.720 85.505 15.890 85.650 ;
        RECT 15.265 84.575 15.535 85.480 ;
        RECT 15.720 85.335 16.385 85.505 ;
        RECT 18.465 85.495 20.155 86.015 ;
        RECT 15.705 84.405 16.035 85.165 ;
        RECT 16.215 84.575 16.385 85.335 ;
        RECT 16.645 84.405 20.155 85.495 ;
        RECT 20.785 85.125 21.035 86.495 ;
        RECT 22.385 86.325 22.715 86.685 ;
        RECT 21.325 86.135 22.715 86.325 ;
        RECT 23.285 86.325 23.615 86.685 ;
        RECT 24.235 86.495 24.485 86.955 ;
        RECT 24.655 86.495 25.215 86.785 ;
        RECT 23.285 86.135 24.675 86.325 ;
        RECT 21.325 86.045 21.495 86.135 ;
        RECT 21.205 85.715 21.495 86.045 ;
        RECT 24.505 86.045 24.675 86.135 ;
        RECT 21.665 85.715 22.005 85.965 ;
        RECT 22.225 85.715 22.900 85.965 ;
        RECT 21.325 85.465 21.495 85.715 ;
        RECT 21.325 85.295 22.265 85.465 ;
        RECT 22.635 85.355 22.900 85.715 ;
        RECT 23.100 85.715 23.775 85.965 ;
        RECT 23.995 85.715 24.335 85.965 ;
        RECT 24.505 85.715 24.795 86.045 ;
        RECT 23.100 85.355 23.365 85.715 ;
        RECT 24.505 85.465 24.675 85.715 ;
        RECT 20.785 84.575 21.245 85.125 ;
        RECT 21.435 84.405 21.765 85.125 ;
        RECT 21.965 84.745 22.265 85.295 ;
        RECT 23.735 85.295 24.675 85.465 ;
        RECT 22.435 84.405 22.715 85.075 ;
        RECT 23.285 84.405 23.565 85.075 ;
        RECT 23.735 84.745 24.035 85.295 ;
        RECT 24.965 85.125 25.215 86.495 ;
        RECT 25.385 86.410 30.730 86.955 ;
        RECT 26.970 85.580 27.310 86.410 ;
        RECT 31.365 86.230 31.655 86.955 ;
        RECT 32.375 86.405 32.545 86.785 ;
        RECT 32.725 86.575 33.055 86.955 ;
        RECT 32.375 86.235 33.040 86.405 ;
        RECT 33.235 86.280 33.495 86.785 ;
        RECT 24.235 84.405 24.565 85.125 ;
        RECT 24.755 84.575 25.215 85.125 ;
        RECT 28.790 84.840 29.140 86.090 ;
        RECT 32.305 85.685 32.635 86.055 ;
        RECT 32.870 85.980 33.040 86.235 ;
        RECT 32.870 85.650 33.155 85.980 ;
        RECT 25.385 84.405 30.730 84.840 ;
        RECT 31.365 84.405 31.655 85.570 ;
        RECT 32.870 85.505 33.040 85.650 ;
        RECT 32.375 85.335 33.040 85.505 ;
        RECT 33.325 85.480 33.495 86.280 ;
        RECT 33.665 86.185 35.335 86.955 ;
        RECT 33.665 85.665 34.415 86.185 ;
        RECT 35.545 86.135 35.775 86.955 ;
        RECT 35.945 86.155 36.275 86.785 ;
        RECT 34.585 85.495 35.335 86.015 ;
        RECT 35.525 85.715 35.855 85.965 ;
        RECT 36.025 85.555 36.275 86.155 ;
        RECT 36.445 86.135 36.655 86.955 ;
        RECT 36.975 86.405 37.145 86.695 ;
        RECT 37.315 86.575 37.645 86.955 ;
        RECT 36.975 86.235 37.640 86.405 ;
        RECT 32.375 84.575 32.545 85.335 ;
        RECT 32.725 84.405 33.055 85.165 ;
        RECT 33.225 84.575 33.495 85.480 ;
        RECT 33.665 84.405 35.335 85.495 ;
        RECT 35.545 84.405 35.775 85.545 ;
        RECT 35.945 84.575 36.275 85.555 ;
        RECT 36.445 84.405 36.655 85.545 ;
        RECT 36.890 85.415 37.240 86.065 ;
        RECT 37.410 85.245 37.640 86.235 ;
        RECT 36.975 85.075 37.640 85.245 ;
        RECT 36.975 84.575 37.145 85.075 ;
        RECT 37.315 84.405 37.645 84.905 ;
        RECT 37.815 84.575 38.040 86.695 ;
        RECT 38.255 86.575 38.585 86.955 ;
        RECT 38.755 86.405 38.925 86.735 ;
        RECT 39.225 86.575 40.240 86.775 ;
        RECT 38.230 86.215 38.925 86.405 ;
        RECT 38.230 85.245 38.400 86.215 ;
        RECT 38.570 85.415 38.980 86.035 ;
        RECT 39.150 85.465 39.370 86.335 ;
        RECT 39.550 86.025 39.900 86.395 ;
        RECT 40.070 85.845 40.240 86.575 ;
        RECT 40.410 86.515 40.820 86.955 ;
        RECT 41.110 86.315 41.360 86.745 ;
        RECT 41.560 86.495 41.880 86.955 ;
        RECT 42.440 86.565 43.290 86.735 ;
        RECT 40.410 85.975 40.820 86.305 ;
        RECT 41.110 85.975 41.530 86.315 ;
        RECT 39.820 85.805 40.240 85.845 ;
        RECT 39.820 85.635 41.170 85.805 ;
        RECT 38.230 85.075 38.925 85.245 ;
        RECT 39.150 85.085 39.650 85.465 ;
        RECT 38.255 84.405 38.585 84.905 ;
        RECT 38.755 84.575 38.925 85.075 ;
        RECT 39.820 84.790 39.990 85.635 ;
        RECT 40.920 85.475 41.170 85.635 ;
        RECT 40.160 85.205 40.410 85.465 ;
        RECT 41.340 85.205 41.530 85.975 ;
        RECT 40.160 84.955 41.530 85.205 ;
        RECT 41.700 86.145 42.950 86.315 ;
        RECT 41.700 85.385 41.870 86.145 ;
        RECT 42.620 86.025 42.950 86.145 ;
        RECT 42.040 85.565 42.220 85.975 ;
        RECT 43.120 85.805 43.290 86.565 ;
        RECT 43.490 86.475 44.150 86.955 ;
        RECT 44.330 86.360 44.650 86.690 ;
        RECT 43.480 86.035 44.140 86.305 ;
        RECT 43.480 85.975 43.810 86.035 ;
        RECT 43.960 85.805 44.290 85.865 ;
        RECT 42.390 85.635 44.290 85.805 ;
        RECT 41.700 85.075 42.220 85.385 ;
        RECT 42.390 85.125 42.560 85.635 ;
        RECT 44.460 85.465 44.650 86.360 ;
        RECT 42.730 85.295 44.650 85.465 ;
        RECT 44.330 85.275 44.650 85.295 ;
        RECT 44.850 86.045 45.100 86.695 ;
        RECT 45.280 86.495 45.565 86.955 ;
        RECT 45.745 86.245 46.000 86.775 ;
        RECT 44.850 85.715 45.650 86.045 ;
        RECT 42.390 84.955 43.600 85.125 ;
        RECT 39.160 84.620 39.990 84.790 ;
        RECT 40.230 84.405 40.610 84.785 ;
        RECT 40.790 84.665 40.960 84.955 ;
        RECT 42.390 84.875 42.560 84.955 ;
        RECT 41.130 84.405 41.460 84.785 ;
        RECT 41.930 84.625 42.560 84.875 ;
        RECT 42.740 84.405 43.160 84.785 ;
        RECT 43.360 84.665 43.600 84.955 ;
        RECT 43.830 84.405 44.160 85.095 ;
        RECT 44.330 84.665 44.500 85.275 ;
        RECT 44.850 85.125 45.100 85.715 ;
        RECT 45.820 85.385 46.000 86.245 ;
        RECT 44.770 84.615 45.100 85.125 ;
        RECT 45.280 84.405 45.565 85.205 ;
        RECT 45.745 84.915 46.000 85.385 ;
        RECT 46.550 86.215 46.805 86.785 ;
        RECT 46.975 86.555 47.305 86.955 ;
        RECT 47.730 86.420 48.260 86.785 ;
        RECT 47.730 86.385 47.905 86.420 ;
        RECT 46.975 86.215 47.905 86.385 ;
        RECT 46.550 85.545 46.720 86.215 ;
        RECT 46.975 86.045 47.145 86.215 ;
        RECT 46.890 85.715 47.145 86.045 ;
        RECT 47.370 85.715 47.565 86.045 ;
        RECT 45.745 84.745 46.085 84.915 ;
        RECT 45.745 84.715 46.000 84.745 ;
        RECT 46.550 84.575 46.885 85.545 ;
        RECT 47.055 84.405 47.225 85.545 ;
        RECT 47.395 84.745 47.565 85.715 ;
        RECT 47.735 85.085 47.905 86.215 ;
        RECT 48.075 85.425 48.245 86.225 ;
        RECT 48.450 85.935 48.725 86.785 ;
        RECT 48.445 85.765 48.725 85.935 ;
        RECT 48.450 85.625 48.725 85.765 ;
        RECT 48.895 85.425 49.085 86.785 ;
        RECT 49.265 86.420 49.775 86.955 ;
        RECT 49.995 86.145 50.240 86.750 ;
        RECT 50.890 86.175 51.390 86.785 ;
        RECT 49.285 85.975 50.515 86.145 ;
        RECT 48.075 85.255 49.085 85.425 ;
        RECT 49.255 85.410 50.005 85.600 ;
        RECT 47.735 84.915 48.860 85.085 ;
        RECT 49.255 84.745 49.425 85.410 ;
        RECT 50.175 85.165 50.515 85.975 ;
        RECT 50.685 85.715 51.035 85.965 ;
        RECT 51.220 85.545 51.390 86.175 ;
        RECT 52.020 86.305 52.350 86.785 ;
        RECT 52.520 86.495 52.745 86.955 ;
        RECT 52.915 86.305 53.245 86.785 ;
        RECT 52.020 86.135 53.245 86.305 ;
        RECT 53.435 86.155 53.685 86.955 ;
        RECT 53.855 86.155 54.195 86.785 ;
        RECT 54.375 86.455 54.705 86.955 ;
        RECT 54.905 86.385 55.075 86.735 ;
        RECT 55.275 86.555 55.605 86.955 ;
        RECT 55.775 86.385 55.945 86.735 ;
        RECT 56.115 86.555 56.495 86.955 ;
        RECT 53.965 86.105 54.195 86.155 ;
        RECT 51.560 85.765 51.890 85.965 ;
        RECT 52.060 85.765 52.390 85.965 ;
        RECT 52.560 85.765 52.980 85.965 ;
        RECT 53.155 85.795 53.850 85.965 ;
        RECT 53.155 85.545 53.325 85.795 ;
        RECT 54.020 85.545 54.195 86.105 ;
        RECT 54.370 85.715 54.720 86.285 ;
        RECT 54.905 86.215 56.515 86.385 ;
        RECT 56.685 86.280 56.955 86.625 ;
        RECT 56.345 86.045 56.515 86.215 ;
        RECT 47.395 84.575 49.425 84.745 ;
        RECT 49.595 84.405 49.765 85.165 ;
        RECT 50.000 84.755 50.515 85.165 ;
        RECT 50.890 85.375 53.325 85.545 ;
        RECT 50.890 84.575 51.220 85.375 ;
        RECT 51.390 84.405 51.720 85.205 ;
        RECT 52.020 84.575 52.350 85.375 ;
        RECT 52.995 84.405 53.245 85.205 ;
        RECT 53.515 84.405 53.685 85.545 ;
        RECT 53.855 84.575 54.195 85.545 ;
        RECT 54.370 85.255 54.690 85.545 ;
        RECT 54.890 85.425 55.600 86.045 ;
        RECT 55.770 85.715 56.175 86.045 ;
        RECT 56.345 85.715 56.615 86.045 ;
        RECT 56.345 85.545 56.515 85.715 ;
        RECT 56.785 85.545 56.955 86.280 ;
        RECT 57.125 86.230 57.415 86.955 ;
        RECT 57.585 86.280 57.845 86.785 ;
        RECT 58.025 86.575 58.355 86.955 ;
        RECT 58.535 86.405 58.705 86.785 ;
        RECT 55.790 85.375 56.515 85.545 ;
        RECT 55.790 85.255 55.960 85.375 ;
        RECT 54.370 85.085 55.960 85.255 ;
        RECT 54.370 84.625 56.025 84.915 ;
        RECT 56.195 84.405 56.475 85.205 ;
        RECT 56.685 84.575 56.955 85.545 ;
        RECT 57.125 84.405 57.415 85.570 ;
        RECT 57.585 85.480 57.755 86.280 ;
        RECT 58.040 86.235 58.705 86.405 ;
        RECT 58.040 85.980 58.210 86.235 ;
        RECT 58.970 86.215 59.225 86.785 ;
        RECT 59.395 86.555 59.725 86.955 ;
        RECT 60.150 86.420 60.680 86.785 ;
        RECT 60.150 86.385 60.325 86.420 ;
        RECT 59.395 86.215 60.325 86.385 ;
        RECT 60.870 86.275 61.145 86.785 ;
        RECT 57.925 85.650 58.210 85.980 ;
        RECT 58.445 85.685 58.775 86.055 ;
        RECT 58.040 85.505 58.210 85.650 ;
        RECT 58.970 85.545 59.140 86.215 ;
        RECT 59.395 86.045 59.565 86.215 ;
        RECT 59.310 85.715 59.565 86.045 ;
        RECT 59.790 85.715 59.985 86.045 ;
        RECT 57.585 84.575 57.855 85.480 ;
        RECT 58.040 85.335 58.705 85.505 ;
        RECT 58.025 84.405 58.355 85.165 ;
        RECT 58.535 84.575 58.705 85.335 ;
        RECT 58.970 84.575 59.305 85.545 ;
        RECT 59.475 84.405 59.645 85.545 ;
        RECT 59.815 84.745 59.985 85.715 ;
        RECT 60.155 85.085 60.325 86.215 ;
        RECT 60.495 85.425 60.665 86.225 ;
        RECT 60.865 86.105 61.145 86.275 ;
        RECT 60.870 85.625 61.145 86.105 ;
        RECT 61.315 85.425 61.505 86.785 ;
        RECT 61.685 86.420 62.195 86.955 ;
        RECT 62.415 86.145 62.660 86.750 ;
        RECT 64.115 86.405 64.285 86.695 ;
        RECT 64.455 86.575 64.785 86.955 ;
        RECT 64.115 86.235 64.780 86.405 ;
        RECT 61.705 85.975 62.935 86.145 ;
        RECT 60.495 85.255 61.505 85.425 ;
        RECT 61.675 85.410 62.425 85.600 ;
        RECT 60.155 84.915 61.280 85.085 ;
        RECT 61.675 84.745 61.845 85.410 ;
        RECT 62.595 85.165 62.935 85.975 ;
        RECT 64.030 85.415 64.380 86.065 ;
        RECT 64.550 85.245 64.780 86.235 ;
        RECT 59.815 84.575 61.845 84.745 ;
        RECT 62.015 84.405 62.185 85.165 ;
        RECT 62.420 84.755 62.935 85.165 ;
        RECT 64.115 85.075 64.780 85.245 ;
        RECT 64.115 84.575 64.285 85.075 ;
        RECT 64.455 84.405 64.785 84.905 ;
        RECT 64.955 84.575 65.180 86.695 ;
        RECT 65.395 86.575 65.725 86.955 ;
        RECT 65.895 86.405 66.065 86.735 ;
        RECT 66.365 86.575 67.380 86.775 ;
        RECT 65.370 86.215 66.065 86.405 ;
        RECT 65.370 85.245 65.540 86.215 ;
        RECT 65.710 85.415 66.120 86.035 ;
        RECT 66.290 85.465 66.510 86.335 ;
        RECT 66.690 86.025 67.040 86.395 ;
        RECT 67.210 85.845 67.380 86.575 ;
        RECT 67.550 86.515 67.960 86.955 ;
        RECT 68.250 86.315 68.500 86.745 ;
        RECT 68.700 86.495 69.020 86.955 ;
        RECT 69.580 86.565 70.430 86.735 ;
        RECT 67.550 85.975 67.960 86.305 ;
        RECT 68.250 85.975 68.670 86.315 ;
        RECT 66.960 85.805 67.380 85.845 ;
        RECT 66.960 85.635 68.310 85.805 ;
        RECT 65.370 85.075 66.065 85.245 ;
        RECT 66.290 85.085 66.790 85.465 ;
        RECT 65.395 84.405 65.725 84.905 ;
        RECT 65.895 84.575 66.065 85.075 ;
        RECT 66.960 84.790 67.130 85.635 ;
        RECT 68.060 85.475 68.310 85.635 ;
        RECT 67.300 85.205 67.550 85.465 ;
        RECT 68.480 85.205 68.670 85.975 ;
        RECT 67.300 84.955 68.670 85.205 ;
        RECT 68.840 86.145 70.090 86.315 ;
        RECT 68.840 85.385 69.010 86.145 ;
        RECT 69.760 86.025 70.090 86.145 ;
        RECT 69.180 85.565 69.360 85.975 ;
        RECT 70.260 85.805 70.430 86.565 ;
        RECT 70.630 86.475 71.290 86.955 ;
        RECT 71.470 86.360 71.790 86.690 ;
        RECT 70.620 86.035 71.280 86.305 ;
        RECT 70.620 85.975 70.950 86.035 ;
        RECT 71.100 85.805 71.430 85.865 ;
        RECT 69.530 85.635 71.430 85.805 ;
        RECT 68.840 85.075 69.360 85.385 ;
        RECT 69.530 85.125 69.700 85.635 ;
        RECT 71.600 85.465 71.790 86.360 ;
        RECT 69.870 85.295 71.790 85.465 ;
        RECT 71.470 85.275 71.790 85.295 ;
        RECT 71.990 86.045 72.240 86.695 ;
        RECT 72.420 86.495 72.705 86.955 ;
        RECT 72.885 86.275 73.140 86.775 ;
        RECT 72.885 86.245 73.225 86.275 ;
        RECT 72.960 86.105 73.225 86.245 ;
        RECT 73.690 86.215 73.945 86.785 ;
        RECT 74.115 86.555 74.445 86.955 ;
        RECT 74.870 86.420 75.400 86.785 ;
        RECT 74.870 86.385 75.045 86.420 ;
        RECT 74.115 86.215 75.045 86.385 ;
        RECT 71.990 85.715 72.790 86.045 ;
        RECT 69.530 84.955 70.740 85.125 ;
        RECT 66.300 84.620 67.130 84.790 ;
        RECT 67.370 84.405 67.750 84.785 ;
        RECT 67.930 84.665 68.100 84.955 ;
        RECT 69.530 84.875 69.700 84.955 ;
        RECT 68.270 84.405 68.600 84.785 ;
        RECT 69.070 84.625 69.700 84.875 ;
        RECT 69.880 84.405 70.300 84.785 ;
        RECT 70.500 84.665 70.740 84.955 ;
        RECT 70.970 84.405 71.300 85.095 ;
        RECT 71.470 84.665 71.640 85.275 ;
        RECT 71.990 85.125 72.240 85.715 ;
        RECT 72.960 85.385 73.140 86.105 ;
        RECT 71.910 84.615 72.240 85.125 ;
        RECT 72.420 84.405 72.705 85.205 ;
        RECT 72.885 84.715 73.140 85.385 ;
        RECT 73.690 85.545 73.860 86.215 ;
        RECT 74.115 86.045 74.285 86.215 ;
        RECT 74.030 85.715 74.285 86.045 ;
        RECT 74.510 85.715 74.705 86.045 ;
        RECT 73.690 84.575 74.025 85.545 ;
        RECT 74.195 84.405 74.365 85.545 ;
        RECT 74.535 84.745 74.705 85.715 ;
        RECT 74.875 85.085 75.045 86.215 ;
        RECT 75.215 85.425 75.385 86.225 ;
        RECT 75.590 85.935 75.865 86.785 ;
        RECT 75.585 85.765 75.865 85.935 ;
        RECT 75.590 85.625 75.865 85.765 ;
        RECT 76.035 85.425 76.225 86.785 ;
        RECT 76.405 86.420 76.915 86.955 ;
        RECT 77.135 86.145 77.380 86.750 ;
        RECT 77.825 86.155 78.165 86.785 ;
        RECT 78.335 86.155 78.585 86.955 ;
        RECT 78.775 86.305 79.105 86.785 ;
        RECT 79.275 86.495 79.500 86.955 ;
        RECT 79.670 86.305 80.000 86.785 ;
        RECT 76.425 85.975 77.655 86.145 ;
        RECT 75.215 85.255 76.225 85.425 ;
        RECT 76.395 85.410 77.145 85.600 ;
        RECT 74.875 84.915 76.000 85.085 ;
        RECT 76.395 84.745 76.565 85.410 ;
        RECT 77.315 85.165 77.655 85.975 ;
        RECT 74.535 84.575 76.565 84.745 ;
        RECT 76.735 84.405 76.905 85.165 ;
        RECT 77.140 84.755 77.655 85.165 ;
        RECT 77.825 85.545 78.000 86.155 ;
        RECT 78.775 86.135 80.000 86.305 ;
        RECT 80.630 86.175 81.130 86.785 ;
        RECT 81.505 86.205 82.715 86.955 ;
        RECT 82.885 86.230 83.175 86.955 ;
        RECT 83.345 86.410 88.690 86.955 ;
        RECT 88.865 86.410 94.210 86.955 ;
        RECT 94.385 86.410 99.730 86.955 ;
        RECT 99.905 86.410 105.250 86.955 ;
        RECT 78.170 85.795 78.865 85.965 ;
        RECT 78.695 85.545 78.865 85.795 ;
        RECT 79.040 85.765 79.460 85.965 ;
        RECT 79.630 85.765 79.960 85.965 ;
        RECT 80.130 85.765 80.460 85.965 ;
        RECT 80.630 85.545 80.800 86.175 ;
        RECT 80.985 85.715 81.335 85.965 ;
        RECT 81.505 85.665 82.025 86.205 ;
        RECT 77.825 84.575 78.165 85.545 ;
        RECT 78.335 84.405 78.505 85.545 ;
        RECT 78.695 85.375 81.130 85.545 ;
        RECT 82.195 85.495 82.715 86.035 ;
        RECT 84.930 85.580 85.270 86.410 ;
        RECT 78.775 84.405 79.025 85.205 ;
        RECT 79.670 84.575 80.000 85.375 ;
        RECT 80.300 84.405 80.630 85.205 ;
        RECT 80.800 84.575 81.130 85.375 ;
        RECT 81.505 84.405 82.715 85.495 ;
        RECT 82.885 84.405 83.175 85.570 ;
        RECT 86.750 84.840 87.100 86.090 ;
        RECT 90.450 85.580 90.790 86.410 ;
        RECT 92.270 84.840 92.620 86.090 ;
        RECT 95.970 85.580 96.310 86.410 ;
        RECT 97.790 84.840 98.140 86.090 ;
        RECT 101.490 85.580 101.830 86.410 ;
        RECT 105.425 86.185 108.015 86.955 ;
        RECT 108.645 86.230 108.935 86.955 ;
        RECT 109.105 86.185 111.695 86.955 ;
        RECT 112.325 86.205 113.535 86.955 ;
        RECT 103.310 84.840 103.660 86.090 ;
        RECT 105.425 85.665 106.635 86.185 ;
        RECT 106.805 85.495 108.015 86.015 ;
        RECT 109.105 85.665 110.315 86.185 ;
        RECT 83.345 84.405 88.690 84.840 ;
        RECT 88.865 84.405 94.210 84.840 ;
        RECT 94.385 84.405 99.730 84.840 ;
        RECT 99.905 84.405 105.250 84.840 ;
        RECT 105.425 84.405 108.015 85.495 ;
        RECT 108.645 84.405 108.935 85.570 ;
        RECT 110.485 85.495 111.695 86.015 ;
        RECT 109.105 84.405 111.695 85.495 ;
        RECT 112.325 85.495 112.845 86.035 ;
        RECT 113.015 85.665 113.535 86.205 ;
        RECT 112.325 84.405 113.535 85.495 ;
        RECT 5.520 84.235 113.620 84.405 ;
        RECT 5.605 83.145 6.815 84.235 ;
        RECT 6.985 83.800 12.330 84.235 ;
        RECT 12.505 83.800 17.850 84.235 ;
        RECT 5.605 82.435 6.125 82.975 ;
        RECT 6.295 82.605 6.815 83.145 ;
        RECT 5.605 81.685 6.815 82.435 ;
        RECT 8.570 82.230 8.910 83.060 ;
        RECT 10.390 82.550 10.740 83.800 ;
        RECT 14.090 82.230 14.430 83.060 ;
        RECT 15.910 82.550 16.260 83.800 ;
        RECT 18.485 83.070 18.775 84.235 ;
        RECT 18.945 83.145 20.615 84.235 ;
        RECT 21.335 83.565 21.505 84.065 ;
        RECT 21.675 83.735 22.005 84.235 ;
        RECT 21.335 83.395 22.000 83.565 ;
        RECT 18.945 82.455 19.695 82.975 ;
        RECT 19.865 82.625 20.615 83.145 ;
        RECT 21.250 82.575 21.600 83.225 ;
        RECT 6.985 81.685 12.330 82.230 ;
        RECT 12.505 81.685 17.850 82.230 ;
        RECT 18.485 81.685 18.775 82.410 ;
        RECT 18.945 81.685 20.615 82.455 ;
        RECT 21.770 82.405 22.000 83.395 ;
        RECT 21.335 82.235 22.000 82.405 ;
        RECT 21.335 81.945 21.505 82.235 ;
        RECT 21.675 81.685 22.005 82.065 ;
        RECT 22.175 81.945 22.400 84.065 ;
        RECT 22.615 83.735 22.945 84.235 ;
        RECT 23.115 83.565 23.285 84.065 ;
        RECT 23.520 83.850 24.350 84.020 ;
        RECT 24.590 83.855 24.970 84.235 ;
        RECT 22.590 83.395 23.285 83.565 ;
        RECT 22.590 82.425 22.760 83.395 ;
        RECT 22.930 82.605 23.340 83.225 ;
        RECT 23.510 83.175 24.010 83.555 ;
        RECT 22.590 82.235 23.285 82.425 ;
        RECT 23.510 82.305 23.730 83.175 ;
        RECT 24.180 83.005 24.350 83.850 ;
        RECT 25.150 83.685 25.320 83.975 ;
        RECT 25.490 83.855 25.820 84.235 ;
        RECT 26.290 83.765 26.920 84.015 ;
        RECT 27.100 83.855 27.520 84.235 ;
        RECT 26.750 83.685 26.920 83.765 ;
        RECT 27.720 83.685 27.960 83.975 ;
        RECT 24.520 83.435 25.890 83.685 ;
        RECT 24.520 83.175 24.770 83.435 ;
        RECT 25.280 83.005 25.530 83.165 ;
        RECT 24.180 82.835 25.530 83.005 ;
        RECT 24.180 82.795 24.600 82.835 ;
        RECT 23.910 82.245 24.260 82.615 ;
        RECT 22.615 81.685 22.945 82.065 ;
        RECT 23.115 81.905 23.285 82.235 ;
        RECT 24.430 82.065 24.600 82.795 ;
        RECT 25.700 82.665 25.890 83.435 ;
        RECT 24.770 82.335 25.180 82.665 ;
        RECT 25.470 82.325 25.890 82.665 ;
        RECT 26.060 83.255 26.580 83.565 ;
        RECT 26.750 83.515 27.960 83.685 ;
        RECT 28.190 83.545 28.520 84.235 ;
        RECT 26.060 82.495 26.230 83.255 ;
        RECT 26.400 82.665 26.580 83.075 ;
        RECT 26.750 83.005 26.920 83.515 ;
        RECT 28.690 83.365 28.860 83.975 ;
        RECT 29.130 83.515 29.460 84.025 ;
        RECT 28.690 83.345 29.010 83.365 ;
        RECT 27.090 83.175 29.010 83.345 ;
        RECT 26.750 82.835 28.650 83.005 ;
        RECT 26.980 82.495 27.310 82.615 ;
        RECT 26.060 82.325 27.310 82.495 ;
        RECT 23.585 81.865 24.600 82.065 ;
        RECT 24.770 81.685 25.180 82.125 ;
        RECT 25.470 81.895 25.720 82.325 ;
        RECT 25.920 81.685 26.240 82.145 ;
        RECT 27.480 82.075 27.650 82.835 ;
        RECT 28.320 82.775 28.650 82.835 ;
        RECT 27.840 82.605 28.170 82.665 ;
        RECT 27.840 82.335 28.500 82.605 ;
        RECT 28.820 82.280 29.010 83.175 ;
        RECT 26.800 81.905 27.650 82.075 ;
        RECT 27.850 81.685 28.510 82.165 ;
        RECT 28.690 81.950 29.010 82.280 ;
        RECT 29.210 82.925 29.460 83.515 ;
        RECT 29.640 83.435 29.925 84.235 ;
        RECT 30.105 83.255 30.360 83.925 ;
        RECT 30.995 83.565 31.165 84.065 ;
        RECT 31.335 83.735 31.665 84.235 ;
        RECT 30.995 83.395 31.660 83.565 ;
        RECT 29.210 82.595 30.010 82.925 ;
        RECT 29.210 81.945 29.460 82.595 ;
        RECT 30.180 82.395 30.360 83.255 ;
        RECT 30.910 82.575 31.260 83.225 ;
        RECT 31.430 82.405 31.660 83.395 ;
        RECT 30.105 82.195 30.360 82.395 ;
        RECT 30.995 82.235 31.660 82.405 ;
        RECT 29.640 81.685 29.925 82.145 ;
        RECT 30.105 82.025 30.445 82.195 ;
        RECT 30.105 81.865 30.360 82.025 ;
        RECT 30.995 81.945 31.165 82.235 ;
        RECT 31.335 81.685 31.665 82.065 ;
        RECT 31.835 81.945 32.060 84.065 ;
        RECT 32.275 83.735 32.605 84.235 ;
        RECT 32.775 83.565 32.945 84.065 ;
        RECT 33.180 83.850 34.010 84.020 ;
        RECT 34.250 83.855 34.630 84.235 ;
        RECT 32.250 83.395 32.945 83.565 ;
        RECT 32.250 82.425 32.420 83.395 ;
        RECT 32.590 82.605 33.000 83.225 ;
        RECT 33.170 83.175 33.670 83.555 ;
        RECT 32.250 82.235 32.945 82.425 ;
        RECT 33.170 82.305 33.390 83.175 ;
        RECT 33.840 83.005 34.010 83.850 ;
        RECT 34.810 83.685 34.980 83.975 ;
        RECT 35.150 83.855 35.480 84.235 ;
        RECT 35.950 83.765 36.580 84.015 ;
        RECT 36.760 83.855 37.180 84.235 ;
        RECT 36.410 83.685 36.580 83.765 ;
        RECT 37.380 83.685 37.620 83.975 ;
        RECT 34.180 83.435 35.550 83.685 ;
        RECT 34.180 83.175 34.430 83.435 ;
        RECT 34.940 83.005 35.190 83.165 ;
        RECT 33.840 82.835 35.190 83.005 ;
        RECT 33.840 82.795 34.260 82.835 ;
        RECT 33.570 82.245 33.920 82.615 ;
        RECT 32.275 81.685 32.605 82.065 ;
        RECT 32.775 81.905 32.945 82.235 ;
        RECT 34.090 82.065 34.260 82.795 ;
        RECT 35.360 82.665 35.550 83.435 ;
        RECT 34.430 82.335 34.840 82.665 ;
        RECT 35.130 82.325 35.550 82.665 ;
        RECT 35.720 83.255 36.240 83.565 ;
        RECT 36.410 83.515 37.620 83.685 ;
        RECT 37.850 83.545 38.180 84.235 ;
        RECT 35.720 82.495 35.890 83.255 ;
        RECT 36.060 82.665 36.240 83.075 ;
        RECT 36.410 83.005 36.580 83.515 ;
        RECT 38.350 83.365 38.520 83.975 ;
        RECT 38.790 83.515 39.120 84.025 ;
        RECT 38.350 83.345 38.670 83.365 ;
        RECT 36.750 83.175 38.670 83.345 ;
        RECT 36.410 82.835 38.310 83.005 ;
        RECT 36.640 82.495 36.970 82.615 ;
        RECT 35.720 82.325 36.970 82.495 ;
        RECT 33.245 81.865 34.260 82.065 ;
        RECT 34.430 81.685 34.840 82.125 ;
        RECT 35.130 81.895 35.380 82.325 ;
        RECT 35.580 81.685 35.900 82.145 ;
        RECT 37.140 82.075 37.310 82.835 ;
        RECT 37.980 82.775 38.310 82.835 ;
        RECT 37.500 82.605 37.830 82.665 ;
        RECT 37.500 82.335 38.160 82.605 ;
        RECT 38.480 82.280 38.670 83.175 ;
        RECT 36.460 81.905 37.310 82.075 ;
        RECT 37.510 81.685 38.170 82.165 ;
        RECT 38.350 81.950 38.670 82.280 ;
        RECT 38.870 82.925 39.120 83.515 ;
        RECT 39.300 83.435 39.585 84.235 ;
        RECT 39.765 83.895 40.020 83.925 ;
        RECT 39.765 83.725 40.105 83.895 ;
        RECT 39.765 83.255 40.020 83.725 ;
        RECT 38.870 82.595 39.670 82.925 ;
        RECT 38.870 81.945 39.120 82.595 ;
        RECT 39.840 82.395 40.020 83.255 ;
        RECT 41.065 83.095 41.295 84.235 ;
        RECT 41.465 83.085 41.795 84.065 ;
        RECT 41.965 83.095 42.175 84.235 ;
        RECT 42.405 83.145 44.075 84.235 ;
        RECT 41.045 82.675 41.375 82.925 ;
        RECT 39.300 81.685 39.585 82.145 ;
        RECT 39.765 81.865 40.020 82.395 ;
        RECT 41.065 81.685 41.295 82.505 ;
        RECT 41.545 82.485 41.795 83.085 ;
        RECT 41.465 81.855 41.795 82.485 ;
        RECT 41.965 81.685 42.175 82.505 ;
        RECT 42.405 82.455 43.155 82.975 ;
        RECT 43.325 82.625 44.075 83.145 ;
        RECT 44.245 83.070 44.535 84.235 ;
        RECT 44.705 83.145 46.375 84.235 ;
        RECT 44.705 82.455 45.455 82.975 ;
        RECT 45.625 82.625 46.375 83.145 ;
        RECT 47.005 83.095 47.345 84.065 ;
        RECT 47.515 83.095 47.685 84.235 ;
        RECT 47.955 83.435 48.205 84.235 ;
        RECT 48.850 83.265 49.180 84.065 ;
        RECT 49.480 83.435 49.810 84.235 ;
        RECT 49.980 83.265 50.310 84.065 ;
        RECT 50.685 83.800 56.030 84.235 ;
        RECT 47.875 83.095 50.310 83.265 ;
        RECT 47.005 82.485 47.180 83.095 ;
        RECT 47.875 82.845 48.045 83.095 ;
        RECT 47.350 82.675 48.045 82.845 ;
        RECT 48.220 82.675 48.640 82.875 ;
        RECT 48.810 82.675 49.140 82.875 ;
        RECT 49.310 82.675 49.640 82.875 ;
        RECT 42.405 81.685 44.075 82.455 ;
        RECT 44.245 81.685 44.535 82.410 ;
        RECT 44.705 81.685 46.375 82.455 ;
        RECT 47.005 81.855 47.345 82.485 ;
        RECT 47.515 81.685 47.765 82.485 ;
        RECT 47.955 82.335 49.180 82.505 ;
        RECT 47.955 81.855 48.285 82.335 ;
        RECT 48.455 81.685 48.680 82.145 ;
        RECT 48.850 81.855 49.180 82.335 ;
        RECT 49.810 82.465 49.980 83.095 ;
        RECT 50.165 82.675 50.515 82.925 ;
        RECT 49.810 81.855 50.310 82.465 ;
        RECT 52.270 82.230 52.610 83.060 ;
        RECT 54.090 82.550 54.440 83.800 ;
        RECT 56.205 83.145 59.715 84.235 ;
        RECT 59.890 83.810 60.225 84.235 ;
        RECT 60.395 83.630 60.580 84.035 ;
        RECT 56.205 82.455 57.855 82.975 ;
        RECT 58.025 82.625 59.715 83.145 ;
        RECT 59.915 83.455 60.580 83.630 ;
        RECT 60.785 83.455 61.115 84.235 ;
        RECT 50.685 81.685 56.030 82.230 ;
        RECT 56.205 81.685 59.715 82.455 ;
        RECT 59.915 82.425 60.255 83.455 ;
        RECT 61.285 83.265 61.555 84.035 ;
        RECT 61.725 83.800 67.070 84.235 ;
        RECT 60.425 83.095 61.555 83.265 ;
        RECT 60.425 82.595 60.675 83.095 ;
        RECT 59.915 82.255 60.600 82.425 ;
        RECT 60.855 82.345 61.215 82.925 ;
        RECT 59.890 81.685 60.225 82.085 ;
        RECT 60.395 81.855 60.600 82.255 ;
        RECT 61.385 82.185 61.555 83.095 ;
        RECT 63.310 82.230 63.650 83.060 ;
        RECT 65.130 82.550 65.480 83.800 ;
        RECT 67.245 83.145 69.835 84.235 ;
        RECT 67.245 82.455 68.455 82.975 ;
        RECT 68.625 82.625 69.835 83.145 ;
        RECT 70.005 83.070 70.295 84.235 ;
        RECT 70.525 83.095 70.735 84.235 ;
        RECT 70.905 83.085 71.235 84.065 ;
        RECT 71.405 83.095 71.635 84.235 ;
        RECT 72.395 83.305 72.565 84.065 ;
        RECT 72.745 83.475 73.075 84.235 ;
        RECT 72.395 83.135 73.060 83.305 ;
        RECT 73.245 83.160 73.515 84.065 ;
        RECT 73.775 83.565 73.945 84.065 ;
        RECT 74.115 83.735 74.445 84.235 ;
        RECT 73.775 83.395 74.440 83.565 ;
        RECT 60.810 81.685 61.085 82.165 ;
        RECT 61.295 81.855 61.555 82.185 ;
        RECT 61.725 81.685 67.070 82.230 ;
        RECT 67.245 81.685 69.835 82.455 ;
        RECT 70.005 81.685 70.295 82.410 ;
        RECT 70.525 81.685 70.735 82.505 ;
        RECT 70.905 82.485 71.155 83.085 ;
        RECT 72.890 82.990 73.060 83.135 ;
        RECT 71.325 82.675 71.655 82.925 ;
        RECT 72.325 82.585 72.655 82.955 ;
        RECT 72.890 82.660 73.175 82.990 ;
        RECT 70.905 81.855 71.235 82.485 ;
        RECT 71.405 81.685 71.635 82.505 ;
        RECT 72.890 82.405 73.060 82.660 ;
        RECT 72.395 82.235 73.060 82.405 ;
        RECT 73.345 82.360 73.515 83.160 ;
        RECT 73.690 82.575 74.040 83.225 ;
        RECT 74.210 82.405 74.440 83.395 ;
        RECT 72.395 81.855 72.565 82.235 ;
        RECT 72.745 81.685 73.075 82.065 ;
        RECT 73.255 81.855 73.515 82.360 ;
        RECT 73.775 82.235 74.440 82.405 ;
        RECT 73.775 81.945 73.945 82.235 ;
        RECT 74.115 81.685 74.445 82.065 ;
        RECT 74.615 81.945 74.840 84.065 ;
        RECT 75.055 83.735 75.385 84.235 ;
        RECT 75.555 83.565 75.725 84.065 ;
        RECT 75.960 83.850 76.790 84.020 ;
        RECT 77.030 83.855 77.410 84.235 ;
        RECT 75.030 83.395 75.725 83.565 ;
        RECT 75.030 82.425 75.200 83.395 ;
        RECT 75.370 82.605 75.780 83.225 ;
        RECT 75.950 83.175 76.450 83.555 ;
        RECT 75.030 82.235 75.725 82.425 ;
        RECT 75.950 82.305 76.170 83.175 ;
        RECT 76.620 83.005 76.790 83.850 ;
        RECT 77.590 83.685 77.760 83.975 ;
        RECT 77.930 83.855 78.260 84.235 ;
        RECT 78.730 83.765 79.360 84.015 ;
        RECT 79.540 83.855 79.960 84.235 ;
        RECT 79.190 83.685 79.360 83.765 ;
        RECT 80.160 83.685 80.400 83.975 ;
        RECT 76.960 83.435 78.330 83.685 ;
        RECT 76.960 83.175 77.210 83.435 ;
        RECT 77.720 83.005 77.970 83.165 ;
        RECT 76.620 82.835 77.970 83.005 ;
        RECT 76.620 82.795 77.040 82.835 ;
        RECT 76.350 82.245 76.700 82.615 ;
        RECT 75.055 81.685 75.385 82.065 ;
        RECT 75.555 81.905 75.725 82.235 ;
        RECT 76.870 82.065 77.040 82.795 ;
        RECT 78.140 82.665 78.330 83.435 ;
        RECT 77.210 82.335 77.620 82.665 ;
        RECT 77.910 82.325 78.330 82.665 ;
        RECT 78.500 83.255 79.020 83.565 ;
        RECT 79.190 83.515 80.400 83.685 ;
        RECT 80.630 83.545 80.960 84.235 ;
        RECT 78.500 82.495 78.670 83.255 ;
        RECT 78.840 82.665 79.020 83.075 ;
        RECT 79.190 83.005 79.360 83.515 ;
        RECT 81.130 83.365 81.300 83.975 ;
        RECT 81.570 83.515 81.900 84.025 ;
        RECT 81.130 83.345 81.450 83.365 ;
        RECT 79.530 83.175 81.450 83.345 ;
        RECT 79.190 82.835 81.090 83.005 ;
        RECT 79.420 82.495 79.750 82.615 ;
        RECT 78.500 82.325 79.750 82.495 ;
        RECT 76.025 81.865 77.040 82.065 ;
        RECT 77.210 81.685 77.620 82.125 ;
        RECT 77.910 81.895 78.160 82.325 ;
        RECT 78.360 81.685 78.680 82.145 ;
        RECT 79.920 82.075 80.090 82.835 ;
        RECT 80.760 82.775 81.090 82.835 ;
        RECT 80.280 82.605 80.610 82.665 ;
        RECT 80.280 82.335 80.940 82.605 ;
        RECT 81.260 82.280 81.450 83.175 ;
        RECT 79.240 81.905 80.090 82.075 ;
        RECT 80.290 81.685 80.950 82.165 ;
        RECT 81.130 81.950 81.450 82.280 ;
        RECT 81.650 82.925 81.900 83.515 ;
        RECT 82.080 83.435 82.365 84.235 ;
        RECT 82.545 83.895 82.800 83.925 ;
        RECT 82.545 83.725 82.885 83.895 ;
        RECT 83.345 83.800 88.690 84.235 ;
        RECT 82.545 83.255 82.800 83.725 ;
        RECT 81.650 82.595 82.450 82.925 ;
        RECT 81.650 81.945 81.900 82.595 ;
        RECT 82.620 82.395 82.800 83.255 ;
        RECT 82.080 81.685 82.365 82.145 ;
        RECT 82.545 81.865 82.800 82.395 ;
        RECT 84.930 82.230 85.270 83.060 ;
        RECT 86.750 82.550 87.100 83.800 ;
        RECT 88.865 83.145 92.375 84.235 ;
        RECT 93.205 83.565 93.485 84.235 ;
        RECT 93.655 83.345 93.955 83.895 ;
        RECT 94.155 83.515 94.485 84.235 ;
        RECT 94.675 83.515 95.135 84.065 ;
        RECT 88.865 82.455 90.515 82.975 ;
        RECT 90.685 82.625 92.375 83.145 ;
        RECT 93.020 82.925 93.285 83.285 ;
        RECT 93.655 83.175 94.595 83.345 ;
        RECT 94.425 82.925 94.595 83.175 ;
        RECT 93.020 82.675 93.695 82.925 ;
        RECT 93.915 82.675 94.255 82.925 ;
        RECT 94.425 82.595 94.715 82.925 ;
        RECT 94.425 82.505 94.595 82.595 ;
        RECT 83.345 81.685 88.690 82.230 ;
        RECT 88.865 81.685 92.375 82.455 ;
        RECT 93.205 82.315 94.595 82.505 ;
        RECT 93.205 81.955 93.535 82.315 ;
        RECT 94.885 82.145 95.135 83.515 ;
        RECT 95.765 83.070 96.055 84.235 ;
        RECT 96.285 83.095 96.495 84.235 ;
        RECT 96.665 83.085 96.995 84.065 ;
        RECT 97.165 83.095 97.395 84.235 ;
        RECT 97.605 83.145 101.115 84.235 ;
        RECT 102.295 83.565 102.465 84.065 ;
        RECT 102.635 83.735 102.965 84.235 ;
        RECT 102.295 83.395 102.960 83.565 ;
        RECT 94.155 81.685 94.405 82.145 ;
        RECT 94.575 81.855 95.135 82.145 ;
        RECT 95.765 81.685 96.055 82.410 ;
        RECT 96.285 81.685 96.495 82.505 ;
        RECT 96.665 82.485 96.915 83.085 ;
        RECT 97.085 82.675 97.415 82.925 ;
        RECT 96.665 81.855 96.995 82.485 ;
        RECT 97.165 81.685 97.395 82.505 ;
        RECT 97.605 82.455 99.255 82.975 ;
        RECT 99.425 82.625 101.115 83.145 ;
        RECT 102.210 82.575 102.560 83.225 ;
        RECT 97.605 81.685 101.115 82.455 ;
        RECT 102.730 82.405 102.960 83.395 ;
        RECT 102.295 82.235 102.960 82.405 ;
        RECT 102.295 81.945 102.465 82.235 ;
        RECT 102.635 81.685 102.965 82.065 ;
        RECT 103.135 81.945 103.360 84.065 ;
        RECT 103.575 83.735 103.905 84.235 ;
        RECT 104.075 83.565 104.245 84.065 ;
        RECT 104.480 83.850 105.310 84.020 ;
        RECT 105.550 83.855 105.930 84.235 ;
        RECT 103.550 83.395 104.245 83.565 ;
        RECT 103.550 82.425 103.720 83.395 ;
        RECT 103.890 82.605 104.300 83.225 ;
        RECT 104.470 83.175 104.970 83.555 ;
        RECT 103.550 82.235 104.245 82.425 ;
        RECT 104.470 82.305 104.690 83.175 ;
        RECT 105.140 83.005 105.310 83.850 ;
        RECT 106.110 83.685 106.280 83.975 ;
        RECT 106.450 83.855 106.780 84.235 ;
        RECT 107.250 83.765 107.880 84.015 ;
        RECT 108.060 83.855 108.480 84.235 ;
        RECT 107.710 83.685 107.880 83.765 ;
        RECT 108.680 83.685 108.920 83.975 ;
        RECT 105.480 83.435 106.850 83.685 ;
        RECT 105.480 83.175 105.730 83.435 ;
        RECT 106.240 83.005 106.490 83.165 ;
        RECT 105.140 82.835 106.490 83.005 ;
        RECT 105.140 82.795 105.560 82.835 ;
        RECT 104.870 82.245 105.220 82.615 ;
        RECT 103.575 81.685 103.905 82.065 ;
        RECT 104.075 81.905 104.245 82.235 ;
        RECT 105.390 82.065 105.560 82.795 ;
        RECT 106.660 82.665 106.850 83.435 ;
        RECT 105.730 82.335 106.140 82.665 ;
        RECT 106.430 82.325 106.850 82.665 ;
        RECT 107.020 83.255 107.540 83.565 ;
        RECT 107.710 83.515 108.920 83.685 ;
        RECT 109.150 83.545 109.480 84.235 ;
        RECT 107.020 82.495 107.190 83.255 ;
        RECT 107.360 82.665 107.540 83.075 ;
        RECT 107.710 83.005 107.880 83.515 ;
        RECT 109.650 83.365 109.820 83.975 ;
        RECT 110.090 83.515 110.420 84.025 ;
        RECT 109.650 83.345 109.970 83.365 ;
        RECT 108.050 83.175 109.970 83.345 ;
        RECT 107.710 82.835 109.610 83.005 ;
        RECT 107.940 82.495 108.270 82.615 ;
        RECT 107.020 82.325 108.270 82.495 ;
        RECT 104.545 81.865 105.560 82.065 ;
        RECT 105.730 81.685 106.140 82.125 ;
        RECT 106.430 81.895 106.680 82.325 ;
        RECT 106.880 81.685 107.200 82.145 ;
        RECT 108.440 82.075 108.610 82.835 ;
        RECT 109.280 82.775 109.610 82.835 ;
        RECT 108.800 82.605 109.130 82.665 ;
        RECT 108.800 82.335 109.460 82.605 ;
        RECT 109.780 82.280 109.970 83.175 ;
        RECT 107.760 81.905 108.610 82.075 ;
        RECT 108.810 81.685 109.470 82.165 ;
        RECT 109.650 81.950 109.970 82.280 ;
        RECT 110.170 82.925 110.420 83.515 ;
        RECT 110.600 83.435 110.885 84.235 ;
        RECT 111.065 83.895 111.320 83.925 ;
        RECT 111.065 83.725 111.405 83.895 ;
        RECT 111.065 83.255 111.320 83.725 ;
        RECT 110.170 82.595 110.970 82.925 ;
        RECT 110.170 81.945 110.420 82.595 ;
        RECT 111.140 82.395 111.320 83.255 ;
        RECT 112.325 83.145 113.535 84.235 ;
        RECT 112.325 82.605 112.845 83.145 ;
        RECT 113.015 82.435 113.535 82.975 ;
        RECT 110.600 81.685 110.885 82.145 ;
        RECT 111.065 81.865 111.320 82.395 ;
        RECT 112.325 81.685 113.535 82.435 ;
        RECT 5.520 81.515 113.620 81.685 ;
        RECT 5.605 80.765 6.815 81.515 ;
        RECT 5.605 80.225 6.125 80.765 ;
        RECT 6.985 80.745 9.575 81.515 ;
        RECT 10.205 80.840 10.465 81.345 ;
        RECT 10.645 81.135 10.975 81.515 ;
        RECT 11.155 80.965 11.325 81.345 ;
        RECT 6.295 80.055 6.815 80.595 ;
        RECT 6.985 80.225 8.195 80.745 ;
        RECT 8.365 80.055 9.575 80.575 ;
        RECT 5.605 78.965 6.815 80.055 ;
        RECT 6.985 78.965 9.575 80.055 ;
        RECT 10.205 80.040 10.375 80.840 ;
        RECT 10.660 80.795 11.325 80.965 ;
        RECT 11.585 80.840 11.845 81.345 ;
        RECT 12.025 81.135 12.355 81.515 ;
        RECT 12.535 80.965 12.705 81.345 ;
        RECT 10.660 80.540 10.830 80.795 ;
        RECT 10.545 80.210 10.830 80.540 ;
        RECT 11.065 80.245 11.395 80.615 ;
        RECT 10.660 80.065 10.830 80.210 ;
        RECT 10.205 79.135 10.475 80.040 ;
        RECT 10.660 79.895 11.325 80.065 ;
        RECT 10.645 78.965 10.975 79.725 ;
        RECT 11.155 79.135 11.325 79.895 ;
        RECT 11.585 80.040 11.755 80.840 ;
        RECT 12.040 80.795 12.705 80.965 ;
        RECT 12.040 80.540 12.210 80.795 ;
        RECT 12.965 80.765 14.175 81.515 ;
        RECT 14.350 80.775 14.605 81.345 ;
        RECT 14.775 81.115 15.105 81.515 ;
        RECT 15.530 80.980 16.060 81.345 ;
        RECT 15.530 80.945 15.705 80.980 ;
        RECT 14.775 80.775 15.705 80.945 ;
        RECT 11.925 80.210 12.210 80.540 ;
        RECT 12.445 80.245 12.775 80.615 ;
        RECT 12.965 80.225 13.485 80.765 ;
        RECT 12.040 80.065 12.210 80.210 ;
        RECT 11.585 79.135 11.855 80.040 ;
        RECT 12.040 79.895 12.705 80.065 ;
        RECT 13.655 80.055 14.175 80.595 ;
        RECT 12.025 78.965 12.355 79.725 ;
        RECT 12.535 79.135 12.705 79.895 ;
        RECT 12.965 78.965 14.175 80.055 ;
        RECT 14.350 80.105 14.520 80.775 ;
        RECT 14.775 80.605 14.945 80.775 ;
        RECT 14.690 80.275 14.945 80.605 ;
        RECT 15.170 80.275 15.365 80.605 ;
        RECT 14.350 79.135 14.685 80.105 ;
        RECT 14.855 78.965 15.025 80.105 ;
        RECT 15.195 79.305 15.365 80.275 ;
        RECT 15.535 79.645 15.705 80.775 ;
        RECT 15.875 79.985 16.045 80.785 ;
        RECT 16.250 80.495 16.525 81.345 ;
        RECT 16.245 80.325 16.525 80.495 ;
        RECT 16.250 80.185 16.525 80.325 ;
        RECT 16.695 79.985 16.885 81.345 ;
        RECT 17.065 80.980 17.575 81.515 ;
        RECT 17.795 80.705 18.040 81.310 ;
        RECT 18.485 80.745 21.995 81.515 ;
        RECT 23.085 80.840 23.345 81.345 ;
        RECT 23.525 81.135 23.855 81.515 ;
        RECT 24.035 80.965 24.205 81.345 ;
        RECT 17.085 80.535 18.315 80.705 ;
        RECT 15.875 79.815 16.885 79.985 ;
        RECT 17.055 79.970 17.805 80.160 ;
        RECT 15.535 79.475 16.660 79.645 ;
        RECT 17.055 79.305 17.225 79.970 ;
        RECT 17.975 79.725 18.315 80.535 ;
        RECT 18.485 80.225 20.135 80.745 ;
        RECT 20.305 80.055 21.995 80.575 ;
        RECT 15.195 79.135 17.225 79.305 ;
        RECT 17.395 78.965 17.565 79.725 ;
        RECT 17.800 79.315 18.315 79.725 ;
        RECT 18.485 78.965 21.995 80.055 ;
        RECT 23.085 80.040 23.255 80.840 ;
        RECT 23.540 80.795 24.205 80.965 ;
        RECT 23.540 80.540 23.710 80.795 ;
        RECT 24.470 80.775 24.725 81.345 ;
        RECT 24.895 81.115 25.225 81.515 ;
        RECT 25.650 80.980 26.180 81.345 ;
        RECT 25.650 80.945 25.825 80.980 ;
        RECT 24.895 80.775 25.825 80.945 ;
        RECT 23.425 80.210 23.710 80.540 ;
        RECT 23.945 80.245 24.275 80.615 ;
        RECT 23.540 80.065 23.710 80.210 ;
        RECT 24.470 80.105 24.640 80.775 ;
        RECT 24.895 80.605 25.065 80.775 ;
        RECT 24.810 80.275 25.065 80.605 ;
        RECT 25.290 80.275 25.485 80.605 ;
        RECT 23.085 79.135 23.355 80.040 ;
        RECT 23.540 79.895 24.205 80.065 ;
        RECT 23.525 78.965 23.855 79.725 ;
        RECT 24.035 79.135 24.205 79.895 ;
        RECT 24.470 79.135 24.805 80.105 ;
        RECT 24.975 78.965 25.145 80.105 ;
        RECT 25.315 79.305 25.485 80.275 ;
        RECT 25.655 79.645 25.825 80.775 ;
        RECT 25.995 79.985 26.165 80.785 ;
        RECT 26.370 80.495 26.645 81.345 ;
        RECT 26.365 80.325 26.645 80.495 ;
        RECT 26.370 80.185 26.645 80.325 ;
        RECT 26.815 79.985 27.005 81.345 ;
        RECT 27.185 80.980 27.695 81.515 ;
        RECT 27.915 80.705 28.160 81.310 ;
        RECT 27.205 80.535 28.435 80.705 ;
        RECT 28.665 80.695 28.875 81.515 ;
        RECT 29.045 80.715 29.375 81.345 ;
        RECT 25.995 79.815 27.005 79.985 ;
        RECT 27.175 79.970 27.925 80.160 ;
        RECT 25.655 79.475 26.780 79.645 ;
        RECT 27.175 79.305 27.345 79.970 ;
        RECT 28.095 79.725 28.435 80.535 ;
        RECT 29.045 80.115 29.295 80.715 ;
        RECT 29.545 80.695 29.775 81.515 ;
        RECT 29.985 80.765 31.195 81.515 ;
        RECT 31.365 80.790 31.655 81.515 ;
        RECT 32.290 80.775 32.545 81.345 ;
        RECT 32.715 81.115 33.045 81.515 ;
        RECT 33.470 80.980 34.000 81.345 ;
        RECT 33.470 80.945 33.645 80.980 ;
        RECT 32.715 80.775 33.645 80.945 ;
        RECT 29.465 80.275 29.795 80.525 ;
        RECT 29.985 80.225 30.505 80.765 ;
        RECT 25.315 79.135 27.345 79.305 ;
        RECT 27.515 78.965 27.685 79.725 ;
        RECT 27.920 79.315 28.435 79.725 ;
        RECT 28.665 78.965 28.875 80.105 ;
        RECT 29.045 79.135 29.375 80.115 ;
        RECT 29.545 78.965 29.775 80.105 ;
        RECT 30.675 80.055 31.195 80.595 ;
        RECT 29.985 78.965 31.195 80.055 ;
        RECT 31.365 78.965 31.655 80.130 ;
        RECT 32.290 80.105 32.460 80.775 ;
        RECT 32.715 80.605 32.885 80.775 ;
        RECT 32.630 80.275 32.885 80.605 ;
        RECT 33.110 80.275 33.305 80.605 ;
        RECT 32.290 79.135 32.625 80.105 ;
        RECT 32.795 78.965 32.965 80.105 ;
        RECT 33.135 79.305 33.305 80.275 ;
        RECT 33.475 79.645 33.645 80.775 ;
        RECT 33.815 79.985 33.985 80.785 ;
        RECT 34.190 80.495 34.465 81.345 ;
        RECT 34.185 80.325 34.465 80.495 ;
        RECT 34.190 80.185 34.465 80.325 ;
        RECT 34.635 79.985 34.825 81.345 ;
        RECT 35.005 80.980 35.515 81.515 ;
        RECT 35.735 80.705 35.980 81.310 ;
        RECT 36.425 80.745 39.935 81.515 ;
        RECT 41.025 80.840 41.285 81.345 ;
        RECT 41.465 81.135 41.795 81.515 ;
        RECT 41.975 80.965 42.145 81.345 ;
        RECT 35.025 80.535 36.255 80.705 ;
        RECT 33.815 79.815 34.825 79.985 ;
        RECT 34.995 79.970 35.745 80.160 ;
        RECT 33.475 79.475 34.600 79.645 ;
        RECT 34.995 79.305 35.165 79.970 ;
        RECT 35.915 79.725 36.255 80.535 ;
        RECT 36.425 80.225 38.075 80.745 ;
        RECT 38.245 80.055 39.935 80.575 ;
        RECT 33.135 79.135 35.165 79.305 ;
        RECT 35.335 78.965 35.505 79.725 ;
        RECT 35.740 79.315 36.255 79.725 ;
        RECT 36.425 78.965 39.935 80.055 ;
        RECT 41.025 80.040 41.195 80.840 ;
        RECT 41.480 80.795 42.145 80.965 ;
        RECT 41.480 80.540 41.650 80.795 ;
        RECT 42.870 80.775 43.125 81.345 ;
        RECT 43.295 81.115 43.625 81.515 ;
        RECT 44.050 80.980 44.580 81.345 ;
        RECT 44.770 81.175 45.045 81.345 ;
        RECT 44.765 81.005 45.045 81.175 ;
        RECT 44.050 80.945 44.225 80.980 ;
        RECT 43.295 80.775 44.225 80.945 ;
        RECT 41.365 80.210 41.650 80.540 ;
        RECT 41.885 80.245 42.215 80.615 ;
        RECT 41.480 80.065 41.650 80.210 ;
        RECT 42.870 80.105 43.040 80.775 ;
        RECT 43.295 80.605 43.465 80.775 ;
        RECT 43.210 80.275 43.465 80.605 ;
        RECT 43.690 80.275 43.885 80.605 ;
        RECT 41.025 79.135 41.295 80.040 ;
        RECT 41.480 79.895 42.145 80.065 ;
        RECT 41.465 78.965 41.795 79.725 ;
        RECT 41.975 79.135 42.145 79.895 ;
        RECT 42.870 79.135 43.205 80.105 ;
        RECT 43.375 78.965 43.545 80.105 ;
        RECT 43.715 79.305 43.885 80.275 ;
        RECT 44.055 79.645 44.225 80.775 ;
        RECT 44.395 79.985 44.565 80.785 ;
        RECT 44.770 80.185 45.045 81.005 ;
        RECT 45.215 79.985 45.405 81.345 ;
        RECT 45.585 80.980 46.095 81.515 ;
        RECT 46.315 80.705 46.560 81.310 ;
        RECT 47.005 80.970 52.350 81.515 ;
        RECT 45.605 80.535 46.835 80.705 ;
        RECT 44.395 79.815 45.405 79.985 ;
        RECT 45.575 79.970 46.325 80.160 ;
        RECT 44.055 79.475 45.180 79.645 ;
        RECT 45.575 79.305 45.745 79.970 ;
        RECT 46.495 79.725 46.835 80.535 ;
        RECT 48.590 80.140 48.930 80.970 ;
        RECT 52.525 80.745 56.035 81.515 ;
        RECT 57.125 80.790 57.415 81.515 ;
        RECT 57.585 80.970 62.930 81.515 ;
        RECT 63.105 80.970 68.450 81.515 ;
        RECT 68.625 80.970 73.970 81.515 ;
        RECT 43.715 79.135 45.745 79.305 ;
        RECT 45.915 78.965 46.085 79.725 ;
        RECT 46.320 79.315 46.835 79.725 ;
        RECT 50.410 79.400 50.760 80.650 ;
        RECT 52.525 80.225 54.175 80.745 ;
        RECT 54.345 80.055 56.035 80.575 ;
        RECT 59.170 80.140 59.510 80.970 ;
        RECT 47.005 78.965 52.350 79.400 ;
        RECT 52.525 78.965 56.035 80.055 ;
        RECT 57.125 78.965 57.415 80.130 ;
        RECT 60.990 79.400 61.340 80.650 ;
        RECT 64.690 80.140 65.030 80.970 ;
        RECT 66.510 79.400 66.860 80.650 ;
        RECT 70.210 80.140 70.550 80.970 ;
        RECT 75.070 80.775 75.325 81.345 ;
        RECT 75.495 81.115 75.825 81.515 ;
        RECT 76.250 80.980 76.780 81.345 ;
        RECT 76.250 80.945 76.425 80.980 ;
        RECT 75.495 80.775 76.425 80.945 ;
        RECT 72.030 79.400 72.380 80.650 ;
        RECT 75.070 80.105 75.240 80.775 ;
        RECT 75.495 80.605 75.665 80.775 ;
        RECT 75.410 80.275 75.665 80.605 ;
        RECT 75.890 80.275 76.085 80.605 ;
        RECT 57.585 78.965 62.930 79.400 ;
        RECT 63.105 78.965 68.450 79.400 ;
        RECT 68.625 78.965 73.970 79.400 ;
        RECT 75.070 79.135 75.405 80.105 ;
        RECT 75.575 78.965 75.745 80.105 ;
        RECT 75.915 79.305 76.085 80.275 ;
        RECT 76.255 79.645 76.425 80.775 ;
        RECT 76.595 79.985 76.765 80.785 ;
        RECT 76.970 80.495 77.245 81.345 ;
        RECT 76.965 80.325 77.245 80.495 ;
        RECT 76.970 80.185 77.245 80.325 ;
        RECT 77.415 79.985 77.605 81.345 ;
        RECT 77.785 80.980 78.295 81.515 ;
        RECT 78.515 80.705 78.760 81.310 ;
        RECT 77.805 80.535 79.035 80.705 ;
        RECT 79.265 80.695 79.475 81.515 ;
        RECT 79.645 80.715 79.975 81.345 ;
        RECT 76.595 79.815 77.605 79.985 ;
        RECT 77.775 79.970 78.525 80.160 ;
        RECT 76.255 79.475 77.380 79.645 ;
        RECT 77.775 79.305 77.945 79.970 ;
        RECT 78.695 79.725 79.035 80.535 ;
        RECT 79.645 80.115 79.895 80.715 ;
        RECT 80.145 80.695 80.375 81.515 ;
        RECT 80.585 80.745 82.255 81.515 ;
        RECT 82.885 80.790 83.175 81.515 ;
        RECT 83.345 80.970 88.690 81.515 ;
        RECT 80.065 80.275 80.395 80.525 ;
        RECT 80.585 80.225 81.335 80.745 ;
        RECT 75.915 79.135 77.945 79.305 ;
        RECT 78.115 78.965 78.285 79.725 ;
        RECT 78.520 79.315 79.035 79.725 ;
        RECT 79.265 78.965 79.475 80.105 ;
        RECT 79.645 79.135 79.975 80.115 ;
        RECT 80.145 78.965 80.375 80.105 ;
        RECT 81.505 80.055 82.255 80.575 ;
        RECT 84.930 80.140 85.270 80.970 ;
        RECT 89.875 80.965 90.045 81.345 ;
        RECT 90.225 81.135 90.555 81.515 ;
        RECT 89.875 80.795 90.540 80.965 ;
        RECT 90.735 80.840 90.995 81.345 ;
        RECT 80.585 78.965 82.255 80.055 ;
        RECT 82.885 78.965 83.175 80.130 ;
        RECT 86.750 79.400 87.100 80.650 ;
        RECT 89.805 80.245 90.135 80.615 ;
        RECT 90.370 80.540 90.540 80.795 ;
        RECT 90.370 80.210 90.655 80.540 ;
        RECT 90.370 80.065 90.540 80.210 ;
        RECT 89.875 79.895 90.540 80.065 ;
        RECT 90.825 80.040 90.995 80.840 ;
        RECT 91.255 80.965 91.425 81.255 ;
        RECT 91.595 81.135 91.925 81.515 ;
        RECT 91.255 80.795 91.920 80.965 ;
        RECT 83.345 78.965 88.690 79.400 ;
        RECT 89.875 79.135 90.045 79.895 ;
        RECT 90.225 78.965 90.555 79.725 ;
        RECT 90.725 79.135 90.995 80.040 ;
        RECT 91.170 79.975 91.520 80.625 ;
        RECT 91.690 79.805 91.920 80.795 ;
        RECT 91.255 79.635 91.920 79.805 ;
        RECT 91.255 79.135 91.425 79.635 ;
        RECT 91.595 78.965 91.925 79.465 ;
        RECT 92.095 79.135 92.320 81.255 ;
        RECT 92.535 81.135 92.865 81.515 ;
        RECT 93.035 80.965 93.205 81.295 ;
        RECT 93.505 81.135 94.520 81.335 ;
        RECT 92.510 80.775 93.205 80.965 ;
        RECT 92.510 79.805 92.680 80.775 ;
        RECT 92.850 79.975 93.260 80.595 ;
        RECT 93.430 80.025 93.650 80.895 ;
        RECT 93.830 80.585 94.180 80.955 ;
        RECT 94.350 80.405 94.520 81.135 ;
        RECT 94.690 81.075 95.100 81.515 ;
        RECT 95.390 80.875 95.640 81.305 ;
        RECT 95.840 81.055 96.160 81.515 ;
        RECT 96.720 81.125 97.570 81.295 ;
        RECT 94.690 80.535 95.100 80.865 ;
        RECT 95.390 80.535 95.810 80.875 ;
        RECT 94.100 80.365 94.520 80.405 ;
        RECT 94.100 80.195 95.450 80.365 ;
        RECT 92.510 79.635 93.205 79.805 ;
        RECT 93.430 79.645 93.930 80.025 ;
        RECT 92.535 78.965 92.865 79.465 ;
        RECT 93.035 79.135 93.205 79.635 ;
        RECT 94.100 79.350 94.270 80.195 ;
        RECT 95.200 80.035 95.450 80.195 ;
        RECT 94.440 79.765 94.690 80.025 ;
        RECT 95.620 79.765 95.810 80.535 ;
        RECT 94.440 79.515 95.810 79.765 ;
        RECT 95.980 80.705 97.230 80.875 ;
        RECT 95.980 79.945 96.150 80.705 ;
        RECT 96.900 80.585 97.230 80.705 ;
        RECT 96.320 80.125 96.500 80.535 ;
        RECT 97.400 80.365 97.570 81.125 ;
        RECT 97.770 81.035 98.430 81.515 ;
        RECT 98.610 80.920 98.930 81.250 ;
        RECT 97.760 80.595 98.420 80.865 ;
        RECT 97.760 80.535 98.090 80.595 ;
        RECT 98.240 80.365 98.570 80.425 ;
        RECT 96.670 80.195 98.570 80.365 ;
        RECT 95.980 79.635 96.500 79.945 ;
        RECT 96.670 79.685 96.840 80.195 ;
        RECT 98.740 80.025 98.930 80.920 ;
        RECT 97.010 79.855 98.930 80.025 ;
        RECT 98.610 79.835 98.930 79.855 ;
        RECT 99.130 80.605 99.380 81.255 ;
        RECT 99.560 81.055 99.845 81.515 ;
        RECT 100.025 80.805 100.280 81.335 ;
        RECT 99.130 80.275 99.930 80.605 ;
        RECT 96.670 79.515 97.880 79.685 ;
        RECT 93.440 79.180 94.270 79.350 ;
        RECT 94.510 78.965 94.890 79.345 ;
        RECT 95.070 79.225 95.240 79.515 ;
        RECT 96.670 79.435 96.840 79.515 ;
        RECT 95.410 78.965 95.740 79.345 ;
        RECT 96.210 79.185 96.840 79.435 ;
        RECT 97.020 78.965 97.440 79.345 ;
        RECT 97.640 79.225 97.880 79.515 ;
        RECT 98.110 78.965 98.440 79.655 ;
        RECT 98.610 79.225 98.780 79.835 ;
        RECT 99.130 79.685 99.380 80.275 ;
        RECT 100.100 79.945 100.280 80.805 ;
        RECT 101.100 80.705 101.345 81.310 ;
        RECT 101.565 80.980 102.075 81.515 ;
        RECT 99.050 79.175 99.380 79.685 ;
        RECT 99.560 78.965 99.845 79.765 ;
        RECT 100.025 79.475 100.280 79.945 ;
        RECT 100.825 80.535 102.055 80.705 ;
        RECT 100.825 79.725 101.165 80.535 ;
        RECT 101.335 79.970 102.085 80.160 ;
        RECT 100.025 79.305 100.365 79.475 ;
        RECT 100.825 79.315 101.340 79.725 ;
        RECT 100.025 79.275 100.280 79.305 ;
        RECT 101.575 78.965 101.745 79.725 ;
        RECT 101.915 79.305 102.085 79.970 ;
        RECT 102.255 79.985 102.445 81.345 ;
        RECT 102.615 80.495 102.890 81.345 ;
        RECT 103.080 80.980 103.610 81.345 ;
        RECT 104.035 81.115 104.365 81.515 ;
        RECT 103.435 80.945 103.610 80.980 ;
        RECT 102.615 80.325 102.895 80.495 ;
        RECT 102.615 80.185 102.890 80.325 ;
        RECT 103.095 79.985 103.265 80.785 ;
        RECT 102.255 79.815 103.265 79.985 ;
        RECT 103.435 80.775 104.365 80.945 ;
        RECT 104.535 80.775 104.790 81.345 ;
        RECT 103.435 79.645 103.605 80.775 ;
        RECT 104.195 80.605 104.365 80.775 ;
        RECT 102.480 79.475 103.605 79.645 ;
        RECT 103.775 80.275 103.970 80.605 ;
        RECT 104.195 80.275 104.450 80.605 ;
        RECT 103.775 79.305 103.945 80.275 ;
        RECT 104.620 80.105 104.790 80.775 ;
        RECT 101.915 79.135 103.945 79.305 ;
        RECT 104.115 78.965 104.285 80.105 ;
        RECT 104.455 79.135 104.790 80.105 ;
        RECT 104.965 80.840 105.225 81.345 ;
        RECT 105.405 81.135 105.735 81.515 ;
        RECT 105.915 80.965 106.085 81.345 ;
        RECT 104.965 80.040 105.135 80.840 ;
        RECT 105.420 80.795 106.085 80.965 ;
        RECT 106.345 80.840 106.605 81.345 ;
        RECT 106.785 81.135 107.115 81.515 ;
        RECT 107.295 80.965 107.465 81.345 ;
        RECT 105.420 80.540 105.590 80.795 ;
        RECT 105.305 80.210 105.590 80.540 ;
        RECT 105.825 80.245 106.155 80.615 ;
        RECT 105.420 80.065 105.590 80.210 ;
        RECT 104.965 79.135 105.235 80.040 ;
        RECT 105.420 79.895 106.085 80.065 ;
        RECT 105.405 78.965 105.735 79.725 ;
        RECT 105.915 79.135 106.085 79.895 ;
        RECT 106.345 80.040 106.515 80.840 ;
        RECT 106.800 80.795 107.465 80.965 ;
        RECT 106.800 80.540 106.970 80.795 ;
        RECT 108.645 80.790 108.935 81.515 ;
        RECT 109.165 80.695 109.375 81.515 ;
        RECT 109.545 80.715 109.875 81.345 ;
        RECT 106.685 80.210 106.970 80.540 ;
        RECT 107.205 80.245 107.535 80.615 ;
        RECT 106.800 80.065 106.970 80.210 ;
        RECT 106.345 79.135 106.615 80.040 ;
        RECT 106.800 79.895 107.465 80.065 ;
        RECT 106.785 78.965 107.115 79.725 ;
        RECT 107.295 79.135 107.465 79.895 ;
        RECT 108.645 78.965 108.935 80.130 ;
        RECT 109.545 80.115 109.795 80.715 ;
        RECT 110.045 80.695 110.275 81.515 ;
        RECT 110.525 80.695 110.755 81.515 ;
        RECT 110.925 80.715 111.255 81.345 ;
        RECT 109.965 80.275 110.295 80.525 ;
        RECT 110.505 80.275 110.835 80.525 ;
        RECT 111.005 80.115 111.255 80.715 ;
        RECT 111.425 80.695 111.635 81.515 ;
        RECT 112.325 80.765 113.535 81.515 ;
        RECT 109.165 78.965 109.375 80.105 ;
        RECT 109.545 79.135 109.875 80.115 ;
        RECT 110.045 78.965 110.275 80.105 ;
        RECT 110.525 78.965 110.755 80.105 ;
        RECT 110.925 79.135 111.255 80.115 ;
        RECT 111.425 78.965 111.635 80.105 ;
        RECT 112.325 80.055 112.845 80.595 ;
        RECT 113.015 80.225 113.535 80.765 ;
        RECT 112.325 78.965 113.535 80.055 ;
        RECT 5.520 78.795 113.620 78.965 ;
        RECT 5.605 77.705 6.815 78.795 ;
        RECT 6.985 77.705 8.655 78.795 ;
        RECT 8.915 78.125 9.085 78.625 ;
        RECT 9.255 78.295 9.585 78.795 ;
        RECT 8.915 77.955 9.580 78.125 ;
        RECT 5.605 76.995 6.125 77.535 ;
        RECT 6.295 77.165 6.815 77.705 ;
        RECT 6.985 77.015 7.735 77.535 ;
        RECT 7.905 77.185 8.655 77.705 ;
        RECT 8.830 77.135 9.180 77.785 ;
        RECT 5.605 76.245 6.815 76.995 ;
        RECT 6.985 76.245 8.655 77.015 ;
        RECT 9.350 76.965 9.580 77.955 ;
        RECT 8.915 76.795 9.580 76.965 ;
        RECT 8.915 76.505 9.085 76.795 ;
        RECT 9.255 76.245 9.585 76.625 ;
        RECT 9.755 76.505 9.980 78.625 ;
        RECT 10.195 78.295 10.525 78.795 ;
        RECT 10.695 78.125 10.865 78.625 ;
        RECT 11.100 78.410 11.930 78.580 ;
        RECT 12.170 78.415 12.550 78.795 ;
        RECT 10.170 77.955 10.865 78.125 ;
        RECT 10.170 76.985 10.340 77.955 ;
        RECT 10.510 77.165 10.920 77.785 ;
        RECT 11.090 77.735 11.590 78.115 ;
        RECT 10.170 76.795 10.865 76.985 ;
        RECT 11.090 76.865 11.310 77.735 ;
        RECT 11.760 77.565 11.930 78.410 ;
        RECT 12.730 78.245 12.900 78.535 ;
        RECT 13.070 78.415 13.400 78.795 ;
        RECT 13.870 78.325 14.500 78.575 ;
        RECT 14.680 78.415 15.100 78.795 ;
        RECT 14.330 78.245 14.500 78.325 ;
        RECT 15.300 78.245 15.540 78.535 ;
        RECT 12.100 77.995 13.470 78.245 ;
        RECT 12.100 77.735 12.350 77.995 ;
        RECT 12.860 77.565 13.110 77.725 ;
        RECT 11.760 77.395 13.110 77.565 ;
        RECT 11.760 77.355 12.180 77.395 ;
        RECT 11.490 76.805 11.840 77.175 ;
        RECT 10.195 76.245 10.525 76.625 ;
        RECT 10.695 76.465 10.865 76.795 ;
        RECT 12.010 76.625 12.180 77.355 ;
        RECT 13.280 77.225 13.470 77.995 ;
        RECT 12.350 76.895 12.760 77.225 ;
        RECT 13.050 76.885 13.470 77.225 ;
        RECT 13.640 77.815 14.160 78.125 ;
        RECT 14.330 78.075 15.540 78.245 ;
        RECT 15.770 78.105 16.100 78.795 ;
        RECT 13.640 77.055 13.810 77.815 ;
        RECT 13.980 77.225 14.160 77.635 ;
        RECT 14.330 77.565 14.500 78.075 ;
        RECT 16.270 77.925 16.440 78.535 ;
        RECT 16.710 78.075 17.040 78.585 ;
        RECT 16.270 77.905 16.590 77.925 ;
        RECT 14.670 77.735 16.590 77.905 ;
        RECT 14.330 77.395 16.230 77.565 ;
        RECT 14.560 77.055 14.890 77.175 ;
        RECT 13.640 76.885 14.890 77.055 ;
        RECT 11.165 76.425 12.180 76.625 ;
        RECT 12.350 76.245 12.760 76.685 ;
        RECT 13.050 76.455 13.300 76.885 ;
        RECT 13.500 76.245 13.820 76.705 ;
        RECT 15.060 76.635 15.230 77.395 ;
        RECT 15.900 77.335 16.230 77.395 ;
        RECT 15.420 77.165 15.750 77.225 ;
        RECT 15.420 76.895 16.080 77.165 ;
        RECT 16.400 76.840 16.590 77.735 ;
        RECT 14.380 76.465 15.230 76.635 ;
        RECT 15.430 76.245 16.090 76.725 ;
        RECT 16.270 76.510 16.590 76.840 ;
        RECT 16.790 77.485 17.040 78.075 ;
        RECT 17.220 77.995 17.505 78.795 ;
        RECT 17.685 77.815 17.940 78.485 ;
        RECT 16.790 77.155 17.590 77.485 ;
        RECT 16.790 76.505 17.040 77.155 ;
        RECT 17.760 76.955 17.940 77.815 ;
        RECT 18.485 77.630 18.775 78.795 ;
        RECT 19.005 77.655 19.215 78.795 ;
        RECT 19.385 77.645 19.715 78.625 ;
        RECT 19.885 77.655 20.115 78.795 ;
        RECT 20.325 77.705 21.995 78.795 ;
        RECT 22.170 78.285 23.825 78.575 ;
        RECT 17.685 76.755 17.940 76.955 ;
        RECT 17.220 76.245 17.505 76.705 ;
        RECT 17.685 76.585 18.025 76.755 ;
        RECT 17.685 76.425 17.940 76.585 ;
        RECT 18.485 76.245 18.775 76.970 ;
        RECT 19.005 76.245 19.215 77.065 ;
        RECT 19.385 77.045 19.635 77.645 ;
        RECT 19.805 77.235 20.135 77.485 ;
        RECT 19.385 76.415 19.715 77.045 ;
        RECT 19.885 76.245 20.115 77.065 ;
        RECT 20.325 77.015 21.075 77.535 ;
        RECT 21.245 77.185 21.995 77.705 ;
        RECT 22.170 77.945 23.760 78.115 ;
        RECT 23.995 77.995 24.275 78.795 ;
        RECT 22.170 77.655 22.490 77.945 ;
        RECT 23.590 77.825 23.760 77.945 ;
        RECT 22.685 77.605 23.400 77.775 ;
        RECT 23.590 77.655 24.315 77.825 ;
        RECT 24.485 77.655 24.755 78.625 ;
        RECT 24.930 78.285 26.585 78.575 ;
        RECT 24.930 77.945 26.520 78.115 ;
        RECT 26.755 77.995 27.035 78.795 ;
        RECT 24.930 77.655 25.250 77.945 ;
        RECT 26.350 77.825 26.520 77.945 ;
        RECT 20.325 76.245 21.995 77.015 ;
        RECT 22.170 76.915 22.520 77.485 ;
        RECT 22.690 77.155 23.400 77.605 ;
        RECT 24.145 77.485 24.315 77.655 ;
        RECT 23.570 77.155 23.975 77.485 ;
        RECT 24.145 77.155 24.415 77.485 ;
        RECT 24.145 76.985 24.315 77.155 ;
        RECT 22.705 76.815 24.315 76.985 ;
        RECT 24.585 76.920 24.755 77.655 ;
        RECT 25.445 77.605 26.160 77.775 ;
        RECT 26.350 77.655 27.075 77.825 ;
        RECT 27.245 77.655 27.515 78.625 ;
        RECT 27.685 78.360 33.030 78.795 ;
        RECT 33.205 78.360 38.550 78.795 ;
        RECT 22.175 76.245 22.505 76.745 ;
        RECT 22.705 76.465 22.875 76.815 ;
        RECT 23.075 76.245 23.405 76.645 ;
        RECT 23.575 76.465 23.745 76.815 ;
        RECT 23.915 76.245 24.295 76.645 ;
        RECT 24.485 76.575 24.755 76.920 ;
        RECT 24.930 76.915 25.280 77.485 ;
        RECT 25.450 77.155 26.160 77.605 ;
        RECT 26.905 77.485 27.075 77.655 ;
        RECT 26.330 77.155 26.735 77.485 ;
        RECT 26.905 77.155 27.175 77.485 ;
        RECT 26.905 76.985 27.075 77.155 ;
        RECT 25.465 76.815 27.075 76.985 ;
        RECT 27.345 76.920 27.515 77.655 ;
        RECT 24.935 76.245 25.265 76.745 ;
        RECT 25.465 76.465 25.635 76.815 ;
        RECT 25.835 76.245 26.165 76.645 ;
        RECT 26.335 76.465 26.505 76.815 ;
        RECT 26.675 76.245 27.055 76.645 ;
        RECT 27.245 76.575 27.515 76.920 ;
        RECT 29.270 76.790 29.610 77.620 ;
        RECT 31.090 77.110 31.440 78.360 ;
        RECT 34.790 76.790 35.130 77.620 ;
        RECT 36.610 77.110 36.960 78.360 ;
        RECT 38.725 77.705 41.315 78.795 ;
        RECT 38.725 77.015 39.935 77.535 ;
        RECT 40.105 77.185 41.315 77.705 ;
        RECT 41.525 77.655 41.755 78.795 ;
        RECT 41.925 77.645 42.255 78.625 ;
        RECT 42.425 77.655 42.635 78.795 ;
        RECT 42.865 77.705 44.075 78.795 ;
        RECT 41.505 77.235 41.835 77.485 ;
        RECT 27.685 76.245 33.030 76.790 ;
        RECT 33.205 76.245 38.550 76.790 ;
        RECT 38.725 76.245 41.315 77.015 ;
        RECT 41.525 76.245 41.755 77.065 ;
        RECT 42.005 77.045 42.255 77.645 ;
        RECT 41.925 76.415 42.255 77.045 ;
        RECT 42.425 76.245 42.635 77.065 ;
        RECT 42.865 76.995 43.385 77.535 ;
        RECT 43.555 77.165 44.075 77.705 ;
        RECT 44.245 77.630 44.535 78.795 ;
        RECT 44.705 78.360 50.050 78.795 ;
        RECT 42.865 76.245 44.075 76.995 ;
        RECT 44.245 76.245 44.535 76.970 ;
        RECT 46.290 76.790 46.630 77.620 ;
        RECT 48.110 77.110 48.460 78.360 ;
        RECT 51.235 78.125 51.405 78.625 ;
        RECT 51.575 78.295 51.905 78.795 ;
        RECT 51.235 77.955 51.900 78.125 ;
        RECT 51.150 77.135 51.500 77.785 ;
        RECT 51.670 76.965 51.900 77.955 ;
        RECT 51.235 76.795 51.900 76.965 ;
        RECT 44.705 76.245 50.050 76.790 ;
        RECT 51.235 76.505 51.405 76.795 ;
        RECT 51.575 76.245 51.905 76.625 ;
        RECT 52.075 76.505 52.300 78.625 ;
        RECT 52.515 78.295 52.845 78.795 ;
        RECT 53.015 78.125 53.185 78.625 ;
        RECT 53.420 78.410 54.250 78.580 ;
        RECT 54.490 78.415 54.870 78.795 ;
        RECT 52.490 77.955 53.185 78.125 ;
        RECT 52.490 76.985 52.660 77.955 ;
        RECT 52.830 77.165 53.240 77.785 ;
        RECT 53.410 77.735 53.910 78.115 ;
        RECT 52.490 76.795 53.185 76.985 ;
        RECT 53.410 76.865 53.630 77.735 ;
        RECT 54.080 77.565 54.250 78.410 ;
        RECT 55.050 78.245 55.220 78.535 ;
        RECT 55.390 78.415 55.720 78.795 ;
        RECT 56.190 78.325 56.820 78.575 ;
        RECT 57.000 78.415 57.420 78.795 ;
        RECT 56.650 78.245 56.820 78.325 ;
        RECT 57.620 78.245 57.860 78.535 ;
        RECT 54.420 77.995 55.790 78.245 ;
        RECT 54.420 77.735 54.670 77.995 ;
        RECT 55.180 77.565 55.430 77.725 ;
        RECT 54.080 77.395 55.430 77.565 ;
        RECT 54.080 77.355 54.500 77.395 ;
        RECT 53.810 76.805 54.160 77.175 ;
        RECT 52.515 76.245 52.845 76.625 ;
        RECT 53.015 76.465 53.185 76.795 ;
        RECT 54.330 76.625 54.500 77.355 ;
        RECT 55.600 77.225 55.790 77.995 ;
        RECT 54.670 76.895 55.080 77.225 ;
        RECT 55.370 76.885 55.790 77.225 ;
        RECT 55.960 77.815 56.480 78.125 ;
        RECT 56.650 78.075 57.860 78.245 ;
        RECT 58.090 78.105 58.420 78.795 ;
        RECT 55.960 77.055 56.130 77.815 ;
        RECT 56.300 77.225 56.480 77.635 ;
        RECT 56.650 77.565 56.820 78.075 ;
        RECT 58.590 77.925 58.760 78.535 ;
        RECT 59.030 78.075 59.360 78.585 ;
        RECT 58.590 77.905 58.910 77.925 ;
        RECT 56.990 77.735 58.910 77.905 ;
        RECT 56.650 77.395 58.550 77.565 ;
        RECT 56.880 77.055 57.210 77.175 ;
        RECT 55.960 76.885 57.210 77.055 ;
        RECT 53.485 76.425 54.500 76.625 ;
        RECT 54.670 76.245 55.080 76.685 ;
        RECT 55.370 76.455 55.620 76.885 ;
        RECT 55.820 76.245 56.140 76.705 ;
        RECT 57.380 76.635 57.550 77.395 ;
        RECT 58.220 77.335 58.550 77.395 ;
        RECT 57.740 77.165 58.070 77.225 ;
        RECT 57.740 76.895 58.400 77.165 ;
        RECT 58.720 76.840 58.910 77.735 ;
        RECT 56.700 76.465 57.550 76.635 ;
        RECT 57.750 76.245 58.410 76.725 ;
        RECT 58.590 76.510 58.910 76.840 ;
        RECT 59.110 77.485 59.360 78.075 ;
        RECT 59.540 77.995 59.825 78.795 ;
        RECT 60.005 77.815 60.260 78.485 ;
        RECT 60.080 77.775 60.260 77.815 ;
        RECT 60.080 77.605 60.345 77.775 ;
        RECT 60.810 77.655 61.145 78.625 ;
        RECT 61.315 77.655 61.485 78.795 ;
        RECT 61.655 78.455 63.685 78.625 ;
        RECT 59.110 77.155 59.910 77.485 ;
        RECT 59.110 76.505 59.360 77.155 ;
        RECT 60.080 76.955 60.260 77.605 ;
        RECT 59.540 76.245 59.825 76.705 ;
        RECT 60.005 76.425 60.260 76.955 ;
        RECT 60.810 76.985 60.980 77.655 ;
        RECT 61.655 77.485 61.825 78.455 ;
        RECT 61.150 77.155 61.405 77.485 ;
        RECT 61.630 77.155 61.825 77.485 ;
        RECT 61.995 78.115 63.120 78.285 ;
        RECT 61.235 76.985 61.405 77.155 ;
        RECT 61.995 76.985 62.165 78.115 ;
        RECT 60.810 76.415 61.065 76.985 ;
        RECT 61.235 76.815 62.165 76.985 ;
        RECT 62.335 77.775 63.345 77.945 ;
        RECT 62.335 76.975 62.505 77.775 ;
        RECT 62.710 77.435 62.985 77.575 ;
        RECT 62.705 77.265 62.985 77.435 ;
        RECT 61.990 76.780 62.165 76.815 ;
        RECT 61.235 76.245 61.565 76.645 ;
        RECT 61.990 76.415 62.520 76.780 ;
        RECT 62.710 76.415 62.985 77.265 ;
        RECT 63.155 76.415 63.345 77.775 ;
        RECT 63.515 77.790 63.685 78.455 ;
        RECT 63.855 78.035 64.025 78.795 ;
        RECT 64.260 78.035 64.775 78.445 ;
        RECT 63.515 77.600 64.265 77.790 ;
        RECT 64.435 77.225 64.775 78.035 ;
        RECT 65.150 77.825 65.480 78.625 ;
        RECT 65.650 77.995 65.980 78.795 ;
        RECT 66.280 77.825 66.610 78.625 ;
        RECT 67.255 77.995 67.505 78.795 ;
        RECT 65.150 77.655 67.585 77.825 ;
        RECT 67.775 77.655 67.945 78.795 ;
        RECT 68.115 77.655 68.455 78.625 ;
        RECT 68.685 77.655 68.895 78.795 ;
        RECT 64.945 77.235 65.295 77.485 ;
        RECT 63.545 77.055 64.775 77.225 ;
        RECT 63.525 76.245 64.035 76.780 ;
        RECT 64.255 76.450 64.500 77.055 ;
        RECT 65.480 77.025 65.650 77.655 ;
        RECT 65.820 77.235 66.150 77.435 ;
        RECT 66.320 77.235 66.650 77.435 ;
        RECT 66.820 77.235 67.240 77.435 ;
        RECT 67.415 77.405 67.585 77.655 ;
        RECT 67.415 77.235 68.110 77.405 ;
        RECT 65.150 76.415 65.650 77.025 ;
        RECT 66.280 76.895 67.505 77.065 ;
        RECT 68.280 77.045 68.455 77.655 ;
        RECT 69.065 77.645 69.395 78.625 ;
        RECT 69.565 77.655 69.795 78.795 ;
        RECT 66.280 76.415 66.610 76.895 ;
        RECT 66.780 76.245 67.005 76.705 ;
        RECT 67.175 76.415 67.505 76.895 ;
        RECT 67.695 76.245 67.945 77.045 ;
        RECT 68.115 76.415 68.455 77.045 ;
        RECT 68.685 76.245 68.895 77.065 ;
        RECT 69.065 77.045 69.315 77.645 ;
        RECT 70.005 77.630 70.295 78.795 ;
        RECT 70.465 78.360 75.810 78.795 ;
        RECT 69.485 77.235 69.815 77.485 ;
        RECT 69.065 76.415 69.395 77.045 ;
        RECT 69.565 76.245 69.795 77.065 ;
        RECT 70.005 76.245 70.295 76.970 ;
        RECT 72.050 76.790 72.390 77.620 ;
        RECT 73.870 77.110 74.220 78.360 ;
        RECT 76.995 77.865 77.165 78.625 ;
        RECT 77.345 78.035 77.675 78.795 ;
        RECT 76.995 77.695 77.660 77.865 ;
        RECT 77.845 77.720 78.115 78.625 ;
        RECT 77.490 77.550 77.660 77.695 ;
        RECT 76.925 77.145 77.255 77.515 ;
        RECT 77.490 77.220 77.775 77.550 ;
        RECT 77.490 76.965 77.660 77.220 ;
        RECT 76.995 76.795 77.660 76.965 ;
        RECT 77.945 76.920 78.115 77.720 ;
        RECT 70.465 76.245 75.810 76.790 ;
        RECT 76.995 76.415 77.165 76.795 ;
        RECT 77.345 76.245 77.675 76.625 ;
        RECT 77.855 76.415 78.115 76.920 ;
        RECT 78.745 77.655 79.015 78.625 ;
        RECT 79.225 77.995 79.505 78.795 ;
        RECT 79.675 78.285 81.330 78.575 ;
        RECT 81.505 78.360 86.850 78.795 ;
        RECT 79.740 77.945 81.330 78.115 ;
        RECT 79.740 77.825 79.910 77.945 ;
        RECT 79.185 77.655 79.910 77.825 ;
        RECT 78.745 76.920 78.915 77.655 ;
        RECT 79.185 77.485 79.355 77.655 ;
        RECT 79.085 77.155 79.355 77.485 ;
        RECT 79.525 77.155 79.930 77.485 ;
        RECT 80.100 77.155 80.810 77.775 ;
        RECT 81.010 77.655 81.330 77.945 ;
        RECT 79.185 76.985 79.355 77.155 ;
        RECT 78.745 76.575 79.015 76.920 ;
        RECT 79.185 76.815 80.795 76.985 ;
        RECT 80.980 76.915 81.330 77.485 ;
        RECT 79.205 76.245 79.585 76.645 ;
        RECT 79.755 76.465 79.925 76.815 ;
        RECT 80.095 76.245 80.425 76.645 ;
        RECT 80.625 76.465 80.795 76.815 ;
        RECT 83.090 76.790 83.430 77.620 ;
        RECT 84.910 77.110 85.260 78.360 ;
        RECT 87.025 77.705 88.695 78.795 ;
        RECT 87.025 77.015 87.775 77.535 ;
        RECT 87.945 77.185 88.695 77.705 ;
        RECT 89.325 78.075 89.785 78.625 ;
        RECT 89.975 78.075 90.305 78.795 ;
        RECT 80.995 76.245 81.325 76.745 ;
        RECT 81.505 76.245 86.850 76.790 ;
        RECT 87.025 76.245 88.695 77.015 ;
        RECT 89.325 76.705 89.575 78.075 ;
        RECT 90.505 77.905 90.805 78.455 ;
        RECT 90.975 78.125 91.255 78.795 ;
        RECT 89.865 77.735 90.805 77.905 ;
        RECT 91.625 78.075 92.085 78.625 ;
        RECT 92.275 78.075 92.605 78.795 ;
        RECT 89.865 77.485 90.035 77.735 ;
        RECT 91.175 77.485 91.440 77.845 ;
        RECT 89.745 77.155 90.035 77.485 ;
        RECT 90.205 77.235 90.545 77.485 ;
        RECT 90.765 77.235 91.440 77.485 ;
        RECT 89.865 77.065 90.035 77.155 ;
        RECT 89.865 76.875 91.255 77.065 ;
        RECT 89.325 76.415 89.885 76.705 ;
        RECT 90.055 76.245 90.305 76.705 ;
        RECT 90.925 76.515 91.255 76.875 ;
        RECT 91.625 76.705 91.875 78.075 ;
        RECT 92.805 77.905 93.105 78.455 ;
        RECT 93.275 78.125 93.555 78.795 ;
        RECT 92.165 77.735 93.105 77.905 ;
        RECT 92.165 77.485 92.335 77.735 ;
        RECT 93.475 77.485 93.740 77.845 ;
        RECT 93.925 77.705 95.595 78.795 ;
        RECT 92.045 77.155 92.335 77.485 ;
        RECT 92.505 77.235 92.845 77.485 ;
        RECT 93.065 77.235 93.740 77.485 ;
        RECT 92.165 77.065 92.335 77.155 ;
        RECT 92.165 76.875 93.555 77.065 ;
        RECT 91.625 76.415 92.185 76.705 ;
        RECT 92.355 76.245 92.605 76.705 ;
        RECT 93.225 76.515 93.555 76.875 ;
        RECT 93.925 77.015 94.675 77.535 ;
        RECT 94.845 77.185 95.595 77.705 ;
        RECT 95.765 77.630 96.055 78.795 ;
        RECT 96.230 77.655 96.565 78.625 ;
        RECT 96.735 77.655 96.905 78.795 ;
        RECT 97.075 78.455 99.105 78.625 ;
        RECT 93.925 76.245 95.595 77.015 ;
        RECT 96.230 76.985 96.400 77.655 ;
        RECT 97.075 77.485 97.245 78.455 ;
        RECT 96.570 77.155 96.825 77.485 ;
        RECT 97.050 77.155 97.245 77.485 ;
        RECT 97.415 78.115 98.540 78.285 ;
        RECT 96.655 76.985 96.825 77.155 ;
        RECT 97.415 76.985 97.585 78.115 ;
        RECT 95.765 76.245 96.055 76.970 ;
        RECT 96.230 76.415 96.485 76.985 ;
        RECT 96.655 76.815 97.585 76.985 ;
        RECT 97.755 77.775 98.765 77.945 ;
        RECT 97.755 76.975 97.925 77.775 ;
        RECT 97.410 76.780 97.585 76.815 ;
        RECT 96.655 76.245 96.985 76.645 ;
        RECT 97.410 76.415 97.940 76.780 ;
        RECT 98.130 76.755 98.405 77.575 ;
        RECT 98.125 76.585 98.405 76.755 ;
        RECT 98.130 76.415 98.405 76.585 ;
        RECT 98.575 76.415 98.765 77.775 ;
        RECT 98.935 77.790 99.105 78.455 ;
        RECT 99.275 78.035 99.445 78.795 ;
        RECT 99.680 78.035 100.195 78.445 ;
        RECT 98.935 77.600 99.685 77.790 ;
        RECT 99.855 77.225 100.195 78.035 ;
        RECT 100.915 78.125 101.085 78.625 ;
        RECT 101.255 78.295 101.585 78.795 ;
        RECT 100.915 77.955 101.580 78.125 ;
        RECT 98.965 77.055 100.195 77.225 ;
        RECT 100.830 77.135 101.180 77.785 ;
        RECT 98.945 76.245 99.455 76.780 ;
        RECT 99.675 76.450 99.920 77.055 ;
        RECT 101.350 76.965 101.580 77.955 ;
        RECT 100.915 76.795 101.580 76.965 ;
        RECT 100.915 76.505 101.085 76.795 ;
        RECT 101.255 76.245 101.585 76.625 ;
        RECT 101.755 76.505 101.980 78.625 ;
        RECT 102.195 78.295 102.525 78.795 ;
        RECT 102.695 78.125 102.865 78.625 ;
        RECT 103.100 78.410 103.930 78.580 ;
        RECT 104.170 78.415 104.550 78.795 ;
        RECT 102.170 77.955 102.865 78.125 ;
        RECT 102.170 76.985 102.340 77.955 ;
        RECT 102.510 77.165 102.920 77.785 ;
        RECT 103.090 77.735 103.590 78.115 ;
        RECT 102.170 76.795 102.865 76.985 ;
        RECT 103.090 76.865 103.310 77.735 ;
        RECT 103.760 77.565 103.930 78.410 ;
        RECT 104.730 78.245 104.900 78.535 ;
        RECT 105.070 78.415 105.400 78.795 ;
        RECT 105.870 78.325 106.500 78.575 ;
        RECT 106.680 78.415 107.100 78.795 ;
        RECT 106.330 78.245 106.500 78.325 ;
        RECT 107.300 78.245 107.540 78.535 ;
        RECT 104.100 77.995 105.470 78.245 ;
        RECT 104.100 77.735 104.350 77.995 ;
        RECT 104.860 77.565 105.110 77.725 ;
        RECT 103.760 77.395 105.110 77.565 ;
        RECT 103.760 77.355 104.180 77.395 ;
        RECT 103.490 76.805 103.840 77.175 ;
        RECT 102.195 76.245 102.525 76.625 ;
        RECT 102.695 76.465 102.865 76.795 ;
        RECT 104.010 76.625 104.180 77.355 ;
        RECT 105.280 77.225 105.470 77.995 ;
        RECT 104.350 76.895 104.760 77.225 ;
        RECT 105.050 76.885 105.470 77.225 ;
        RECT 105.640 77.815 106.160 78.125 ;
        RECT 106.330 78.075 107.540 78.245 ;
        RECT 107.770 78.105 108.100 78.795 ;
        RECT 105.640 77.055 105.810 77.815 ;
        RECT 105.980 77.225 106.160 77.635 ;
        RECT 106.330 77.565 106.500 78.075 ;
        RECT 108.270 77.925 108.440 78.535 ;
        RECT 108.710 78.075 109.040 78.585 ;
        RECT 108.270 77.905 108.590 77.925 ;
        RECT 106.670 77.735 108.590 77.905 ;
        RECT 106.330 77.395 108.230 77.565 ;
        RECT 106.560 77.055 106.890 77.175 ;
        RECT 105.640 76.885 106.890 77.055 ;
        RECT 103.165 76.425 104.180 76.625 ;
        RECT 104.350 76.245 104.760 76.685 ;
        RECT 105.050 76.455 105.300 76.885 ;
        RECT 105.500 76.245 105.820 76.705 ;
        RECT 107.060 76.635 107.230 77.395 ;
        RECT 107.900 77.335 108.230 77.395 ;
        RECT 107.420 77.165 107.750 77.225 ;
        RECT 107.420 76.895 108.080 77.165 ;
        RECT 108.400 76.840 108.590 77.735 ;
        RECT 106.380 76.465 107.230 76.635 ;
        RECT 107.430 76.245 108.090 76.725 ;
        RECT 108.270 76.510 108.590 76.840 ;
        RECT 108.790 77.485 109.040 78.075 ;
        RECT 109.220 77.995 109.505 78.795 ;
        RECT 109.685 77.815 109.940 78.485 ;
        RECT 109.760 77.775 109.940 77.815 ;
        RECT 109.760 77.605 110.025 77.775 ;
        RECT 110.485 77.705 112.155 78.795 ;
        RECT 108.790 77.155 109.590 77.485 ;
        RECT 108.790 76.505 109.040 77.155 ;
        RECT 109.760 76.955 109.940 77.605 ;
        RECT 109.220 76.245 109.505 76.705 ;
        RECT 109.685 76.425 109.940 76.955 ;
        RECT 110.485 77.015 111.235 77.535 ;
        RECT 111.405 77.185 112.155 77.705 ;
        RECT 112.325 77.705 113.535 78.795 ;
        RECT 112.325 77.165 112.845 77.705 ;
        RECT 110.485 76.245 112.155 77.015 ;
        RECT 113.015 76.995 113.535 77.535 ;
        RECT 112.325 76.245 113.535 76.995 ;
        RECT 5.520 76.075 113.620 76.245 ;
        RECT 5.605 75.325 6.815 76.075 ;
        RECT 7.075 75.525 7.245 75.815 ;
        RECT 7.415 75.695 7.745 76.075 ;
        RECT 7.075 75.355 7.740 75.525 ;
        RECT 5.605 74.785 6.125 75.325 ;
        RECT 6.295 74.615 6.815 75.155 ;
        RECT 5.605 73.525 6.815 74.615 ;
        RECT 6.990 74.535 7.340 75.185 ;
        RECT 7.510 74.365 7.740 75.355 ;
        RECT 7.075 74.195 7.740 74.365 ;
        RECT 7.075 73.695 7.245 74.195 ;
        RECT 7.415 73.525 7.745 74.025 ;
        RECT 7.915 73.695 8.140 75.815 ;
        RECT 8.355 75.695 8.685 76.075 ;
        RECT 8.855 75.525 9.025 75.855 ;
        RECT 9.325 75.695 10.340 75.895 ;
        RECT 8.330 75.335 9.025 75.525 ;
        RECT 8.330 74.365 8.500 75.335 ;
        RECT 8.670 74.535 9.080 75.155 ;
        RECT 9.250 74.585 9.470 75.455 ;
        RECT 9.650 75.145 10.000 75.515 ;
        RECT 10.170 74.965 10.340 75.695 ;
        RECT 10.510 75.635 10.920 76.075 ;
        RECT 11.210 75.435 11.460 75.865 ;
        RECT 11.660 75.615 11.980 76.075 ;
        RECT 12.540 75.685 13.390 75.855 ;
        RECT 10.510 75.095 10.920 75.425 ;
        RECT 11.210 75.095 11.630 75.435 ;
        RECT 9.920 74.925 10.340 74.965 ;
        RECT 9.920 74.755 11.270 74.925 ;
        RECT 8.330 74.195 9.025 74.365 ;
        RECT 9.250 74.205 9.750 74.585 ;
        RECT 8.355 73.525 8.685 74.025 ;
        RECT 8.855 73.695 9.025 74.195 ;
        RECT 9.920 73.910 10.090 74.755 ;
        RECT 11.020 74.595 11.270 74.755 ;
        RECT 10.260 74.325 10.510 74.585 ;
        RECT 11.440 74.325 11.630 75.095 ;
        RECT 10.260 74.075 11.630 74.325 ;
        RECT 11.800 75.265 13.050 75.435 ;
        RECT 11.800 74.505 11.970 75.265 ;
        RECT 12.720 75.145 13.050 75.265 ;
        RECT 12.140 74.685 12.320 75.095 ;
        RECT 13.220 74.925 13.390 75.685 ;
        RECT 13.590 75.595 14.250 76.075 ;
        RECT 14.430 75.480 14.750 75.810 ;
        RECT 13.580 75.155 14.240 75.425 ;
        RECT 13.580 75.095 13.910 75.155 ;
        RECT 14.060 74.925 14.390 74.985 ;
        RECT 12.490 74.755 14.390 74.925 ;
        RECT 11.800 74.195 12.320 74.505 ;
        RECT 12.490 74.245 12.660 74.755 ;
        RECT 14.560 74.585 14.750 75.480 ;
        RECT 12.830 74.415 14.750 74.585 ;
        RECT 14.430 74.395 14.750 74.415 ;
        RECT 14.950 75.165 15.200 75.815 ;
        RECT 15.380 75.615 15.665 76.075 ;
        RECT 15.845 75.395 16.100 75.895 ;
        RECT 15.845 75.365 16.185 75.395 ;
        RECT 15.920 75.225 16.185 75.365 ;
        RECT 16.650 75.335 16.905 75.905 ;
        RECT 17.075 75.675 17.405 76.075 ;
        RECT 17.830 75.540 18.360 75.905 ;
        RECT 17.830 75.505 18.005 75.540 ;
        RECT 17.075 75.335 18.005 75.505 ;
        RECT 14.950 74.835 15.750 75.165 ;
        RECT 12.490 74.075 13.700 74.245 ;
        RECT 9.260 73.740 10.090 73.910 ;
        RECT 10.330 73.525 10.710 73.905 ;
        RECT 10.890 73.785 11.060 74.075 ;
        RECT 12.490 73.995 12.660 74.075 ;
        RECT 11.230 73.525 11.560 73.905 ;
        RECT 12.030 73.745 12.660 73.995 ;
        RECT 12.840 73.525 13.260 73.905 ;
        RECT 13.460 73.785 13.700 74.075 ;
        RECT 13.930 73.525 14.260 74.215 ;
        RECT 14.430 73.785 14.600 74.395 ;
        RECT 14.950 74.245 15.200 74.835 ;
        RECT 15.920 74.505 16.100 75.225 ;
        RECT 14.870 73.735 15.200 74.245 ;
        RECT 15.380 73.525 15.665 74.325 ;
        RECT 15.845 73.835 16.100 74.505 ;
        RECT 16.650 74.665 16.820 75.335 ;
        RECT 17.075 75.165 17.245 75.335 ;
        RECT 16.990 74.835 17.245 75.165 ;
        RECT 17.470 74.835 17.665 75.165 ;
        RECT 16.650 73.695 16.985 74.665 ;
        RECT 17.155 73.525 17.325 74.665 ;
        RECT 17.495 73.865 17.665 74.835 ;
        RECT 17.835 74.205 18.005 75.335 ;
        RECT 18.175 74.545 18.345 75.345 ;
        RECT 18.550 75.055 18.825 75.905 ;
        RECT 18.545 74.885 18.825 75.055 ;
        RECT 18.550 74.745 18.825 74.885 ;
        RECT 18.995 74.545 19.185 75.905 ;
        RECT 19.365 75.540 19.875 76.075 ;
        RECT 20.095 75.265 20.340 75.870 ;
        RECT 20.785 75.305 22.455 76.075 ;
        RECT 19.385 75.095 20.615 75.265 ;
        RECT 18.175 74.375 19.185 74.545 ;
        RECT 19.355 74.530 20.105 74.720 ;
        RECT 17.835 74.035 18.960 74.205 ;
        RECT 19.355 73.865 19.525 74.530 ;
        RECT 20.275 74.285 20.615 75.095 ;
        RECT 20.785 74.785 21.535 75.305 ;
        RECT 22.830 75.295 23.330 75.905 ;
        RECT 21.705 74.615 22.455 75.135 ;
        RECT 22.625 74.835 22.975 75.085 ;
        RECT 23.160 74.665 23.330 75.295 ;
        RECT 23.960 75.425 24.290 75.905 ;
        RECT 24.460 75.615 24.685 76.075 ;
        RECT 24.855 75.425 25.185 75.905 ;
        RECT 23.960 75.255 25.185 75.425 ;
        RECT 25.375 75.275 25.625 76.075 ;
        RECT 25.795 75.275 26.135 75.905 ;
        RECT 23.500 74.885 23.830 75.085 ;
        RECT 24.000 74.885 24.330 75.085 ;
        RECT 24.500 74.885 24.920 75.085 ;
        RECT 25.095 74.915 25.790 75.085 ;
        RECT 25.095 74.665 25.265 74.915 ;
        RECT 25.960 74.665 26.135 75.275 ;
        RECT 26.305 75.305 29.815 76.075 ;
        RECT 29.985 75.325 31.195 76.075 ;
        RECT 31.365 75.350 31.655 76.075 ;
        RECT 26.305 74.785 27.955 75.305 ;
        RECT 17.495 73.695 19.525 73.865 ;
        RECT 19.695 73.525 19.865 74.285 ;
        RECT 20.100 73.875 20.615 74.285 ;
        RECT 20.785 73.525 22.455 74.615 ;
        RECT 22.830 74.495 25.265 74.665 ;
        RECT 22.830 73.695 23.160 74.495 ;
        RECT 23.330 73.525 23.660 74.325 ;
        RECT 23.960 73.695 24.290 74.495 ;
        RECT 24.935 73.525 25.185 74.325 ;
        RECT 25.455 73.525 25.625 74.665 ;
        RECT 25.795 73.695 26.135 74.665 ;
        RECT 28.125 74.615 29.815 75.135 ;
        RECT 29.985 74.785 30.505 75.325 ;
        RECT 31.825 75.275 32.165 75.905 ;
        RECT 32.335 75.275 32.585 76.075 ;
        RECT 32.775 75.425 33.105 75.905 ;
        RECT 33.275 75.615 33.500 76.075 ;
        RECT 33.670 75.425 34.000 75.905 ;
        RECT 30.675 74.615 31.195 75.155 ;
        RECT 26.305 73.525 29.815 74.615 ;
        RECT 29.985 73.525 31.195 74.615 ;
        RECT 31.365 73.525 31.655 74.690 ;
        RECT 31.825 74.665 32.000 75.275 ;
        RECT 32.775 75.255 34.000 75.425 ;
        RECT 34.630 75.295 35.130 75.905 ;
        RECT 35.505 75.305 37.175 76.075 ;
        RECT 37.895 75.525 38.065 75.815 ;
        RECT 38.235 75.695 38.565 76.075 ;
        RECT 37.895 75.355 38.560 75.525 ;
        RECT 32.170 74.915 32.865 75.085 ;
        RECT 32.695 74.665 32.865 74.915 ;
        RECT 33.040 74.885 33.460 75.085 ;
        RECT 33.630 74.885 33.960 75.085 ;
        RECT 34.130 74.885 34.460 75.085 ;
        RECT 34.630 74.665 34.800 75.295 ;
        RECT 34.985 74.835 35.335 75.085 ;
        RECT 35.505 74.785 36.255 75.305 ;
        RECT 31.825 73.695 32.165 74.665 ;
        RECT 32.335 73.525 32.505 74.665 ;
        RECT 32.695 74.495 35.130 74.665 ;
        RECT 36.425 74.615 37.175 75.135 ;
        RECT 32.775 73.525 33.025 74.325 ;
        RECT 33.670 73.695 34.000 74.495 ;
        RECT 34.300 73.525 34.630 74.325 ;
        RECT 34.800 73.695 35.130 74.495 ;
        RECT 35.505 73.525 37.175 74.615 ;
        RECT 37.810 74.535 38.160 75.185 ;
        RECT 38.330 74.365 38.560 75.355 ;
        RECT 37.895 74.195 38.560 74.365 ;
        RECT 37.895 73.695 38.065 74.195 ;
        RECT 38.235 73.525 38.565 74.025 ;
        RECT 38.735 73.695 38.960 75.815 ;
        RECT 39.175 75.695 39.505 76.075 ;
        RECT 39.675 75.525 39.845 75.855 ;
        RECT 40.145 75.695 41.160 75.895 ;
        RECT 39.150 75.335 39.845 75.525 ;
        RECT 39.150 74.365 39.320 75.335 ;
        RECT 39.490 74.535 39.900 75.155 ;
        RECT 40.070 74.585 40.290 75.455 ;
        RECT 40.470 75.145 40.820 75.515 ;
        RECT 40.990 74.965 41.160 75.695 ;
        RECT 41.330 75.635 41.740 76.075 ;
        RECT 42.030 75.435 42.280 75.865 ;
        RECT 42.480 75.615 42.800 76.075 ;
        RECT 43.360 75.685 44.210 75.855 ;
        RECT 41.330 75.095 41.740 75.425 ;
        RECT 42.030 75.095 42.450 75.435 ;
        RECT 40.740 74.925 41.160 74.965 ;
        RECT 40.740 74.755 42.090 74.925 ;
        RECT 39.150 74.195 39.845 74.365 ;
        RECT 40.070 74.205 40.570 74.585 ;
        RECT 39.175 73.525 39.505 74.025 ;
        RECT 39.675 73.695 39.845 74.195 ;
        RECT 40.740 73.910 40.910 74.755 ;
        RECT 41.840 74.595 42.090 74.755 ;
        RECT 41.080 74.325 41.330 74.585 ;
        RECT 42.260 74.325 42.450 75.095 ;
        RECT 41.080 74.075 42.450 74.325 ;
        RECT 42.620 75.265 43.870 75.435 ;
        RECT 42.620 74.505 42.790 75.265 ;
        RECT 43.540 75.145 43.870 75.265 ;
        RECT 42.960 74.685 43.140 75.095 ;
        RECT 44.040 74.925 44.210 75.685 ;
        RECT 44.410 75.595 45.070 76.075 ;
        RECT 45.250 75.480 45.570 75.810 ;
        RECT 44.400 75.155 45.060 75.425 ;
        RECT 44.400 75.095 44.730 75.155 ;
        RECT 44.880 74.925 45.210 74.985 ;
        RECT 43.310 74.755 45.210 74.925 ;
        RECT 42.620 74.195 43.140 74.505 ;
        RECT 43.310 74.245 43.480 74.755 ;
        RECT 45.380 74.585 45.570 75.480 ;
        RECT 43.650 74.415 45.570 74.585 ;
        RECT 45.250 74.395 45.570 74.415 ;
        RECT 45.770 75.165 46.020 75.815 ;
        RECT 46.200 75.615 46.485 76.075 ;
        RECT 46.665 75.365 46.920 75.895 ;
        RECT 45.770 74.835 46.570 75.165 ;
        RECT 43.310 74.075 44.520 74.245 ;
        RECT 40.080 73.740 40.910 73.910 ;
        RECT 41.150 73.525 41.530 73.905 ;
        RECT 41.710 73.785 41.880 74.075 ;
        RECT 43.310 73.995 43.480 74.075 ;
        RECT 42.050 73.525 42.380 73.905 ;
        RECT 42.850 73.745 43.480 73.995 ;
        RECT 43.660 73.525 44.080 73.905 ;
        RECT 44.280 73.785 44.520 74.075 ;
        RECT 44.750 73.525 45.080 74.215 ;
        RECT 45.250 73.785 45.420 74.395 ;
        RECT 45.770 74.245 46.020 74.835 ;
        RECT 46.740 74.715 46.920 75.365 ;
        RECT 48.130 75.295 48.630 75.905 ;
        RECT 47.925 74.835 48.275 75.085 ;
        RECT 46.740 74.545 47.005 74.715 ;
        RECT 48.460 74.665 48.630 75.295 ;
        RECT 49.260 75.425 49.590 75.905 ;
        RECT 49.760 75.615 49.985 76.075 ;
        RECT 50.155 75.425 50.485 75.905 ;
        RECT 49.260 75.255 50.485 75.425 ;
        RECT 50.675 75.275 50.925 76.075 ;
        RECT 51.095 75.275 51.435 75.905 ;
        RECT 51.615 75.575 51.945 76.075 ;
        RECT 52.145 75.505 52.315 75.855 ;
        RECT 52.515 75.675 52.845 76.075 ;
        RECT 53.015 75.505 53.185 75.855 ;
        RECT 53.355 75.675 53.735 76.075 ;
        RECT 51.205 75.225 51.435 75.275 ;
        RECT 48.800 74.885 49.130 75.085 ;
        RECT 49.300 74.885 49.630 75.085 ;
        RECT 49.800 74.885 50.220 75.085 ;
        RECT 50.395 74.915 51.090 75.085 ;
        RECT 50.395 74.665 50.565 74.915 ;
        RECT 51.260 74.665 51.435 75.225 ;
        RECT 51.610 74.835 51.960 75.405 ;
        RECT 52.145 75.335 53.755 75.505 ;
        RECT 53.925 75.400 54.195 75.745 ;
        RECT 53.585 75.165 53.755 75.335 ;
        RECT 52.130 74.715 52.840 75.165 ;
        RECT 53.010 74.835 53.415 75.165 ;
        RECT 53.585 74.835 53.855 75.165 ;
        RECT 46.740 74.505 46.920 74.545 ;
        RECT 45.690 73.735 46.020 74.245 ;
        RECT 46.200 73.525 46.485 74.325 ;
        RECT 46.665 73.835 46.920 74.505 ;
        RECT 48.130 74.495 50.565 74.665 ;
        RECT 48.130 73.695 48.460 74.495 ;
        RECT 48.630 73.525 48.960 74.325 ;
        RECT 49.260 73.695 49.590 74.495 ;
        RECT 50.235 73.525 50.485 74.325 ;
        RECT 50.755 73.525 50.925 74.665 ;
        RECT 51.095 73.695 51.435 74.665 ;
        RECT 51.610 74.375 51.930 74.665 ;
        RECT 52.125 74.545 52.840 74.715 ;
        RECT 53.585 74.665 53.755 74.835 ;
        RECT 54.025 74.665 54.195 75.400 ;
        RECT 53.030 74.495 53.755 74.665 ;
        RECT 53.030 74.375 53.200 74.495 ;
        RECT 51.610 74.205 53.200 74.375 ;
        RECT 51.610 73.745 53.265 74.035 ;
        RECT 53.435 73.525 53.715 74.325 ;
        RECT 53.925 73.695 54.195 74.665 ;
        RECT 54.365 75.400 54.625 75.905 ;
        RECT 54.805 75.695 55.135 76.075 ;
        RECT 55.315 75.525 55.485 75.905 ;
        RECT 54.365 74.600 54.535 75.400 ;
        RECT 54.820 75.355 55.485 75.525 ;
        RECT 54.820 75.100 54.990 75.355 ;
        RECT 55.785 75.255 56.015 76.075 ;
        RECT 56.185 75.275 56.515 75.905 ;
        RECT 54.705 74.770 54.990 75.100 ;
        RECT 55.225 74.805 55.555 75.175 ;
        RECT 55.765 74.835 56.095 75.085 ;
        RECT 54.820 74.625 54.990 74.770 ;
        RECT 56.265 74.675 56.515 75.275 ;
        RECT 56.685 75.255 56.895 76.075 ;
        RECT 57.125 75.350 57.415 76.075 ;
        RECT 57.585 75.305 60.175 76.075 ;
        RECT 60.435 75.525 60.605 75.815 ;
        RECT 60.775 75.695 61.105 76.075 ;
        RECT 60.435 75.355 61.100 75.525 ;
        RECT 57.585 74.785 58.795 75.305 ;
        RECT 54.365 73.695 54.635 74.600 ;
        RECT 54.820 74.455 55.485 74.625 ;
        RECT 54.805 73.525 55.135 74.285 ;
        RECT 55.315 73.695 55.485 74.455 ;
        RECT 55.785 73.525 56.015 74.665 ;
        RECT 56.185 73.695 56.515 74.675 ;
        RECT 56.685 73.525 56.895 74.665 ;
        RECT 57.125 73.525 57.415 74.690 ;
        RECT 58.965 74.615 60.175 75.135 ;
        RECT 57.585 73.525 60.175 74.615 ;
        RECT 60.350 74.535 60.700 75.185 ;
        RECT 60.870 74.365 61.100 75.355 ;
        RECT 60.435 74.195 61.100 74.365 ;
        RECT 60.435 73.695 60.605 74.195 ;
        RECT 60.775 73.525 61.105 74.025 ;
        RECT 61.275 73.695 61.500 75.815 ;
        RECT 61.715 75.695 62.045 76.075 ;
        RECT 62.215 75.525 62.385 75.855 ;
        RECT 62.685 75.695 63.700 75.895 ;
        RECT 61.690 75.335 62.385 75.525 ;
        RECT 61.690 74.365 61.860 75.335 ;
        RECT 62.030 74.535 62.440 75.155 ;
        RECT 62.610 74.585 62.830 75.455 ;
        RECT 63.010 75.145 63.360 75.515 ;
        RECT 63.530 74.965 63.700 75.695 ;
        RECT 63.870 75.635 64.280 76.075 ;
        RECT 64.570 75.435 64.820 75.865 ;
        RECT 65.020 75.615 65.340 76.075 ;
        RECT 65.900 75.685 66.750 75.855 ;
        RECT 63.870 75.095 64.280 75.425 ;
        RECT 64.570 75.095 64.990 75.435 ;
        RECT 63.280 74.925 63.700 74.965 ;
        RECT 63.280 74.755 64.630 74.925 ;
        RECT 61.690 74.195 62.385 74.365 ;
        RECT 62.610 74.205 63.110 74.585 ;
        RECT 61.715 73.525 62.045 74.025 ;
        RECT 62.215 73.695 62.385 74.195 ;
        RECT 63.280 73.910 63.450 74.755 ;
        RECT 64.380 74.595 64.630 74.755 ;
        RECT 63.620 74.325 63.870 74.585 ;
        RECT 64.800 74.325 64.990 75.095 ;
        RECT 63.620 74.075 64.990 74.325 ;
        RECT 65.160 75.265 66.410 75.435 ;
        RECT 65.160 74.505 65.330 75.265 ;
        RECT 66.080 75.145 66.410 75.265 ;
        RECT 65.500 74.685 65.680 75.095 ;
        RECT 66.580 74.925 66.750 75.685 ;
        RECT 66.950 75.595 67.610 76.075 ;
        RECT 67.790 75.480 68.110 75.810 ;
        RECT 66.940 75.155 67.600 75.425 ;
        RECT 66.940 75.095 67.270 75.155 ;
        RECT 67.420 74.925 67.750 74.985 ;
        RECT 65.850 74.755 67.750 74.925 ;
        RECT 65.160 74.195 65.680 74.505 ;
        RECT 65.850 74.245 66.020 74.755 ;
        RECT 67.920 74.585 68.110 75.480 ;
        RECT 66.190 74.415 68.110 74.585 ;
        RECT 67.790 74.395 68.110 74.415 ;
        RECT 68.310 75.165 68.560 75.815 ;
        RECT 68.740 75.615 69.025 76.075 ;
        RECT 69.205 75.365 69.460 75.895 ;
        RECT 68.310 74.835 69.110 75.165 ;
        RECT 65.850 74.075 67.060 74.245 ;
        RECT 62.620 73.740 63.450 73.910 ;
        RECT 63.690 73.525 64.070 73.905 ;
        RECT 64.250 73.785 64.420 74.075 ;
        RECT 65.850 73.995 66.020 74.075 ;
        RECT 64.590 73.525 64.920 73.905 ;
        RECT 65.390 73.745 66.020 73.995 ;
        RECT 66.200 73.525 66.620 73.905 ;
        RECT 66.820 73.785 67.060 74.075 ;
        RECT 67.290 73.525 67.620 74.215 ;
        RECT 67.790 73.785 67.960 74.395 ;
        RECT 68.310 74.245 68.560 74.835 ;
        RECT 69.280 74.505 69.460 75.365 ;
        RECT 69.205 74.375 69.460 74.505 ;
        RECT 70.010 75.335 70.265 75.905 ;
        RECT 70.435 75.675 70.765 76.075 ;
        RECT 71.190 75.540 71.720 75.905 ;
        RECT 71.190 75.505 71.365 75.540 ;
        RECT 70.435 75.335 71.365 75.505 ;
        RECT 70.010 74.665 70.180 75.335 ;
        RECT 70.435 75.165 70.605 75.335 ;
        RECT 70.350 74.835 70.605 75.165 ;
        RECT 70.830 74.835 71.025 75.165 ;
        RECT 68.230 73.735 68.560 74.245 ;
        RECT 68.740 73.525 69.025 74.325 ;
        RECT 69.205 74.205 69.545 74.375 ;
        RECT 69.205 73.835 69.460 74.205 ;
        RECT 70.010 73.695 70.345 74.665 ;
        RECT 70.515 73.525 70.685 74.665 ;
        RECT 70.855 73.865 71.025 74.835 ;
        RECT 71.195 74.205 71.365 75.335 ;
        RECT 71.535 74.545 71.705 75.345 ;
        RECT 71.910 75.055 72.185 75.905 ;
        RECT 71.905 74.885 72.185 75.055 ;
        RECT 71.910 74.745 72.185 74.885 ;
        RECT 72.355 74.545 72.545 75.905 ;
        RECT 72.725 75.540 73.235 76.075 ;
        RECT 73.455 75.265 73.700 75.870 ;
        RECT 75.340 75.265 75.585 75.870 ;
        RECT 75.805 75.540 76.315 76.075 ;
        RECT 72.745 75.095 73.975 75.265 ;
        RECT 71.535 74.375 72.545 74.545 ;
        RECT 72.715 74.530 73.465 74.720 ;
        RECT 71.195 74.035 72.320 74.205 ;
        RECT 72.715 73.865 72.885 74.530 ;
        RECT 73.635 74.285 73.975 75.095 ;
        RECT 70.855 73.695 72.885 73.865 ;
        RECT 73.055 73.525 73.225 74.285 ;
        RECT 73.460 73.875 73.975 74.285 ;
        RECT 75.065 75.095 76.295 75.265 ;
        RECT 75.065 74.285 75.405 75.095 ;
        RECT 75.575 74.530 76.325 74.720 ;
        RECT 75.065 73.875 75.580 74.285 ;
        RECT 75.815 73.525 75.985 74.285 ;
        RECT 76.155 73.865 76.325 74.530 ;
        RECT 76.495 74.545 76.685 75.905 ;
        RECT 76.855 75.055 77.130 75.905 ;
        RECT 77.320 75.540 77.850 75.905 ;
        RECT 78.275 75.675 78.605 76.075 ;
        RECT 77.675 75.505 77.850 75.540 ;
        RECT 76.855 74.885 77.135 75.055 ;
        RECT 76.855 74.745 77.130 74.885 ;
        RECT 77.335 74.545 77.505 75.345 ;
        RECT 76.495 74.375 77.505 74.545 ;
        RECT 77.675 75.335 78.605 75.505 ;
        RECT 78.775 75.335 79.030 75.905 ;
        RECT 77.675 74.205 77.845 75.335 ;
        RECT 78.435 75.165 78.605 75.335 ;
        RECT 76.720 74.035 77.845 74.205 ;
        RECT 78.015 74.835 78.210 75.165 ;
        RECT 78.435 74.835 78.690 75.165 ;
        RECT 78.015 73.865 78.185 74.835 ;
        RECT 78.860 74.665 79.030 75.335 ;
        RECT 76.155 73.695 78.185 73.865 ;
        RECT 78.355 73.525 78.525 74.665 ;
        RECT 78.695 73.695 79.030 74.665 ;
        RECT 79.205 75.275 79.545 75.905 ;
        RECT 79.715 75.275 79.965 76.075 ;
        RECT 80.155 75.425 80.485 75.905 ;
        RECT 80.655 75.615 80.880 76.075 ;
        RECT 81.050 75.425 81.380 75.905 ;
        RECT 79.205 74.665 79.380 75.275 ;
        RECT 80.155 75.255 81.380 75.425 ;
        RECT 82.010 75.295 82.510 75.905 ;
        RECT 82.885 75.350 83.175 76.075 ;
        RECT 79.550 74.915 80.245 75.085 ;
        RECT 80.075 74.665 80.245 74.915 ;
        RECT 80.420 74.885 80.840 75.085 ;
        RECT 81.010 74.885 81.340 75.085 ;
        RECT 81.510 74.885 81.840 75.085 ;
        RECT 82.010 74.665 82.180 75.295 ;
        RECT 83.405 75.255 83.615 76.075 ;
        RECT 83.785 75.275 84.115 75.905 ;
        RECT 82.365 74.835 82.715 75.085 ;
        RECT 79.205 73.695 79.545 74.665 ;
        RECT 79.715 73.525 79.885 74.665 ;
        RECT 80.075 74.495 82.510 74.665 ;
        RECT 80.155 73.525 80.405 74.325 ;
        RECT 81.050 73.695 81.380 74.495 ;
        RECT 81.680 73.525 82.010 74.325 ;
        RECT 82.180 73.695 82.510 74.495 ;
        RECT 82.885 73.525 83.175 74.690 ;
        RECT 83.785 74.675 84.035 75.275 ;
        RECT 84.285 75.255 84.515 76.075 ;
        RECT 84.725 75.305 86.395 76.075 ;
        RECT 86.575 75.575 86.905 76.075 ;
        RECT 87.105 75.505 87.275 75.855 ;
        RECT 87.475 75.675 87.805 76.075 ;
        RECT 87.975 75.505 88.145 75.855 ;
        RECT 88.315 75.675 88.695 76.075 ;
        RECT 84.205 74.835 84.535 75.085 ;
        RECT 84.725 74.785 85.475 75.305 ;
        RECT 83.405 73.525 83.615 74.665 ;
        RECT 83.785 73.695 84.115 74.675 ;
        RECT 84.285 73.525 84.515 74.665 ;
        RECT 85.645 74.615 86.395 75.135 ;
        RECT 86.570 74.835 86.920 75.405 ;
        RECT 87.105 75.335 88.715 75.505 ;
        RECT 88.885 75.400 89.155 75.745 ;
        RECT 88.545 75.165 88.715 75.335 ;
        RECT 87.090 74.715 87.800 75.165 ;
        RECT 87.970 74.835 88.375 75.165 ;
        RECT 88.545 74.835 88.815 75.165 ;
        RECT 84.725 73.525 86.395 74.615 ;
        RECT 86.570 74.375 86.890 74.665 ;
        RECT 87.085 74.545 87.800 74.715 ;
        RECT 88.545 74.665 88.715 74.835 ;
        RECT 88.985 74.665 89.155 75.400 ;
        RECT 89.325 75.305 90.995 76.075 ;
        RECT 91.175 75.575 91.505 76.075 ;
        RECT 91.705 75.505 91.875 75.855 ;
        RECT 92.075 75.675 92.405 76.075 ;
        RECT 92.575 75.505 92.745 75.855 ;
        RECT 92.915 75.675 93.295 76.075 ;
        RECT 89.325 74.785 90.075 75.305 ;
        RECT 87.990 74.495 88.715 74.665 ;
        RECT 87.990 74.375 88.160 74.495 ;
        RECT 86.570 74.205 88.160 74.375 ;
        RECT 86.570 73.745 88.225 74.035 ;
        RECT 88.395 73.525 88.675 74.325 ;
        RECT 88.885 73.695 89.155 74.665 ;
        RECT 90.245 74.615 90.995 75.135 ;
        RECT 91.170 74.835 91.520 75.405 ;
        RECT 91.705 75.335 93.315 75.505 ;
        RECT 93.485 75.400 93.755 75.745 ;
        RECT 93.935 75.575 94.265 76.075 ;
        RECT 94.465 75.505 94.635 75.855 ;
        RECT 94.835 75.675 95.165 76.075 ;
        RECT 95.335 75.505 95.505 75.855 ;
        RECT 95.675 75.675 96.055 76.075 ;
        RECT 93.145 75.165 93.315 75.335 ;
        RECT 89.325 73.525 90.995 74.615 ;
        RECT 91.170 74.375 91.490 74.665 ;
        RECT 91.690 74.545 92.400 75.165 ;
        RECT 92.570 74.835 92.975 75.165 ;
        RECT 93.145 74.835 93.415 75.165 ;
        RECT 93.145 74.665 93.315 74.835 ;
        RECT 93.585 74.665 93.755 75.400 ;
        RECT 93.930 74.835 94.280 75.405 ;
        RECT 94.465 75.335 96.075 75.505 ;
        RECT 96.245 75.400 96.515 75.745 ;
        RECT 96.695 75.575 97.025 76.075 ;
        RECT 97.225 75.505 97.395 75.855 ;
        RECT 97.595 75.675 97.925 76.075 ;
        RECT 98.095 75.505 98.265 75.855 ;
        RECT 98.435 75.675 98.815 76.075 ;
        RECT 95.905 75.165 96.075 75.335 ;
        RECT 94.450 74.715 95.160 75.165 ;
        RECT 95.330 74.835 95.735 75.165 ;
        RECT 95.905 74.835 96.175 75.165 ;
        RECT 92.590 74.495 93.315 74.665 ;
        RECT 92.590 74.375 92.760 74.495 ;
        RECT 91.170 74.205 92.760 74.375 ;
        RECT 91.170 73.745 92.825 74.035 ;
        RECT 92.995 73.525 93.275 74.325 ;
        RECT 93.485 73.695 93.755 74.665 ;
        RECT 93.930 74.375 94.250 74.665 ;
        RECT 94.445 74.545 95.160 74.715 ;
        RECT 95.905 74.665 96.075 74.835 ;
        RECT 96.345 74.665 96.515 75.400 ;
        RECT 96.690 74.835 97.040 75.405 ;
        RECT 97.225 75.335 98.835 75.505 ;
        RECT 99.005 75.400 99.275 75.745 ;
        RECT 98.665 75.165 98.835 75.335 ;
        RECT 97.210 74.715 97.920 75.165 ;
        RECT 98.090 74.835 98.495 75.165 ;
        RECT 98.665 74.835 98.935 75.165 ;
        RECT 95.350 74.495 96.075 74.665 ;
        RECT 95.350 74.375 95.520 74.495 ;
        RECT 93.930 74.205 95.520 74.375 ;
        RECT 93.930 73.745 95.585 74.035 ;
        RECT 95.755 73.525 96.035 74.325 ;
        RECT 96.245 73.695 96.515 74.665 ;
        RECT 96.690 74.375 97.010 74.665 ;
        RECT 97.205 74.545 97.920 74.715 ;
        RECT 98.665 74.665 98.835 74.835 ;
        RECT 99.105 74.665 99.275 75.400 ;
        RECT 99.445 75.305 102.955 76.075 ;
        RECT 99.445 74.785 101.095 75.305 ;
        RECT 104.320 75.265 104.565 75.870 ;
        RECT 104.785 75.540 105.295 76.075 ;
        RECT 98.110 74.495 98.835 74.665 ;
        RECT 98.110 74.375 98.280 74.495 ;
        RECT 96.690 74.205 98.280 74.375 ;
        RECT 96.690 73.745 98.345 74.035 ;
        RECT 98.515 73.525 98.795 74.325 ;
        RECT 99.005 73.695 99.275 74.665 ;
        RECT 101.265 74.615 102.955 75.135 ;
        RECT 99.445 73.525 102.955 74.615 ;
        RECT 104.045 75.095 105.275 75.265 ;
        RECT 104.045 74.285 104.385 75.095 ;
        RECT 104.555 74.530 105.305 74.720 ;
        RECT 104.045 73.875 104.560 74.285 ;
        RECT 104.795 73.525 104.965 74.285 ;
        RECT 105.135 73.865 105.305 74.530 ;
        RECT 105.475 74.545 105.665 75.905 ;
        RECT 105.835 75.735 106.110 75.905 ;
        RECT 105.835 75.565 106.115 75.735 ;
        RECT 105.835 74.745 106.110 75.565 ;
        RECT 106.300 75.540 106.830 75.905 ;
        RECT 107.255 75.675 107.585 76.075 ;
        RECT 106.655 75.505 106.830 75.540 ;
        RECT 106.315 74.545 106.485 75.345 ;
        RECT 105.475 74.375 106.485 74.545 ;
        RECT 106.655 75.335 107.585 75.505 ;
        RECT 107.755 75.335 108.010 75.905 ;
        RECT 108.645 75.350 108.935 76.075 ;
        RECT 106.655 74.205 106.825 75.335 ;
        RECT 107.415 75.165 107.585 75.335 ;
        RECT 105.700 74.035 106.825 74.205 ;
        RECT 106.995 74.835 107.190 75.165 ;
        RECT 107.415 74.835 107.670 75.165 ;
        RECT 106.995 73.865 107.165 74.835 ;
        RECT 107.840 74.665 108.010 75.335 ;
        RECT 109.105 75.305 111.695 76.075 ;
        RECT 112.325 75.325 113.535 76.075 ;
        RECT 109.105 74.785 110.315 75.305 ;
        RECT 105.135 73.695 107.165 73.865 ;
        RECT 107.335 73.525 107.505 74.665 ;
        RECT 107.675 73.695 108.010 74.665 ;
        RECT 108.645 73.525 108.935 74.690 ;
        RECT 110.485 74.615 111.695 75.135 ;
        RECT 109.105 73.525 111.695 74.615 ;
        RECT 112.325 74.615 112.845 75.155 ;
        RECT 113.015 74.785 113.535 75.325 ;
        RECT 112.325 73.525 113.535 74.615 ;
        RECT 5.520 73.355 113.620 73.525 ;
        RECT 5.605 72.265 6.815 73.355 ;
        RECT 6.985 72.265 10.495 73.355 ;
        RECT 10.665 72.265 11.875 73.355 ;
        RECT 5.605 71.555 6.125 72.095 ;
        RECT 6.295 71.725 6.815 72.265 ;
        RECT 6.985 71.575 8.635 72.095 ;
        RECT 8.805 71.745 10.495 72.265 ;
        RECT 5.605 70.805 6.815 71.555 ;
        RECT 6.985 70.805 10.495 71.575 ;
        RECT 10.665 71.555 11.185 72.095 ;
        RECT 11.355 71.725 11.875 72.265 ;
        RECT 12.105 72.215 12.315 73.355 ;
        RECT 12.485 72.205 12.815 73.185 ;
        RECT 12.985 72.215 13.215 73.355 ;
        RECT 13.425 72.265 16.935 73.355 ;
        RECT 17.105 72.265 18.315 73.355 ;
        RECT 10.665 70.805 11.875 71.555 ;
        RECT 12.105 70.805 12.315 71.625 ;
        RECT 12.485 71.605 12.735 72.205 ;
        RECT 12.905 71.795 13.235 72.045 ;
        RECT 12.485 70.975 12.815 71.605 ;
        RECT 12.985 70.805 13.215 71.625 ;
        RECT 13.425 71.575 15.075 72.095 ;
        RECT 15.245 71.745 16.935 72.265 ;
        RECT 13.425 70.805 16.935 71.575 ;
        RECT 17.105 71.555 17.625 72.095 ;
        RECT 17.795 71.725 18.315 72.265 ;
        RECT 18.485 72.190 18.775 73.355 ;
        RECT 18.945 72.265 20.615 73.355 ;
        RECT 18.945 71.575 19.695 72.095 ;
        RECT 19.865 71.745 20.615 72.265 ;
        RECT 20.785 72.215 21.125 73.185 ;
        RECT 21.295 72.215 21.465 73.355 ;
        RECT 21.735 72.555 21.985 73.355 ;
        RECT 22.630 72.385 22.960 73.185 ;
        RECT 23.260 72.555 23.590 73.355 ;
        RECT 23.760 72.385 24.090 73.185 ;
        RECT 21.655 72.215 24.090 72.385 ;
        RECT 24.670 72.385 25.000 73.185 ;
        RECT 25.170 72.555 25.500 73.355 ;
        RECT 25.800 72.385 26.130 73.185 ;
        RECT 26.775 72.555 27.025 73.355 ;
        RECT 24.670 72.215 27.105 72.385 ;
        RECT 27.295 72.215 27.465 73.355 ;
        RECT 27.635 72.215 27.975 73.185 ;
        RECT 28.150 72.845 29.805 73.135 ;
        RECT 28.150 72.505 29.740 72.675 ;
        RECT 29.975 72.555 30.255 73.355 ;
        RECT 28.150 72.215 28.470 72.505 ;
        RECT 29.570 72.385 29.740 72.505 ;
        RECT 20.785 71.605 20.960 72.215 ;
        RECT 21.655 71.965 21.825 72.215 ;
        RECT 21.130 71.795 21.825 71.965 ;
        RECT 21.995 71.825 22.420 71.995 ;
        RECT 22.000 71.795 22.420 71.825 ;
        RECT 22.590 71.795 22.920 71.995 ;
        RECT 23.090 71.795 23.420 71.995 ;
        RECT 17.105 70.805 18.315 71.555 ;
        RECT 18.485 70.805 18.775 71.530 ;
        RECT 18.945 70.805 20.615 71.575 ;
        RECT 20.785 70.975 21.125 71.605 ;
        RECT 21.295 70.805 21.545 71.605 ;
        RECT 21.735 71.455 22.960 71.625 ;
        RECT 21.735 70.975 22.065 71.455 ;
        RECT 22.235 70.805 22.460 71.265 ;
        RECT 22.630 70.975 22.960 71.455 ;
        RECT 23.590 71.585 23.760 72.215 ;
        RECT 23.945 71.795 24.295 72.045 ;
        RECT 24.465 71.795 24.815 72.045 ;
        RECT 25.000 71.585 25.170 72.215 ;
        RECT 25.340 71.795 25.670 71.995 ;
        RECT 25.840 71.795 26.170 71.995 ;
        RECT 26.340 71.795 26.760 71.995 ;
        RECT 26.935 71.965 27.105 72.215 ;
        RECT 26.935 71.795 27.630 71.965 ;
        RECT 27.800 71.655 27.975 72.215 ;
        RECT 23.590 70.975 24.090 71.585 ;
        RECT 24.670 70.975 25.170 71.585 ;
        RECT 25.800 71.455 27.025 71.625 ;
        RECT 27.745 71.605 27.975 71.655 ;
        RECT 25.800 70.975 26.130 71.455 ;
        RECT 26.300 70.805 26.525 71.265 ;
        RECT 26.695 70.975 27.025 71.455 ;
        RECT 27.215 70.805 27.465 71.605 ;
        RECT 27.635 70.975 27.975 71.605 ;
        RECT 28.150 71.475 28.500 72.045 ;
        RECT 28.670 71.715 29.380 72.335 ;
        RECT 29.570 72.215 30.295 72.385 ;
        RECT 30.465 72.215 30.735 73.185 ;
        RECT 31.830 72.845 33.485 73.135 ;
        RECT 31.830 72.505 33.420 72.675 ;
        RECT 33.655 72.555 33.935 73.355 ;
        RECT 31.830 72.215 32.150 72.505 ;
        RECT 33.250 72.385 33.420 72.505 ;
        RECT 30.125 72.045 30.295 72.215 ;
        RECT 29.550 71.715 29.955 72.045 ;
        RECT 30.125 71.715 30.395 72.045 ;
        RECT 30.125 71.545 30.295 71.715 ;
        RECT 28.685 71.375 30.295 71.545 ;
        RECT 30.565 71.480 30.735 72.215 ;
        RECT 32.345 72.165 33.060 72.335 ;
        RECT 33.250 72.215 33.975 72.385 ;
        RECT 34.145 72.215 34.415 73.185 ;
        RECT 34.675 72.685 34.845 73.185 ;
        RECT 35.015 72.855 35.345 73.355 ;
        RECT 34.675 72.515 35.340 72.685 ;
        RECT 28.155 70.805 28.485 71.305 ;
        RECT 28.685 71.025 28.855 71.375 ;
        RECT 29.055 70.805 29.385 71.205 ;
        RECT 29.555 71.025 29.725 71.375 ;
        RECT 29.895 70.805 30.275 71.205 ;
        RECT 30.465 71.135 30.735 71.480 ;
        RECT 31.830 71.475 32.180 72.045 ;
        RECT 32.350 71.715 33.060 72.165 ;
        RECT 33.805 72.045 33.975 72.215 ;
        RECT 33.230 71.715 33.635 72.045 ;
        RECT 33.805 71.715 34.075 72.045 ;
        RECT 33.805 71.545 33.975 71.715 ;
        RECT 32.365 71.375 33.975 71.545 ;
        RECT 34.245 71.480 34.415 72.215 ;
        RECT 34.590 71.695 34.940 72.345 ;
        RECT 35.110 71.525 35.340 72.515 ;
        RECT 31.835 70.805 32.165 71.305 ;
        RECT 32.365 71.025 32.535 71.375 ;
        RECT 32.735 70.805 33.065 71.205 ;
        RECT 33.235 71.025 33.405 71.375 ;
        RECT 33.575 70.805 33.955 71.205 ;
        RECT 34.145 71.135 34.415 71.480 ;
        RECT 34.675 71.355 35.340 71.525 ;
        RECT 34.675 71.065 34.845 71.355 ;
        RECT 35.015 70.805 35.345 71.185 ;
        RECT 35.515 71.065 35.740 73.185 ;
        RECT 35.955 72.855 36.285 73.355 ;
        RECT 36.455 72.685 36.625 73.185 ;
        RECT 36.860 72.970 37.690 73.140 ;
        RECT 37.930 72.975 38.310 73.355 ;
        RECT 35.930 72.515 36.625 72.685 ;
        RECT 35.930 71.545 36.100 72.515 ;
        RECT 36.270 71.725 36.680 72.345 ;
        RECT 36.850 72.295 37.350 72.675 ;
        RECT 35.930 71.355 36.625 71.545 ;
        RECT 36.850 71.425 37.070 72.295 ;
        RECT 37.520 72.125 37.690 72.970 ;
        RECT 38.490 72.805 38.660 73.095 ;
        RECT 38.830 72.975 39.160 73.355 ;
        RECT 39.630 72.885 40.260 73.135 ;
        RECT 40.440 72.975 40.860 73.355 ;
        RECT 40.090 72.805 40.260 72.885 ;
        RECT 41.060 72.805 41.300 73.095 ;
        RECT 37.860 72.555 39.230 72.805 ;
        RECT 37.860 72.295 38.110 72.555 ;
        RECT 38.620 72.125 38.870 72.285 ;
        RECT 37.520 71.955 38.870 72.125 ;
        RECT 37.520 71.915 37.940 71.955 ;
        RECT 37.250 71.365 37.600 71.735 ;
        RECT 35.955 70.805 36.285 71.185 ;
        RECT 36.455 71.025 36.625 71.355 ;
        RECT 37.770 71.185 37.940 71.915 ;
        RECT 39.040 71.785 39.230 72.555 ;
        RECT 38.110 71.455 38.520 71.785 ;
        RECT 38.810 71.445 39.230 71.785 ;
        RECT 39.400 72.375 39.920 72.685 ;
        RECT 40.090 72.635 41.300 72.805 ;
        RECT 41.530 72.665 41.860 73.355 ;
        RECT 39.400 71.615 39.570 72.375 ;
        RECT 39.740 71.785 39.920 72.195 ;
        RECT 40.090 72.125 40.260 72.635 ;
        RECT 42.030 72.485 42.200 73.095 ;
        RECT 42.470 72.635 42.800 73.145 ;
        RECT 42.030 72.465 42.350 72.485 ;
        RECT 40.430 72.295 42.350 72.465 ;
        RECT 40.090 71.955 41.990 72.125 ;
        RECT 40.320 71.615 40.650 71.735 ;
        RECT 39.400 71.445 40.650 71.615 ;
        RECT 36.925 70.985 37.940 71.185 ;
        RECT 38.110 70.805 38.520 71.245 ;
        RECT 38.810 71.015 39.060 71.445 ;
        RECT 39.260 70.805 39.580 71.265 ;
        RECT 40.820 71.195 40.990 71.955 ;
        RECT 41.660 71.895 41.990 71.955 ;
        RECT 41.180 71.725 41.510 71.785 ;
        RECT 41.180 71.455 41.840 71.725 ;
        RECT 42.160 71.400 42.350 72.295 ;
        RECT 40.140 71.025 40.990 71.195 ;
        RECT 41.190 70.805 41.850 71.285 ;
        RECT 42.030 71.070 42.350 71.400 ;
        RECT 42.550 72.045 42.800 72.635 ;
        RECT 42.980 72.555 43.265 73.355 ;
        RECT 43.445 72.375 43.700 73.045 ;
        RECT 42.550 71.715 43.350 72.045 ;
        RECT 42.550 71.065 42.800 71.715 ;
        RECT 43.520 71.655 43.700 72.375 ;
        RECT 44.245 72.190 44.535 73.355 ;
        RECT 44.710 72.215 45.045 73.185 ;
        RECT 45.215 72.215 45.385 73.355 ;
        RECT 45.555 73.015 47.585 73.185 ;
        RECT 43.520 71.515 43.785 71.655 ;
        RECT 44.710 71.545 44.880 72.215 ;
        RECT 45.555 72.045 45.725 73.015 ;
        RECT 45.050 71.715 45.305 72.045 ;
        RECT 45.530 71.715 45.725 72.045 ;
        RECT 45.895 72.675 47.020 72.845 ;
        RECT 45.135 71.545 45.305 71.715 ;
        RECT 45.895 71.545 46.065 72.675 ;
        RECT 43.445 71.485 43.785 71.515 ;
        RECT 42.980 70.805 43.265 71.265 ;
        RECT 43.445 70.985 43.700 71.485 ;
        RECT 44.245 70.805 44.535 71.530 ;
        RECT 44.710 70.975 44.965 71.545 ;
        RECT 45.135 71.375 46.065 71.545 ;
        RECT 46.235 72.335 47.245 72.505 ;
        RECT 46.235 71.535 46.405 72.335 ;
        RECT 46.610 71.995 46.885 72.135 ;
        RECT 46.605 71.825 46.885 71.995 ;
        RECT 45.890 71.340 46.065 71.375 ;
        RECT 45.135 70.805 45.465 71.205 ;
        RECT 45.890 70.975 46.420 71.340 ;
        RECT 46.610 70.975 46.885 71.825 ;
        RECT 47.055 70.975 47.245 72.335 ;
        RECT 47.415 72.350 47.585 73.015 ;
        RECT 47.755 72.595 47.925 73.355 ;
        RECT 48.160 72.595 48.675 73.005 ;
        RECT 47.415 72.160 48.165 72.350 ;
        RECT 48.335 71.785 48.675 72.595 ;
        RECT 49.050 72.385 49.380 73.185 ;
        RECT 49.550 72.555 49.880 73.355 ;
        RECT 50.180 72.385 50.510 73.185 ;
        RECT 51.155 72.555 51.405 73.355 ;
        RECT 49.050 72.215 51.485 72.385 ;
        RECT 51.675 72.215 51.845 73.355 ;
        RECT 52.015 72.215 52.355 73.185 ;
        RECT 52.525 72.265 55.115 73.355 ;
        RECT 48.845 71.795 49.195 72.045 ;
        RECT 47.445 71.615 48.675 71.785 ;
        RECT 47.425 70.805 47.935 71.340 ;
        RECT 48.155 71.010 48.400 71.615 ;
        RECT 49.380 71.585 49.550 72.215 ;
        RECT 49.720 71.795 50.050 71.995 ;
        RECT 50.220 71.795 50.550 71.995 ;
        RECT 50.720 71.795 51.140 71.995 ;
        RECT 51.315 71.965 51.485 72.215 ;
        RECT 51.315 71.795 52.010 71.965 ;
        RECT 49.050 70.975 49.550 71.585 ;
        RECT 50.180 71.455 51.405 71.625 ;
        RECT 52.180 71.605 52.355 72.215 ;
        RECT 50.180 70.975 50.510 71.455 ;
        RECT 50.680 70.805 50.905 71.265 ;
        RECT 51.075 70.975 51.405 71.455 ;
        RECT 51.595 70.805 51.845 71.605 ;
        RECT 52.015 70.975 52.355 71.605 ;
        RECT 52.525 71.575 53.735 72.095 ;
        RECT 53.905 71.745 55.115 72.265 ;
        RECT 55.745 72.385 56.055 73.185 ;
        RECT 56.225 72.555 56.535 73.355 ;
        RECT 56.705 72.725 56.965 73.185 ;
        RECT 57.135 72.895 57.390 73.355 ;
        RECT 57.565 72.725 57.825 73.185 ;
        RECT 56.705 72.555 57.825 72.725 ;
        RECT 55.745 72.215 56.775 72.385 ;
        RECT 52.525 70.805 55.115 71.575 ;
        RECT 55.745 71.305 55.915 72.215 ;
        RECT 56.085 71.475 56.435 72.045 ;
        RECT 56.605 71.965 56.775 72.215 ;
        RECT 57.565 72.305 57.825 72.555 ;
        RECT 57.995 72.485 58.280 73.355 ;
        RECT 58.710 72.385 59.040 73.185 ;
        RECT 59.210 72.555 59.540 73.355 ;
        RECT 59.840 72.385 60.170 73.185 ;
        RECT 60.815 72.555 61.065 73.355 ;
        RECT 57.565 72.135 58.320 72.305 ;
        RECT 58.710 72.215 61.145 72.385 ;
        RECT 61.335 72.215 61.505 73.355 ;
        RECT 61.675 72.215 62.015 73.185 ;
        RECT 62.390 72.385 62.720 73.185 ;
        RECT 62.890 72.555 63.220 73.355 ;
        RECT 63.520 72.385 63.850 73.185 ;
        RECT 64.495 72.555 64.745 73.355 ;
        RECT 62.390 72.215 64.825 72.385 ;
        RECT 65.015 72.215 65.185 73.355 ;
        RECT 65.355 72.215 65.695 73.185 ;
        RECT 66.070 72.385 66.400 73.185 ;
        RECT 66.570 72.555 66.900 73.355 ;
        RECT 67.200 72.385 67.530 73.185 ;
        RECT 68.175 72.555 68.425 73.355 ;
        RECT 66.070 72.215 68.505 72.385 ;
        RECT 68.695 72.215 68.865 73.355 ;
        RECT 69.035 72.215 69.375 73.185 ;
        RECT 56.605 71.795 57.745 71.965 ;
        RECT 57.915 71.625 58.320 72.135 ;
        RECT 58.505 71.795 58.855 72.045 ;
        RECT 56.670 71.455 58.320 71.625 ;
        RECT 59.040 71.585 59.210 72.215 ;
        RECT 59.380 71.795 59.710 71.995 ;
        RECT 59.880 71.795 60.210 71.995 ;
        RECT 60.380 71.795 60.800 71.995 ;
        RECT 60.975 71.965 61.145 72.215 ;
        RECT 60.975 71.795 61.670 71.965 ;
        RECT 55.745 70.975 56.045 71.305 ;
        RECT 56.215 70.805 56.490 71.285 ;
        RECT 56.670 71.065 56.965 71.455 ;
        RECT 57.135 70.805 57.390 71.285 ;
        RECT 57.565 71.065 57.825 71.455 ;
        RECT 57.995 70.805 58.275 71.285 ;
        RECT 58.710 70.975 59.210 71.585 ;
        RECT 59.840 71.455 61.065 71.625 ;
        RECT 61.840 71.605 62.015 72.215 ;
        RECT 62.185 71.795 62.535 72.045 ;
        RECT 59.840 70.975 60.170 71.455 ;
        RECT 60.340 70.805 60.565 71.265 ;
        RECT 60.735 70.975 61.065 71.455 ;
        RECT 61.255 70.805 61.505 71.605 ;
        RECT 61.675 70.975 62.015 71.605 ;
        RECT 62.720 71.585 62.890 72.215 ;
        RECT 63.060 71.795 63.390 71.995 ;
        RECT 63.560 71.795 63.890 71.995 ;
        RECT 64.060 71.795 64.480 71.995 ;
        RECT 64.655 71.965 64.825 72.215 ;
        RECT 64.655 71.795 65.350 71.965 ;
        RECT 62.390 70.975 62.890 71.585 ;
        RECT 63.520 71.455 64.745 71.625 ;
        RECT 65.520 71.605 65.695 72.215 ;
        RECT 65.865 71.795 66.215 72.045 ;
        RECT 63.520 70.975 63.850 71.455 ;
        RECT 64.020 70.805 64.245 71.265 ;
        RECT 64.415 70.975 64.745 71.455 ;
        RECT 64.935 70.805 65.185 71.605 ;
        RECT 65.355 70.975 65.695 71.605 ;
        RECT 66.400 71.585 66.570 72.215 ;
        RECT 66.740 71.795 67.070 71.995 ;
        RECT 67.240 71.795 67.570 71.995 ;
        RECT 67.740 71.795 68.160 71.995 ;
        RECT 68.335 71.965 68.505 72.215 ;
        RECT 69.145 72.165 69.375 72.215 ;
        RECT 70.005 72.190 70.295 73.355 ;
        RECT 70.465 72.280 70.735 73.185 ;
        RECT 70.905 72.595 71.235 73.355 ;
        RECT 71.415 72.425 71.585 73.185 ;
        RECT 68.335 71.795 69.030 71.965 ;
        RECT 66.070 70.975 66.570 71.585 ;
        RECT 67.200 71.455 68.425 71.625 ;
        RECT 69.200 71.605 69.375 72.165 ;
        RECT 67.200 70.975 67.530 71.455 ;
        RECT 67.700 70.805 67.925 71.265 ;
        RECT 68.095 70.975 68.425 71.455 ;
        RECT 68.615 70.805 68.865 71.605 ;
        RECT 69.035 70.975 69.375 71.605 ;
        RECT 70.005 70.805 70.295 71.530 ;
        RECT 70.465 71.480 70.635 72.280 ;
        RECT 70.920 72.255 71.585 72.425 ;
        RECT 72.970 72.385 73.300 73.185 ;
        RECT 73.470 72.555 73.800 73.355 ;
        RECT 74.100 72.385 74.430 73.185 ;
        RECT 75.075 72.555 75.325 73.355 ;
        RECT 70.920 72.110 71.090 72.255 ;
        RECT 72.970 72.215 75.405 72.385 ;
        RECT 75.595 72.215 75.765 73.355 ;
        RECT 75.935 72.215 76.275 73.185 ;
        RECT 76.995 72.685 77.165 73.185 ;
        RECT 77.335 72.855 77.665 73.355 ;
        RECT 76.995 72.515 77.660 72.685 ;
        RECT 70.805 71.780 71.090 72.110 ;
        RECT 70.920 71.525 71.090 71.780 ;
        RECT 71.325 71.705 71.655 72.075 ;
        RECT 72.765 71.795 73.115 72.045 ;
        RECT 73.300 71.585 73.470 72.215 ;
        RECT 73.640 71.795 73.970 71.995 ;
        RECT 74.140 71.795 74.470 71.995 ;
        RECT 74.640 71.795 75.060 71.995 ;
        RECT 75.235 71.965 75.405 72.215 ;
        RECT 75.235 71.795 75.930 71.965 ;
        RECT 70.465 70.975 70.725 71.480 ;
        RECT 70.920 71.355 71.585 71.525 ;
        RECT 70.905 70.805 71.235 71.185 ;
        RECT 71.415 70.975 71.585 71.355 ;
        RECT 72.970 70.975 73.470 71.585 ;
        RECT 74.100 71.455 75.325 71.625 ;
        RECT 76.100 71.605 76.275 72.215 ;
        RECT 76.910 71.695 77.260 72.345 ;
        RECT 74.100 70.975 74.430 71.455 ;
        RECT 74.600 70.805 74.825 71.265 ;
        RECT 74.995 70.975 75.325 71.455 ;
        RECT 75.515 70.805 75.765 71.605 ;
        RECT 75.935 70.975 76.275 71.605 ;
        RECT 77.430 71.525 77.660 72.515 ;
        RECT 76.995 71.355 77.660 71.525 ;
        RECT 76.995 71.065 77.165 71.355 ;
        RECT 77.335 70.805 77.665 71.185 ;
        RECT 77.835 71.065 78.060 73.185 ;
        RECT 78.275 72.855 78.605 73.355 ;
        RECT 78.775 72.685 78.945 73.185 ;
        RECT 79.180 72.970 80.010 73.140 ;
        RECT 80.250 72.975 80.630 73.355 ;
        RECT 78.250 72.515 78.945 72.685 ;
        RECT 78.250 71.545 78.420 72.515 ;
        RECT 78.590 71.725 79.000 72.345 ;
        RECT 79.170 72.295 79.670 72.675 ;
        RECT 78.250 71.355 78.945 71.545 ;
        RECT 79.170 71.425 79.390 72.295 ;
        RECT 79.840 72.125 80.010 72.970 ;
        RECT 80.810 72.805 80.980 73.095 ;
        RECT 81.150 72.975 81.480 73.355 ;
        RECT 81.950 72.885 82.580 73.135 ;
        RECT 82.760 72.975 83.180 73.355 ;
        RECT 82.410 72.805 82.580 72.885 ;
        RECT 83.380 72.805 83.620 73.095 ;
        RECT 80.180 72.555 81.550 72.805 ;
        RECT 80.180 72.295 80.430 72.555 ;
        RECT 80.940 72.125 81.190 72.285 ;
        RECT 79.840 71.955 81.190 72.125 ;
        RECT 79.840 71.915 80.260 71.955 ;
        RECT 79.570 71.365 79.920 71.735 ;
        RECT 78.275 70.805 78.605 71.185 ;
        RECT 78.775 71.025 78.945 71.355 ;
        RECT 80.090 71.185 80.260 71.915 ;
        RECT 81.360 71.785 81.550 72.555 ;
        RECT 80.430 71.455 80.840 71.785 ;
        RECT 81.130 71.445 81.550 71.785 ;
        RECT 81.720 72.375 82.240 72.685 ;
        RECT 82.410 72.635 83.620 72.805 ;
        RECT 83.850 72.665 84.180 73.355 ;
        RECT 81.720 71.615 81.890 72.375 ;
        RECT 82.060 71.785 82.240 72.195 ;
        RECT 82.410 72.125 82.580 72.635 ;
        RECT 84.350 72.485 84.520 73.095 ;
        RECT 84.790 72.635 85.120 73.145 ;
        RECT 84.350 72.465 84.670 72.485 ;
        RECT 82.750 72.295 84.670 72.465 ;
        RECT 82.410 71.955 84.310 72.125 ;
        RECT 82.640 71.615 82.970 71.735 ;
        RECT 81.720 71.445 82.970 71.615 ;
        RECT 79.245 70.985 80.260 71.185 ;
        RECT 80.430 70.805 80.840 71.245 ;
        RECT 81.130 71.015 81.380 71.445 ;
        RECT 81.580 70.805 81.900 71.265 ;
        RECT 83.140 71.195 83.310 71.955 ;
        RECT 83.980 71.895 84.310 71.955 ;
        RECT 83.500 71.725 83.830 71.785 ;
        RECT 83.500 71.455 84.160 71.725 ;
        RECT 84.480 71.400 84.670 72.295 ;
        RECT 82.460 71.025 83.310 71.195 ;
        RECT 83.510 70.805 84.170 71.285 ;
        RECT 84.350 71.070 84.670 71.400 ;
        RECT 84.870 72.045 85.120 72.635 ;
        RECT 85.300 72.555 85.585 73.355 ;
        RECT 85.765 73.015 86.020 73.045 ;
        RECT 85.765 72.845 86.105 73.015 ;
        RECT 86.565 72.920 91.910 73.355 ;
        RECT 85.765 72.375 86.020 72.845 ;
        RECT 84.870 71.715 85.670 72.045 ;
        RECT 84.870 71.065 85.120 71.715 ;
        RECT 85.840 71.515 86.020 72.375 ;
        RECT 85.300 70.805 85.585 71.265 ;
        RECT 85.765 70.985 86.020 71.515 ;
        RECT 88.150 71.350 88.490 72.180 ;
        RECT 89.970 71.670 90.320 72.920 ;
        RECT 92.745 72.685 93.025 73.355 ;
        RECT 93.195 72.465 93.495 73.015 ;
        RECT 93.695 72.635 94.025 73.355 ;
        RECT 94.215 72.635 94.675 73.185 ;
        RECT 92.560 72.045 92.825 72.405 ;
        RECT 93.195 72.295 94.135 72.465 ;
        RECT 93.965 72.045 94.135 72.295 ;
        RECT 92.560 71.795 93.235 72.045 ;
        RECT 93.455 71.795 93.795 72.045 ;
        RECT 93.965 71.715 94.255 72.045 ;
        RECT 93.965 71.625 94.135 71.715 ;
        RECT 92.745 71.435 94.135 71.625 ;
        RECT 86.565 70.805 91.910 71.350 ;
        RECT 92.745 71.075 93.075 71.435 ;
        RECT 94.425 71.265 94.675 72.635 ;
        RECT 95.765 72.190 96.055 73.355 ;
        RECT 96.225 72.920 101.570 73.355 ;
        RECT 101.745 72.920 107.090 73.355 ;
        RECT 93.695 70.805 93.945 71.265 ;
        RECT 94.115 70.975 94.675 71.265 ;
        RECT 95.765 70.805 96.055 71.530 ;
        RECT 97.810 71.350 98.150 72.180 ;
        RECT 99.630 71.670 99.980 72.920 ;
        RECT 103.330 71.350 103.670 72.180 ;
        RECT 105.150 71.670 105.500 72.920 ;
        RECT 107.265 72.265 110.775 73.355 ;
        RECT 110.945 72.265 112.155 73.355 ;
        RECT 107.265 71.575 108.915 72.095 ;
        RECT 109.085 71.745 110.775 72.265 ;
        RECT 96.225 70.805 101.570 71.350 ;
        RECT 101.745 70.805 107.090 71.350 ;
        RECT 107.265 70.805 110.775 71.575 ;
        RECT 110.945 71.555 111.465 72.095 ;
        RECT 111.635 71.725 112.155 72.265 ;
        RECT 112.325 72.265 113.535 73.355 ;
        RECT 112.325 71.725 112.845 72.265 ;
        RECT 113.015 71.555 113.535 72.095 ;
        RECT 110.945 70.805 112.155 71.555 ;
        RECT 112.325 70.805 113.535 71.555 ;
        RECT 5.520 70.635 113.620 70.805 ;
        RECT 5.605 69.885 6.815 70.635 ;
        RECT 6.985 70.090 12.330 70.635 ;
        RECT 5.605 69.345 6.125 69.885 ;
        RECT 6.295 69.175 6.815 69.715 ;
        RECT 8.570 69.260 8.910 70.090 ;
        RECT 12.970 69.895 13.225 70.465 ;
        RECT 13.395 70.235 13.725 70.635 ;
        RECT 14.150 70.100 14.680 70.465 ;
        RECT 14.870 70.295 15.145 70.465 ;
        RECT 14.865 70.125 15.145 70.295 ;
        RECT 14.150 70.065 14.325 70.100 ;
        RECT 13.395 69.895 14.325 70.065 ;
        RECT 5.605 68.085 6.815 69.175 ;
        RECT 10.390 68.520 10.740 69.770 ;
        RECT 12.970 69.225 13.140 69.895 ;
        RECT 13.395 69.725 13.565 69.895 ;
        RECT 13.310 69.395 13.565 69.725 ;
        RECT 13.790 69.395 13.985 69.725 ;
        RECT 6.985 68.085 12.330 68.520 ;
        RECT 12.970 68.255 13.305 69.225 ;
        RECT 13.475 68.085 13.645 69.225 ;
        RECT 13.815 68.425 13.985 69.395 ;
        RECT 14.155 68.765 14.325 69.895 ;
        RECT 14.495 69.105 14.665 69.905 ;
        RECT 14.870 69.305 15.145 70.125 ;
        RECT 15.315 69.105 15.505 70.465 ;
        RECT 15.685 70.100 16.195 70.635 ;
        RECT 16.415 69.825 16.660 70.430 ;
        RECT 18.025 69.960 18.295 70.305 ;
        RECT 18.485 70.235 18.865 70.635 ;
        RECT 19.035 70.065 19.205 70.415 ;
        RECT 19.375 70.235 19.705 70.635 ;
        RECT 19.905 70.065 20.075 70.415 ;
        RECT 20.275 70.135 20.605 70.635 ;
        RECT 15.705 69.655 16.935 69.825 ;
        RECT 14.495 68.935 15.505 69.105 ;
        RECT 15.675 69.090 16.425 69.280 ;
        RECT 14.155 68.595 15.280 68.765 ;
        RECT 15.675 68.425 15.845 69.090 ;
        RECT 16.595 68.845 16.935 69.655 ;
        RECT 13.815 68.255 15.845 68.425 ;
        RECT 16.015 68.085 16.185 68.845 ;
        RECT 16.420 68.435 16.935 68.845 ;
        RECT 18.025 69.225 18.195 69.960 ;
        RECT 18.465 69.895 20.075 70.065 ;
        RECT 18.465 69.725 18.635 69.895 ;
        RECT 18.365 69.395 18.635 69.725 ;
        RECT 18.805 69.395 19.210 69.725 ;
        RECT 18.465 69.225 18.635 69.395 ;
        RECT 19.380 69.275 20.090 69.725 ;
        RECT 20.260 69.395 20.610 69.965 ;
        RECT 20.785 69.835 21.125 70.465 ;
        RECT 21.295 69.835 21.545 70.635 ;
        RECT 21.735 69.985 22.065 70.465 ;
        RECT 22.235 70.175 22.460 70.635 ;
        RECT 22.630 69.985 22.960 70.465 ;
        RECT 20.785 69.785 21.015 69.835 ;
        RECT 21.735 69.815 22.960 69.985 ;
        RECT 23.590 69.855 24.090 70.465 ;
        RECT 25.590 69.855 26.090 70.465 ;
        RECT 18.025 68.255 18.295 69.225 ;
        RECT 18.465 69.055 19.190 69.225 ;
        RECT 19.380 69.105 20.095 69.275 ;
        RECT 20.785 69.225 20.960 69.785 ;
        RECT 21.130 69.475 21.825 69.645 ;
        RECT 21.655 69.225 21.825 69.475 ;
        RECT 22.000 69.445 22.420 69.645 ;
        RECT 22.590 69.445 22.920 69.645 ;
        RECT 23.090 69.445 23.420 69.645 ;
        RECT 23.590 69.225 23.760 69.855 ;
        RECT 23.945 69.395 24.295 69.645 ;
        RECT 25.385 69.395 25.735 69.645 ;
        RECT 25.920 69.225 26.090 69.855 ;
        RECT 26.720 69.985 27.050 70.465 ;
        RECT 27.220 70.175 27.445 70.635 ;
        RECT 27.615 69.985 27.945 70.465 ;
        RECT 26.720 69.815 27.945 69.985 ;
        RECT 28.135 69.835 28.385 70.635 ;
        RECT 28.555 69.835 28.895 70.465 ;
        RECT 28.665 69.785 28.895 69.835 ;
        RECT 26.260 69.445 26.590 69.645 ;
        RECT 26.760 69.445 27.090 69.645 ;
        RECT 27.260 69.445 27.680 69.645 ;
        RECT 27.855 69.475 28.550 69.645 ;
        RECT 27.855 69.225 28.025 69.475 ;
        RECT 28.720 69.225 28.895 69.785 ;
        RECT 29.065 69.865 30.735 70.635 ;
        RECT 31.365 69.910 31.655 70.635 ;
        RECT 31.835 70.135 32.165 70.635 ;
        RECT 32.365 70.065 32.535 70.415 ;
        RECT 32.735 70.235 33.065 70.635 ;
        RECT 33.235 70.065 33.405 70.415 ;
        RECT 33.575 70.235 33.955 70.635 ;
        RECT 29.065 69.345 29.815 69.865 ;
        RECT 19.020 68.935 19.190 69.055 ;
        RECT 20.290 68.935 20.610 69.225 ;
        RECT 18.505 68.085 18.785 68.885 ;
        RECT 19.020 68.765 20.610 68.935 ;
        RECT 18.955 68.305 20.610 68.595 ;
        RECT 20.785 68.255 21.125 69.225 ;
        RECT 21.295 68.085 21.465 69.225 ;
        RECT 21.655 69.055 24.090 69.225 ;
        RECT 21.735 68.085 21.985 68.885 ;
        RECT 22.630 68.255 22.960 69.055 ;
        RECT 23.260 68.085 23.590 68.885 ;
        RECT 23.760 68.255 24.090 69.055 ;
        RECT 25.590 69.055 28.025 69.225 ;
        RECT 25.590 68.255 25.920 69.055 ;
        RECT 26.090 68.085 26.420 68.885 ;
        RECT 26.720 68.255 27.050 69.055 ;
        RECT 27.695 68.085 27.945 68.885 ;
        RECT 28.215 68.085 28.385 69.225 ;
        RECT 28.555 68.255 28.895 69.225 ;
        RECT 29.985 69.175 30.735 69.695 ;
        RECT 31.830 69.395 32.180 69.965 ;
        RECT 32.365 69.895 33.975 70.065 ;
        RECT 34.145 69.960 34.415 70.305 ;
        RECT 33.805 69.725 33.975 69.895 ;
        RECT 32.350 69.275 33.060 69.725 ;
        RECT 33.230 69.395 33.635 69.725 ;
        RECT 33.805 69.395 34.075 69.725 ;
        RECT 29.065 68.085 30.735 69.175 ;
        RECT 31.365 68.085 31.655 69.250 ;
        RECT 31.830 68.935 32.150 69.225 ;
        RECT 32.345 69.105 33.060 69.275 ;
        RECT 33.805 69.225 33.975 69.395 ;
        RECT 34.245 69.225 34.415 69.960 ;
        RECT 34.585 69.865 36.255 70.635 ;
        RECT 36.885 69.960 37.145 70.465 ;
        RECT 37.325 70.255 37.655 70.635 ;
        RECT 37.835 70.085 38.005 70.465 ;
        RECT 34.585 69.345 35.335 69.865 ;
        RECT 33.250 69.055 33.975 69.225 ;
        RECT 33.250 68.935 33.420 69.055 ;
        RECT 31.830 68.765 33.420 68.935 ;
        RECT 31.830 68.305 33.485 68.595 ;
        RECT 33.655 68.085 33.935 68.885 ;
        RECT 34.145 68.255 34.415 69.225 ;
        RECT 35.505 69.175 36.255 69.695 ;
        RECT 34.585 68.085 36.255 69.175 ;
        RECT 36.885 69.160 37.055 69.960 ;
        RECT 37.340 69.915 38.005 70.085 ;
        RECT 37.340 69.660 37.510 69.915 ;
        RECT 39.190 69.895 39.445 70.465 ;
        RECT 39.615 70.235 39.945 70.635 ;
        RECT 40.370 70.100 40.900 70.465 ;
        RECT 41.090 70.295 41.365 70.465 ;
        RECT 41.085 70.125 41.365 70.295 ;
        RECT 40.370 70.065 40.545 70.100 ;
        RECT 39.615 69.895 40.545 70.065 ;
        RECT 37.225 69.330 37.510 69.660 ;
        RECT 37.745 69.365 38.075 69.735 ;
        RECT 37.340 69.185 37.510 69.330 ;
        RECT 39.190 69.225 39.360 69.895 ;
        RECT 39.615 69.725 39.785 69.895 ;
        RECT 39.530 69.395 39.785 69.725 ;
        RECT 40.010 69.395 40.205 69.725 ;
        RECT 36.885 68.255 37.155 69.160 ;
        RECT 37.340 69.015 38.005 69.185 ;
        RECT 37.325 68.085 37.655 68.845 ;
        RECT 37.835 68.255 38.005 69.015 ;
        RECT 39.190 68.255 39.525 69.225 ;
        RECT 39.695 68.085 39.865 69.225 ;
        RECT 40.035 68.425 40.205 69.395 ;
        RECT 40.375 68.765 40.545 69.895 ;
        RECT 40.715 69.105 40.885 69.905 ;
        RECT 41.090 69.305 41.365 70.125 ;
        RECT 41.535 69.105 41.725 70.465 ;
        RECT 41.905 70.100 42.415 70.635 ;
        RECT 42.635 69.825 42.880 70.430 ;
        RECT 43.325 69.960 43.585 70.465 ;
        RECT 43.765 70.255 44.095 70.635 ;
        RECT 44.275 70.085 44.445 70.465 ;
        RECT 41.925 69.655 43.155 69.825 ;
        RECT 40.715 68.935 41.725 69.105 ;
        RECT 41.895 69.090 42.645 69.280 ;
        RECT 40.375 68.595 41.500 68.765 ;
        RECT 41.895 68.425 42.065 69.090 ;
        RECT 42.815 68.845 43.155 69.655 ;
        RECT 40.035 68.255 42.065 68.425 ;
        RECT 42.235 68.085 42.405 68.845 ;
        RECT 42.640 68.435 43.155 68.845 ;
        RECT 43.325 69.160 43.495 69.960 ;
        RECT 43.780 69.915 44.445 70.085 ;
        RECT 43.780 69.660 43.950 69.915 ;
        RECT 44.745 69.815 44.975 70.635 ;
        RECT 45.145 69.835 45.475 70.465 ;
        RECT 43.665 69.330 43.950 69.660 ;
        RECT 44.185 69.365 44.515 69.735 ;
        RECT 44.725 69.395 45.055 69.645 ;
        RECT 43.780 69.185 43.950 69.330 ;
        RECT 45.225 69.235 45.475 69.835 ;
        RECT 45.645 69.815 45.855 70.635 ;
        RECT 46.085 69.865 49.595 70.635 ;
        RECT 50.235 70.135 50.565 70.635 ;
        RECT 50.765 70.065 50.935 70.415 ;
        RECT 51.135 70.235 51.465 70.635 ;
        RECT 51.635 70.065 51.805 70.415 ;
        RECT 51.975 70.235 52.355 70.635 ;
        RECT 46.085 69.345 47.735 69.865 ;
        RECT 43.325 68.255 43.595 69.160 ;
        RECT 43.780 69.015 44.445 69.185 ;
        RECT 43.765 68.085 44.095 68.845 ;
        RECT 44.275 68.255 44.445 69.015 ;
        RECT 44.745 68.085 44.975 69.225 ;
        RECT 45.145 68.255 45.475 69.235 ;
        RECT 45.645 68.085 45.855 69.225 ;
        RECT 47.905 69.175 49.595 69.695 ;
        RECT 50.230 69.395 50.580 69.965 ;
        RECT 50.765 69.895 52.375 70.065 ;
        RECT 52.545 69.960 52.815 70.305 ;
        RECT 53.045 70.155 53.325 70.635 ;
        RECT 53.495 69.985 53.755 70.375 ;
        RECT 53.930 70.155 54.185 70.635 ;
        RECT 54.355 69.985 54.650 70.375 ;
        RECT 54.830 70.155 55.105 70.635 ;
        RECT 55.275 70.135 55.575 70.465 ;
        RECT 52.205 69.725 52.375 69.895 ;
        RECT 46.085 68.085 49.595 69.175 ;
        RECT 50.230 68.935 50.550 69.225 ;
        RECT 50.750 69.105 51.460 69.725 ;
        RECT 51.630 69.395 52.035 69.725 ;
        RECT 52.205 69.395 52.475 69.725 ;
        RECT 52.205 69.225 52.375 69.395 ;
        RECT 52.645 69.225 52.815 69.960 ;
        RECT 51.650 69.055 52.375 69.225 ;
        RECT 51.650 68.935 51.820 69.055 ;
        RECT 50.230 68.765 51.820 68.935 ;
        RECT 50.230 68.305 51.885 68.595 ;
        RECT 52.055 68.085 52.335 68.885 ;
        RECT 52.545 68.255 52.815 69.225 ;
        RECT 53.000 69.815 54.650 69.985 ;
        RECT 53.000 69.305 53.405 69.815 ;
        RECT 53.575 69.475 54.715 69.645 ;
        RECT 53.000 69.135 53.755 69.305 ;
        RECT 53.040 68.085 53.325 68.955 ;
        RECT 53.495 68.885 53.755 69.135 ;
        RECT 54.545 69.225 54.715 69.475 ;
        RECT 54.885 69.395 55.235 69.965 ;
        RECT 55.405 69.225 55.575 70.135 ;
        RECT 55.745 69.885 56.955 70.635 ;
        RECT 57.125 69.910 57.415 70.635 ;
        RECT 57.585 69.885 58.795 70.635 ;
        RECT 55.745 69.345 56.265 69.885 ;
        RECT 54.545 69.055 55.575 69.225 ;
        RECT 56.435 69.175 56.955 69.715 ;
        RECT 57.585 69.345 58.105 69.885 ;
        RECT 58.970 69.795 59.230 70.635 ;
        RECT 59.405 69.890 59.660 70.465 ;
        RECT 59.830 70.255 60.160 70.635 ;
        RECT 60.375 70.085 60.545 70.465 ;
        RECT 59.830 69.915 60.545 70.085 ;
        RECT 61.265 70.135 61.525 70.465 ;
        RECT 61.695 70.275 62.025 70.635 ;
        RECT 62.280 70.255 63.580 70.465 ;
        RECT 61.265 70.125 61.495 70.135 ;
        RECT 53.495 68.715 54.615 68.885 ;
        RECT 53.495 68.255 53.755 68.715 ;
        RECT 53.930 68.085 54.185 68.545 ;
        RECT 54.355 68.255 54.615 68.715 ;
        RECT 54.785 68.085 55.095 68.885 ;
        RECT 55.265 68.255 55.575 69.055 ;
        RECT 55.745 68.085 56.955 69.175 ;
        RECT 57.125 68.085 57.415 69.250 ;
        RECT 58.275 69.175 58.795 69.715 ;
        RECT 57.585 68.085 58.795 69.175 ;
        RECT 58.970 68.085 59.230 69.235 ;
        RECT 59.405 69.160 59.575 69.890 ;
        RECT 59.830 69.725 60.000 69.915 ;
        RECT 59.745 69.395 60.000 69.725 ;
        RECT 59.830 69.185 60.000 69.395 ;
        RECT 60.280 69.365 60.635 69.735 ;
        RECT 59.405 68.255 59.660 69.160 ;
        RECT 59.830 69.015 60.545 69.185 ;
        RECT 59.830 68.085 60.160 68.845 ;
        RECT 60.375 68.255 60.545 69.015 ;
        RECT 61.265 68.935 61.435 70.125 ;
        RECT 62.280 70.105 62.450 70.255 ;
        RECT 61.695 69.980 62.450 70.105 ;
        RECT 61.605 69.935 62.450 69.980 ;
        RECT 61.605 69.815 61.875 69.935 ;
        RECT 61.605 69.240 61.775 69.815 ;
        RECT 62.005 69.375 62.415 69.680 ;
        RECT 62.705 69.645 62.915 70.045 ;
        RECT 62.585 69.435 62.915 69.645 ;
        RECT 63.160 69.645 63.380 70.045 ;
        RECT 63.855 69.870 64.310 70.635 ;
        RECT 64.485 69.865 67.075 70.635 ;
        RECT 67.710 70.085 67.965 70.375 ;
        RECT 68.135 70.255 68.465 70.635 ;
        RECT 67.710 69.915 68.460 70.085 ;
        RECT 63.160 69.435 63.635 69.645 ;
        RECT 63.825 69.445 64.315 69.645 ;
        RECT 64.485 69.345 65.695 69.865 ;
        RECT 61.605 69.205 61.805 69.240 ;
        RECT 63.135 69.205 64.310 69.265 ;
        RECT 61.605 69.095 64.310 69.205 ;
        RECT 65.865 69.175 67.075 69.695 ;
        RECT 61.665 69.035 63.465 69.095 ;
        RECT 63.135 69.005 63.465 69.035 ;
        RECT 61.265 68.255 61.525 68.935 ;
        RECT 61.695 68.085 61.945 68.865 ;
        RECT 62.195 68.835 63.030 68.845 ;
        RECT 63.620 68.835 63.805 68.925 ;
        RECT 62.195 68.635 63.805 68.835 ;
        RECT 62.195 68.255 62.445 68.635 ;
        RECT 63.575 68.595 63.805 68.635 ;
        RECT 64.055 68.475 64.310 69.095 ;
        RECT 62.615 68.085 62.970 68.465 ;
        RECT 63.975 68.255 64.310 68.475 ;
        RECT 64.485 68.085 67.075 69.175 ;
        RECT 67.710 69.095 68.060 69.745 ;
        RECT 68.230 68.925 68.460 69.915 ;
        RECT 67.710 68.755 68.460 68.925 ;
        RECT 67.710 68.255 67.965 68.755 ;
        RECT 68.135 68.085 68.465 68.585 ;
        RECT 68.635 68.255 68.805 70.375 ;
        RECT 69.165 70.275 69.495 70.635 ;
        RECT 69.665 70.245 70.160 70.415 ;
        RECT 70.365 70.245 71.220 70.415 ;
        RECT 69.035 69.055 69.495 70.105 ;
        RECT 68.975 68.270 69.300 69.055 ;
        RECT 69.665 68.885 69.835 70.245 ;
        RECT 70.005 69.335 70.355 69.955 ;
        RECT 70.525 69.735 70.880 69.955 ;
        RECT 70.525 69.145 70.695 69.735 ;
        RECT 71.050 69.535 71.220 70.245 ;
        RECT 72.095 70.175 72.425 70.635 ;
        RECT 72.635 70.275 72.985 70.445 ;
        RECT 71.425 69.705 72.215 69.955 ;
        RECT 72.635 69.885 72.895 70.275 ;
        RECT 73.205 70.185 74.155 70.465 ;
        RECT 74.325 70.195 74.515 70.635 ;
        RECT 74.685 70.255 75.755 70.425 ;
        RECT 72.385 69.535 72.555 69.715 ;
        RECT 69.665 68.715 70.060 68.885 ;
        RECT 70.230 68.755 70.695 69.145 ;
        RECT 70.865 69.365 72.555 69.535 ;
        RECT 69.890 68.585 70.060 68.715 ;
        RECT 70.865 68.585 71.035 69.365 ;
        RECT 72.725 69.195 72.895 69.885 ;
        RECT 71.395 69.025 72.895 69.195 ;
        RECT 73.085 69.225 73.295 70.015 ;
        RECT 73.465 69.395 73.815 70.015 ;
        RECT 73.985 69.405 74.155 70.185 ;
        RECT 74.685 70.025 74.855 70.255 ;
        RECT 74.325 69.855 74.855 70.025 ;
        RECT 74.325 69.575 74.545 69.855 ;
        RECT 75.025 69.685 75.265 70.085 ;
        RECT 73.985 69.235 74.390 69.405 ;
        RECT 74.725 69.315 75.265 69.685 ;
        RECT 75.435 69.900 75.755 70.255 ;
        RECT 76.000 70.175 76.305 70.635 ;
        RECT 76.475 69.925 76.730 70.455 ;
        RECT 75.435 69.725 75.760 69.900 ;
        RECT 75.435 69.425 76.350 69.725 ;
        RECT 75.610 69.395 76.350 69.425 ;
        RECT 73.085 69.065 73.760 69.225 ;
        RECT 74.220 69.145 74.390 69.235 ;
        RECT 73.085 69.055 74.050 69.065 ;
        RECT 72.725 68.885 72.895 69.025 ;
        RECT 69.470 68.085 69.720 68.545 ;
        RECT 69.890 68.255 70.140 68.585 ;
        RECT 70.355 68.255 71.035 68.585 ;
        RECT 71.205 68.685 72.280 68.855 ;
        RECT 72.725 68.715 73.285 68.885 ;
        RECT 73.590 68.765 74.050 69.055 ;
        RECT 74.220 68.975 75.440 69.145 ;
        RECT 71.205 68.345 71.375 68.685 ;
        RECT 71.610 68.085 71.940 68.515 ;
        RECT 72.110 68.345 72.280 68.685 ;
        RECT 72.575 68.085 72.945 68.545 ;
        RECT 73.115 68.255 73.285 68.715 ;
        RECT 74.220 68.595 74.390 68.975 ;
        RECT 75.610 68.805 75.780 69.395 ;
        RECT 76.520 69.275 76.730 69.925 ;
        RECT 73.520 68.255 74.390 68.595 ;
        RECT 74.980 68.635 75.780 68.805 ;
        RECT 74.560 68.085 74.810 68.545 ;
        RECT 74.980 68.345 75.150 68.635 ;
        RECT 75.330 68.085 75.660 68.465 ;
        RECT 76.000 68.085 76.305 69.225 ;
        RECT 76.475 68.395 76.730 69.275 ;
        RECT 76.905 69.960 77.175 70.305 ;
        RECT 77.365 70.235 77.745 70.635 ;
        RECT 77.915 70.065 78.085 70.415 ;
        RECT 78.255 70.235 78.585 70.635 ;
        RECT 78.785 70.065 78.955 70.415 ;
        RECT 79.155 70.135 79.485 70.635 ;
        RECT 76.905 69.225 77.075 69.960 ;
        RECT 77.345 69.895 78.955 70.065 ;
        RECT 77.345 69.725 77.515 69.895 ;
        RECT 77.245 69.395 77.515 69.725 ;
        RECT 77.685 69.395 78.090 69.725 ;
        RECT 77.345 69.225 77.515 69.395 ;
        RECT 78.260 69.275 78.970 69.725 ;
        RECT 79.140 69.395 79.490 69.965 ;
        RECT 79.665 69.865 82.255 70.635 ;
        RECT 82.885 69.910 83.175 70.635 ;
        RECT 83.345 70.090 88.690 70.635 ;
        RECT 79.665 69.345 80.875 69.865 ;
        RECT 76.905 68.255 77.175 69.225 ;
        RECT 77.345 69.055 78.070 69.225 ;
        RECT 78.260 69.105 78.975 69.275 ;
        RECT 77.900 68.935 78.070 69.055 ;
        RECT 79.170 68.935 79.490 69.225 ;
        RECT 81.045 69.175 82.255 69.695 ;
        RECT 84.930 69.260 85.270 70.090 ;
        RECT 88.865 69.885 90.075 70.635 ;
        RECT 77.385 68.085 77.665 68.885 ;
        RECT 77.900 68.765 79.490 68.935 ;
        RECT 77.835 68.305 79.490 68.595 ;
        RECT 79.665 68.085 82.255 69.175 ;
        RECT 82.885 68.085 83.175 69.250 ;
        RECT 86.750 68.520 87.100 69.770 ;
        RECT 88.865 69.345 89.385 69.885 ;
        RECT 90.450 69.855 90.950 70.465 ;
        RECT 89.555 69.175 90.075 69.715 ;
        RECT 90.245 69.395 90.595 69.645 ;
        RECT 90.780 69.225 90.950 69.855 ;
        RECT 91.580 69.985 91.910 70.465 ;
        RECT 92.080 70.175 92.305 70.635 ;
        RECT 92.475 69.985 92.805 70.465 ;
        RECT 91.580 69.815 92.805 69.985 ;
        RECT 92.995 69.835 93.245 70.635 ;
        RECT 93.415 69.835 93.755 70.465 ;
        RECT 93.925 70.090 99.270 70.635 ;
        RECT 91.120 69.445 91.450 69.645 ;
        RECT 91.620 69.445 91.950 69.645 ;
        RECT 92.120 69.445 92.540 69.645 ;
        RECT 92.715 69.475 93.410 69.645 ;
        RECT 92.715 69.225 92.885 69.475 ;
        RECT 93.580 69.225 93.755 69.835 ;
        RECT 95.510 69.260 95.850 70.090 ;
        RECT 99.995 70.085 100.165 70.465 ;
        RECT 100.345 70.255 100.675 70.635 ;
        RECT 99.995 69.915 100.660 70.085 ;
        RECT 100.855 69.960 101.115 70.465 ;
        RECT 83.345 68.085 88.690 68.520 ;
        RECT 88.865 68.085 90.075 69.175 ;
        RECT 90.450 69.055 92.885 69.225 ;
        RECT 90.450 68.255 90.780 69.055 ;
        RECT 90.950 68.085 91.280 68.885 ;
        RECT 91.580 68.255 91.910 69.055 ;
        RECT 92.555 68.085 92.805 68.885 ;
        RECT 93.075 68.085 93.245 69.225 ;
        RECT 93.415 68.255 93.755 69.225 ;
        RECT 97.330 68.520 97.680 69.770 ;
        RECT 99.925 69.365 100.255 69.735 ;
        RECT 100.490 69.660 100.660 69.915 ;
        RECT 100.490 69.330 100.775 69.660 ;
        RECT 100.490 69.185 100.660 69.330 ;
        RECT 99.995 69.015 100.660 69.185 ;
        RECT 100.945 69.160 101.115 69.960 ;
        RECT 101.285 69.865 102.955 70.635 ;
        RECT 103.215 70.085 103.385 70.465 ;
        RECT 103.565 70.255 103.895 70.635 ;
        RECT 103.215 69.915 103.880 70.085 ;
        RECT 104.075 69.960 104.335 70.465 ;
        RECT 101.285 69.345 102.035 69.865 ;
        RECT 102.205 69.175 102.955 69.695 ;
        RECT 103.145 69.365 103.475 69.735 ;
        RECT 103.710 69.660 103.880 69.915 ;
        RECT 103.710 69.330 103.995 69.660 ;
        RECT 103.710 69.185 103.880 69.330 ;
        RECT 93.925 68.085 99.270 68.520 ;
        RECT 99.995 68.255 100.165 69.015 ;
        RECT 100.345 68.085 100.675 68.845 ;
        RECT 100.845 68.255 101.115 69.160 ;
        RECT 101.285 68.085 102.955 69.175 ;
        RECT 103.215 69.015 103.880 69.185 ;
        RECT 104.165 69.160 104.335 69.960 ;
        RECT 105.025 69.815 105.235 70.635 ;
        RECT 105.405 69.835 105.735 70.465 ;
        RECT 105.405 69.235 105.655 69.835 ;
        RECT 105.905 69.815 106.135 70.635 ;
        RECT 106.345 69.865 108.015 70.635 ;
        RECT 108.645 69.910 108.935 70.635 ;
        RECT 109.105 69.865 111.695 70.635 ;
        RECT 112.325 69.885 113.535 70.635 ;
        RECT 105.825 69.395 106.155 69.645 ;
        RECT 106.345 69.345 107.095 69.865 ;
        RECT 103.215 68.255 103.385 69.015 ;
        RECT 103.565 68.085 103.895 68.845 ;
        RECT 104.065 68.255 104.335 69.160 ;
        RECT 105.025 68.085 105.235 69.225 ;
        RECT 105.405 68.255 105.735 69.235 ;
        RECT 105.905 68.085 106.135 69.225 ;
        RECT 107.265 69.175 108.015 69.695 ;
        RECT 109.105 69.345 110.315 69.865 ;
        RECT 106.345 68.085 108.015 69.175 ;
        RECT 108.645 68.085 108.935 69.250 ;
        RECT 110.485 69.175 111.695 69.695 ;
        RECT 109.105 68.085 111.695 69.175 ;
        RECT 112.325 69.175 112.845 69.715 ;
        RECT 113.015 69.345 113.535 69.885 ;
        RECT 112.325 68.085 113.535 69.175 ;
        RECT 5.520 67.915 113.620 68.085 ;
        RECT 5.605 66.825 6.815 67.915 ;
        RECT 6.985 66.825 9.575 67.915 ;
        RECT 5.605 66.115 6.125 66.655 ;
        RECT 6.295 66.285 6.815 66.825 ;
        RECT 6.985 66.135 8.195 66.655 ;
        RECT 8.365 66.305 9.575 66.825 ;
        RECT 9.745 66.840 10.015 67.745 ;
        RECT 10.185 67.155 10.515 67.915 ;
        RECT 10.695 66.985 10.865 67.745 ;
        RECT 5.605 65.365 6.815 66.115 ;
        RECT 6.985 65.365 9.575 66.135 ;
        RECT 9.745 66.040 9.915 66.840 ;
        RECT 10.200 66.815 10.865 66.985 ;
        RECT 11.125 66.840 11.395 67.745 ;
        RECT 11.565 67.155 11.895 67.915 ;
        RECT 12.075 66.985 12.245 67.745 ;
        RECT 10.200 66.670 10.370 66.815 ;
        RECT 10.085 66.340 10.370 66.670 ;
        RECT 10.200 66.085 10.370 66.340 ;
        RECT 10.605 66.265 10.935 66.635 ;
        RECT 9.745 65.535 10.005 66.040 ;
        RECT 10.200 65.915 10.865 66.085 ;
        RECT 10.185 65.365 10.515 65.745 ;
        RECT 10.695 65.535 10.865 65.915 ;
        RECT 11.125 66.040 11.295 66.840 ;
        RECT 11.580 66.815 12.245 66.985 ;
        RECT 11.580 66.670 11.750 66.815 ;
        RECT 12.565 66.775 12.775 67.915 ;
        RECT 11.465 66.340 11.750 66.670 ;
        RECT 12.945 66.765 13.275 67.745 ;
        RECT 13.445 66.775 13.675 67.915 ;
        RECT 14.350 66.775 14.685 67.745 ;
        RECT 14.855 66.775 15.025 67.915 ;
        RECT 15.195 67.575 17.225 67.745 ;
        RECT 11.580 66.085 11.750 66.340 ;
        RECT 11.985 66.265 12.315 66.635 ;
        RECT 11.125 65.535 11.385 66.040 ;
        RECT 11.580 65.915 12.245 66.085 ;
        RECT 11.565 65.365 11.895 65.745 ;
        RECT 12.075 65.535 12.245 65.915 ;
        RECT 12.565 65.365 12.775 66.185 ;
        RECT 12.945 66.165 13.195 66.765 ;
        RECT 13.365 66.355 13.695 66.605 ;
        RECT 12.945 65.535 13.275 66.165 ;
        RECT 13.445 65.365 13.675 66.185 ;
        RECT 14.350 66.105 14.520 66.775 ;
        RECT 15.195 66.605 15.365 67.575 ;
        RECT 14.690 66.275 14.945 66.605 ;
        RECT 15.170 66.275 15.365 66.605 ;
        RECT 15.535 67.235 16.660 67.405 ;
        RECT 14.775 66.105 14.945 66.275 ;
        RECT 15.535 66.105 15.705 67.235 ;
        RECT 14.350 65.535 14.605 66.105 ;
        RECT 14.775 65.935 15.705 66.105 ;
        RECT 15.875 66.895 16.885 67.065 ;
        RECT 15.875 66.095 16.045 66.895 ;
        RECT 15.530 65.900 15.705 65.935 ;
        RECT 14.775 65.365 15.105 65.765 ;
        RECT 15.530 65.535 16.060 65.900 ;
        RECT 16.250 65.875 16.525 66.695 ;
        RECT 16.245 65.705 16.525 65.875 ;
        RECT 16.250 65.535 16.525 65.705 ;
        RECT 16.695 65.535 16.885 66.895 ;
        RECT 17.055 66.910 17.225 67.575 ;
        RECT 17.395 67.155 17.565 67.915 ;
        RECT 17.800 67.155 18.315 67.565 ;
        RECT 17.055 66.720 17.805 66.910 ;
        RECT 17.975 66.345 18.315 67.155 ;
        RECT 18.485 66.750 18.775 67.915 ;
        RECT 18.945 66.825 21.535 67.915 ;
        RECT 17.085 66.175 18.315 66.345 ;
        RECT 17.065 65.365 17.575 65.900 ;
        RECT 17.795 65.570 18.040 66.175 ;
        RECT 18.945 66.135 20.155 66.655 ;
        RECT 20.325 66.305 21.535 66.825 ;
        RECT 21.910 66.945 22.240 67.745 ;
        RECT 22.410 67.115 22.740 67.915 ;
        RECT 23.040 66.945 23.370 67.745 ;
        RECT 24.015 67.115 24.265 67.915 ;
        RECT 21.910 66.775 24.345 66.945 ;
        RECT 24.535 66.775 24.705 67.915 ;
        RECT 24.875 66.775 25.215 67.745 ;
        RECT 25.385 66.825 27.055 67.915 ;
        RECT 21.705 66.355 22.055 66.605 ;
        RECT 22.240 66.145 22.410 66.775 ;
        RECT 22.580 66.355 22.910 66.555 ;
        RECT 23.080 66.355 23.410 66.555 ;
        RECT 23.580 66.355 24.000 66.555 ;
        RECT 24.175 66.525 24.345 66.775 ;
        RECT 24.175 66.355 24.870 66.525 ;
        RECT 18.485 65.365 18.775 66.090 ;
        RECT 18.945 65.365 21.535 66.135 ;
        RECT 21.910 65.535 22.410 66.145 ;
        RECT 23.040 66.015 24.265 66.185 ;
        RECT 25.040 66.165 25.215 66.775 ;
        RECT 23.040 65.535 23.370 66.015 ;
        RECT 23.540 65.365 23.765 65.825 ;
        RECT 23.935 65.535 24.265 66.015 ;
        RECT 24.455 65.365 24.705 66.165 ;
        RECT 24.875 65.535 25.215 66.165 ;
        RECT 25.385 66.135 26.135 66.655 ;
        RECT 26.305 66.305 27.055 66.825 ;
        RECT 27.890 66.945 28.220 67.745 ;
        RECT 28.390 67.115 28.720 67.915 ;
        RECT 29.020 66.945 29.350 67.745 ;
        RECT 29.995 67.115 30.245 67.915 ;
        RECT 27.890 66.775 30.325 66.945 ;
        RECT 30.515 66.775 30.685 67.915 ;
        RECT 30.855 66.775 31.195 67.745 ;
        RECT 31.365 66.825 33.955 67.915 ;
        RECT 34.130 67.245 34.385 67.745 ;
        RECT 34.555 67.415 34.885 67.915 ;
        RECT 34.130 67.075 34.880 67.245 ;
        RECT 27.685 66.355 28.035 66.605 ;
        RECT 28.220 66.145 28.390 66.775 ;
        RECT 28.560 66.355 28.890 66.555 ;
        RECT 29.060 66.355 29.390 66.555 ;
        RECT 29.560 66.355 29.980 66.555 ;
        RECT 30.155 66.525 30.325 66.775 ;
        RECT 30.155 66.355 30.850 66.525 ;
        RECT 25.385 65.365 27.055 66.135 ;
        RECT 27.890 65.535 28.390 66.145 ;
        RECT 29.020 66.015 30.245 66.185 ;
        RECT 31.020 66.165 31.195 66.775 ;
        RECT 29.020 65.535 29.350 66.015 ;
        RECT 29.520 65.365 29.745 65.825 ;
        RECT 29.915 65.535 30.245 66.015 ;
        RECT 30.435 65.365 30.685 66.165 ;
        RECT 30.855 65.535 31.195 66.165 ;
        RECT 31.365 66.135 32.575 66.655 ;
        RECT 32.745 66.305 33.955 66.825 ;
        RECT 34.130 66.255 34.480 66.905 ;
        RECT 31.365 65.365 33.955 66.135 ;
        RECT 34.650 66.085 34.880 67.075 ;
        RECT 34.130 65.915 34.880 66.085 ;
        RECT 34.130 65.625 34.385 65.915 ;
        RECT 34.555 65.365 34.885 65.745 ;
        RECT 35.055 65.625 35.225 67.745 ;
        RECT 35.395 66.945 35.720 67.730 ;
        RECT 35.890 67.455 36.140 67.915 ;
        RECT 36.310 67.415 36.560 67.745 ;
        RECT 36.775 67.415 37.455 67.745 ;
        RECT 36.310 67.285 36.480 67.415 ;
        RECT 36.085 67.115 36.480 67.285 ;
        RECT 35.455 65.895 35.915 66.945 ;
        RECT 36.085 65.755 36.255 67.115 ;
        RECT 36.650 66.855 37.115 67.245 ;
        RECT 36.425 66.045 36.775 66.665 ;
        RECT 36.945 66.265 37.115 66.855 ;
        RECT 37.285 66.635 37.455 67.415 ;
        RECT 37.625 67.315 37.795 67.655 ;
        RECT 38.030 67.485 38.360 67.915 ;
        RECT 38.530 67.315 38.700 67.655 ;
        RECT 38.995 67.455 39.365 67.915 ;
        RECT 37.625 67.145 38.700 67.315 ;
        RECT 39.535 67.285 39.705 67.745 ;
        RECT 39.940 67.405 40.810 67.745 ;
        RECT 40.980 67.455 41.230 67.915 ;
        RECT 39.145 67.115 39.705 67.285 ;
        RECT 39.145 66.975 39.315 67.115 ;
        RECT 37.815 66.805 39.315 66.975 ;
        RECT 40.010 66.945 40.470 67.235 ;
        RECT 37.285 66.465 38.975 66.635 ;
        RECT 36.945 66.045 37.300 66.265 ;
        RECT 37.470 65.755 37.640 66.465 ;
        RECT 37.845 66.045 38.635 66.295 ;
        RECT 38.805 66.285 38.975 66.465 ;
        RECT 39.145 66.115 39.315 66.805 ;
        RECT 35.585 65.365 35.915 65.725 ;
        RECT 36.085 65.585 36.580 65.755 ;
        RECT 36.785 65.585 37.640 65.755 ;
        RECT 38.515 65.365 38.845 65.825 ;
        RECT 39.055 65.725 39.315 66.115 ;
        RECT 39.505 66.935 40.470 66.945 ;
        RECT 40.640 67.025 40.810 67.405 ;
        RECT 41.400 67.365 41.570 67.655 ;
        RECT 41.750 67.535 42.080 67.915 ;
        RECT 41.400 67.195 42.200 67.365 ;
        RECT 39.505 66.775 40.180 66.935 ;
        RECT 40.640 66.855 41.860 67.025 ;
        RECT 39.505 65.985 39.715 66.775 ;
        RECT 40.640 66.765 40.810 66.855 ;
        RECT 39.885 65.985 40.235 66.605 ;
        RECT 40.405 66.595 40.810 66.765 ;
        RECT 40.405 65.815 40.575 66.595 ;
        RECT 40.745 66.145 40.965 66.425 ;
        RECT 41.145 66.315 41.685 66.685 ;
        RECT 42.030 66.605 42.200 67.195 ;
        RECT 42.420 66.775 42.725 67.915 ;
        RECT 42.895 66.725 43.150 67.605 ;
        RECT 44.245 66.750 44.535 67.915 ;
        RECT 44.705 67.480 50.050 67.915 ;
        RECT 42.030 66.575 42.770 66.605 ;
        RECT 40.745 65.975 41.275 66.145 ;
        RECT 39.055 65.555 39.405 65.725 ;
        RECT 39.625 65.535 40.575 65.815 ;
        RECT 40.745 65.365 40.935 65.805 ;
        RECT 41.105 65.745 41.275 65.975 ;
        RECT 41.445 65.915 41.685 66.315 ;
        RECT 41.855 66.275 42.770 66.575 ;
        RECT 41.855 66.100 42.180 66.275 ;
        RECT 41.855 65.745 42.175 66.100 ;
        RECT 42.940 66.075 43.150 66.725 ;
        RECT 41.105 65.575 42.175 65.745 ;
        RECT 42.420 65.365 42.725 65.825 ;
        RECT 42.895 65.545 43.150 66.075 ;
        RECT 44.245 65.365 44.535 66.090 ;
        RECT 46.290 65.910 46.630 66.740 ;
        RECT 48.110 66.230 48.460 67.480 ;
        RECT 50.890 66.945 51.220 67.745 ;
        RECT 51.390 67.115 51.720 67.915 ;
        RECT 52.020 66.945 52.350 67.745 ;
        RECT 52.995 67.115 53.245 67.915 ;
        RECT 50.890 66.775 53.325 66.945 ;
        RECT 53.515 66.775 53.685 67.915 ;
        RECT 53.855 66.775 54.195 67.745 ;
        RECT 50.685 66.355 51.035 66.605 ;
        RECT 51.220 66.145 51.390 66.775 ;
        RECT 51.560 66.355 51.890 66.555 ;
        RECT 52.060 66.355 52.390 66.555 ;
        RECT 52.560 66.355 52.980 66.555 ;
        RECT 53.155 66.525 53.325 66.775 ;
        RECT 53.155 66.355 53.850 66.525 ;
        RECT 44.705 65.365 50.050 65.910 ;
        RECT 50.890 65.535 51.390 66.145 ;
        RECT 52.020 66.015 53.245 66.185 ;
        RECT 54.020 66.165 54.195 66.775 ;
        RECT 52.020 65.535 52.350 66.015 ;
        RECT 52.520 65.365 52.745 65.825 ;
        RECT 52.915 65.535 53.245 66.015 ;
        RECT 53.435 65.365 53.685 66.165 ;
        RECT 53.855 65.535 54.195 66.165 ;
        RECT 54.825 67.325 55.525 67.745 ;
        RECT 55.725 67.555 56.055 67.915 ;
        RECT 56.225 67.325 56.555 67.725 ;
        RECT 54.825 67.095 56.555 67.325 ;
        RECT 54.825 66.125 55.030 67.095 ;
        RECT 55.200 66.355 55.530 66.895 ;
        RECT 55.705 66.605 56.030 66.895 ;
        RECT 56.225 66.875 56.555 67.095 ;
        RECT 56.725 66.605 56.895 67.530 ;
        RECT 57.075 66.855 57.405 67.915 ;
        RECT 57.590 66.765 57.850 67.915 ;
        RECT 58.025 66.840 58.280 67.745 ;
        RECT 58.450 67.155 58.780 67.915 ;
        RECT 58.995 66.985 59.165 67.745 ;
        RECT 59.435 67.105 59.730 67.915 ;
        RECT 55.705 66.275 56.200 66.605 ;
        RECT 56.520 66.275 56.895 66.605 ;
        RECT 57.105 66.275 57.415 66.605 ;
        RECT 54.825 65.535 55.535 66.125 ;
        RECT 56.045 65.895 57.405 66.105 ;
        RECT 56.045 65.535 56.375 65.895 ;
        RECT 56.575 65.365 56.905 65.725 ;
        RECT 57.075 65.535 57.405 65.895 ;
        RECT 57.590 65.365 57.850 66.205 ;
        RECT 58.025 66.110 58.195 66.840 ;
        RECT 58.450 66.815 59.165 66.985 ;
        RECT 58.450 66.605 58.620 66.815 ;
        RECT 58.365 66.275 58.620 66.605 ;
        RECT 58.025 65.535 58.280 66.110 ;
        RECT 58.450 66.085 58.620 66.275 ;
        RECT 58.900 66.265 59.255 66.635 ;
        RECT 59.910 66.605 60.155 67.745 ;
        RECT 60.330 67.105 60.590 67.915 ;
        RECT 61.190 67.910 67.465 67.915 ;
        RECT 60.770 66.605 61.020 67.740 ;
        RECT 61.190 67.115 61.450 67.910 ;
        RECT 61.620 67.015 61.880 67.740 ;
        RECT 62.050 67.185 62.310 67.910 ;
        RECT 62.480 67.015 62.740 67.740 ;
        RECT 62.910 67.185 63.170 67.910 ;
        RECT 63.340 67.015 63.600 67.740 ;
        RECT 63.770 67.185 64.030 67.910 ;
        RECT 64.200 67.015 64.460 67.740 ;
        RECT 64.630 67.185 64.875 67.910 ;
        RECT 65.045 67.015 65.305 67.740 ;
        RECT 65.490 67.185 65.735 67.910 ;
        RECT 65.905 67.015 66.165 67.740 ;
        RECT 66.350 67.185 66.595 67.910 ;
        RECT 66.765 67.015 67.025 67.740 ;
        RECT 67.210 67.185 67.465 67.910 ;
        RECT 61.620 67.000 67.025 67.015 ;
        RECT 67.635 67.000 67.925 67.740 ;
        RECT 68.095 67.170 68.365 67.915 ;
        RECT 61.620 66.895 68.365 67.000 ;
        RECT 61.620 66.775 68.395 66.895 ;
        RECT 68.625 66.825 69.835 67.915 ;
        RECT 67.200 66.725 68.395 66.775 ;
        RECT 58.450 65.915 59.165 66.085 ;
        RECT 59.425 66.045 59.740 66.605 ;
        RECT 59.910 66.355 67.030 66.605 ;
        RECT 58.450 65.365 58.780 65.745 ;
        RECT 58.995 65.535 59.165 65.915 ;
        RECT 59.425 65.365 59.730 65.875 ;
        RECT 59.910 65.545 60.160 66.355 ;
        RECT 60.330 65.365 60.590 65.890 ;
        RECT 60.770 65.545 61.020 66.355 ;
        RECT 67.200 66.185 68.365 66.725 ;
        RECT 61.620 66.015 68.365 66.185 ;
        RECT 68.625 66.115 69.145 66.655 ;
        RECT 69.315 66.285 69.835 66.825 ;
        RECT 70.005 66.750 70.295 67.915 ;
        RECT 70.465 66.825 72.135 67.915 ;
        RECT 70.465 66.135 71.215 66.655 ;
        RECT 71.385 66.305 72.135 66.825 ;
        RECT 72.805 66.775 73.035 67.915 ;
        RECT 73.205 66.765 73.535 67.745 ;
        RECT 73.705 66.775 73.915 67.915 ;
        RECT 74.145 67.480 79.490 67.915 ;
        RECT 72.785 66.355 73.115 66.605 ;
        RECT 61.190 65.365 61.450 65.925 ;
        RECT 61.620 65.560 61.880 66.015 ;
        RECT 62.050 65.365 62.310 65.845 ;
        RECT 62.480 65.560 62.740 66.015 ;
        RECT 62.910 65.365 63.170 65.845 ;
        RECT 63.340 65.560 63.600 66.015 ;
        RECT 63.770 65.365 64.015 65.845 ;
        RECT 64.185 65.560 64.460 66.015 ;
        RECT 64.630 65.365 64.875 65.845 ;
        RECT 65.045 65.560 65.305 66.015 ;
        RECT 65.485 65.365 65.735 65.845 ;
        RECT 65.905 65.560 66.165 66.015 ;
        RECT 66.345 65.365 66.595 65.845 ;
        RECT 66.765 65.560 67.025 66.015 ;
        RECT 67.205 65.365 67.465 65.845 ;
        RECT 67.635 65.560 67.895 66.015 ;
        RECT 68.065 65.365 68.365 65.845 ;
        RECT 68.625 65.365 69.835 66.115 ;
        RECT 70.005 65.365 70.295 66.090 ;
        RECT 70.465 65.365 72.135 66.135 ;
        RECT 72.805 65.365 73.035 66.185 ;
        RECT 73.285 66.165 73.535 66.765 ;
        RECT 73.205 65.535 73.535 66.165 ;
        RECT 73.705 65.365 73.915 66.185 ;
        RECT 75.730 65.910 76.070 66.740 ;
        RECT 77.550 66.230 77.900 67.480 ;
        RECT 79.665 66.825 83.175 67.915 ;
        RECT 79.665 66.135 81.315 66.655 ;
        RECT 81.485 66.305 83.175 66.825 ;
        RECT 84.470 66.945 84.800 67.745 ;
        RECT 84.970 67.115 85.300 67.915 ;
        RECT 85.600 66.945 85.930 67.745 ;
        RECT 86.575 67.115 86.825 67.915 ;
        RECT 84.470 66.775 86.905 66.945 ;
        RECT 87.095 66.775 87.265 67.915 ;
        RECT 87.435 66.775 87.775 67.745 ;
        RECT 87.945 66.825 90.535 67.915 ;
        RECT 84.265 66.355 84.615 66.605 ;
        RECT 84.800 66.145 84.970 66.775 ;
        RECT 85.140 66.355 85.470 66.555 ;
        RECT 85.640 66.355 85.970 66.555 ;
        RECT 86.140 66.355 86.560 66.555 ;
        RECT 86.735 66.525 86.905 66.775 ;
        RECT 86.735 66.355 87.430 66.525 ;
        RECT 74.145 65.365 79.490 65.910 ;
        RECT 79.665 65.365 83.175 66.135 ;
        RECT 84.470 65.535 84.970 66.145 ;
        RECT 85.600 66.015 86.825 66.185 ;
        RECT 87.600 66.165 87.775 66.775 ;
        RECT 85.600 65.535 85.930 66.015 ;
        RECT 86.100 65.365 86.325 65.825 ;
        RECT 86.495 65.535 86.825 66.015 ;
        RECT 87.015 65.365 87.265 66.165 ;
        RECT 87.435 65.535 87.775 66.165 ;
        RECT 87.945 66.135 89.155 66.655 ;
        RECT 89.325 66.305 90.535 66.825 ;
        RECT 90.910 66.945 91.240 67.745 ;
        RECT 91.410 67.115 91.740 67.915 ;
        RECT 92.040 66.945 92.370 67.745 ;
        RECT 93.015 67.115 93.265 67.915 ;
        RECT 90.910 66.775 93.345 66.945 ;
        RECT 93.535 66.775 93.705 67.915 ;
        RECT 93.875 66.775 94.215 67.745 ;
        RECT 94.425 66.775 94.655 67.915 ;
        RECT 90.705 66.355 91.055 66.605 ;
        RECT 91.240 66.145 91.410 66.775 ;
        RECT 91.580 66.355 91.910 66.555 ;
        RECT 92.080 66.355 92.410 66.555 ;
        RECT 92.580 66.355 93.000 66.555 ;
        RECT 93.175 66.525 93.345 66.775 ;
        RECT 93.175 66.355 93.870 66.525 ;
        RECT 87.945 65.365 90.535 66.135 ;
        RECT 90.910 65.535 91.410 66.145 ;
        RECT 92.040 66.015 93.265 66.185 ;
        RECT 94.040 66.165 94.215 66.775 ;
        RECT 94.825 66.765 95.155 67.745 ;
        RECT 95.325 66.775 95.535 67.915 ;
        RECT 94.405 66.355 94.735 66.605 ;
        RECT 92.040 65.535 92.370 66.015 ;
        RECT 92.540 65.365 92.765 65.825 ;
        RECT 92.935 65.535 93.265 66.015 ;
        RECT 93.455 65.365 93.705 66.165 ;
        RECT 93.875 65.535 94.215 66.165 ;
        RECT 94.425 65.365 94.655 66.185 ;
        RECT 94.905 66.165 95.155 66.765 ;
        RECT 95.765 66.750 96.055 67.915 ;
        RECT 96.430 66.945 96.760 67.745 ;
        RECT 96.930 67.115 97.260 67.915 ;
        RECT 97.560 66.945 97.890 67.745 ;
        RECT 98.535 67.115 98.785 67.915 ;
        RECT 96.430 66.775 98.865 66.945 ;
        RECT 99.055 66.775 99.225 67.915 ;
        RECT 99.395 66.775 99.735 67.745 ;
        RECT 99.995 67.245 100.165 67.745 ;
        RECT 100.335 67.415 100.665 67.915 ;
        RECT 99.995 67.075 100.660 67.245 ;
        RECT 96.225 66.355 96.575 66.605 ;
        RECT 94.825 65.535 95.155 66.165 ;
        RECT 95.325 65.365 95.535 66.185 ;
        RECT 96.760 66.145 96.930 66.775 ;
        RECT 97.100 66.355 97.430 66.555 ;
        RECT 97.600 66.355 97.930 66.555 ;
        RECT 98.100 66.355 98.520 66.555 ;
        RECT 98.695 66.525 98.865 66.775 ;
        RECT 98.695 66.355 99.390 66.525 ;
        RECT 95.765 65.365 96.055 66.090 ;
        RECT 96.430 65.535 96.930 66.145 ;
        RECT 97.560 66.015 98.785 66.185 ;
        RECT 99.560 66.165 99.735 66.775 ;
        RECT 99.910 66.255 100.260 66.905 ;
        RECT 97.560 65.535 97.890 66.015 ;
        RECT 98.060 65.365 98.285 65.825 ;
        RECT 98.455 65.535 98.785 66.015 ;
        RECT 98.975 65.365 99.225 66.165 ;
        RECT 99.395 65.535 99.735 66.165 ;
        RECT 100.430 66.085 100.660 67.075 ;
        RECT 99.995 65.915 100.660 66.085 ;
        RECT 99.995 65.625 100.165 65.915 ;
        RECT 100.335 65.365 100.665 65.745 ;
        RECT 100.835 65.625 101.060 67.745 ;
        RECT 101.275 67.415 101.605 67.915 ;
        RECT 101.775 67.245 101.945 67.745 ;
        RECT 102.180 67.530 103.010 67.700 ;
        RECT 103.250 67.535 103.630 67.915 ;
        RECT 101.250 67.075 101.945 67.245 ;
        RECT 101.250 66.105 101.420 67.075 ;
        RECT 101.590 66.285 102.000 66.905 ;
        RECT 102.170 66.855 102.670 67.235 ;
        RECT 101.250 65.915 101.945 66.105 ;
        RECT 102.170 65.985 102.390 66.855 ;
        RECT 102.840 66.685 103.010 67.530 ;
        RECT 103.810 67.365 103.980 67.655 ;
        RECT 104.150 67.535 104.480 67.915 ;
        RECT 104.950 67.445 105.580 67.695 ;
        RECT 105.760 67.535 106.180 67.915 ;
        RECT 105.410 67.365 105.580 67.445 ;
        RECT 106.380 67.365 106.620 67.655 ;
        RECT 103.180 67.115 104.550 67.365 ;
        RECT 103.180 66.855 103.430 67.115 ;
        RECT 103.940 66.685 104.190 66.845 ;
        RECT 102.840 66.515 104.190 66.685 ;
        RECT 102.840 66.475 103.260 66.515 ;
        RECT 102.570 65.925 102.920 66.295 ;
        RECT 101.275 65.365 101.605 65.745 ;
        RECT 101.775 65.585 101.945 65.915 ;
        RECT 103.090 65.745 103.260 66.475 ;
        RECT 104.360 66.345 104.550 67.115 ;
        RECT 103.430 66.015 103.840 66.345 ;
        RECT 104.130 66.005 104.550 66.345 ;
        RECT 104.720 66.935 105.240 67.245 ;
        RECT 105.410 67.195 106.620 67.365 ;
        RECT 106.850 67.225 107.180 67.915 ;
        RECT 104.720 66.175 104.890 66.935 ;
        RECT 105.060 66.345 105.240 66.755 ;
        RECT 105.410 66.685 105.580 67.195 ;
        RECT 107.350 67.045 107.520 67.655 ;
        RECT 107.790 67.195 108.120 67.705 ;
        RECT 107.350 67.025 107.670 67.045 ;
        RECT 105.750 66.855 107.670 67.025 ;
        RECT 105.410 66.515 107.310 66.685 ;
        RECT 105.640 66.175 105.970 66.295 ;
        RECT 104.720 66.005 105.970 66.175 ;
        RECT 102.245 65.545 103.260 65.745 ;
        RECT 103.430 65.365 103.840 65.805 ;
        RECT 104.130 65.575 104.380 66.005 ;
        RECT 104.580 65.365 104.900 65.825 ;
        RECT 106.140 65.755 106.310 66.515 ;
        RECT 106.980 66.455 107.310 66.515 ;
        RECT 106.500 66.285 106.830 66.345 ;
        RECT 106.500 66.015 107.160 66.285 ;
        RECT 107.480 65.960 107.670 66.855 ;
        RECT 105.460 65.585 106.310 65.755 ;
        RECT 106.510 65.365 107.170 65.845 ;
        RECT 107.350 65.630 107.670 65.960 ;
        RECT 107.870 66.605 108.120 67.195 ;
        RECT 108.300 67.115 108.585 67.915 ;
        RECT 108.765 66.935 109.020 67.605 ;
        RECT 107.870 66.275 108.670 66.605 ;
        RECT 107.870 65.625 108.120 66.275 ;
        RECT 108.840 66.075 109.020 66.935 ;
        RECT 109.605 66.775 109.835 67.915 ;
        RECT 110.005 66.765 110.335 67.745 ;
        RECT 110.505 66.775 110.715 67.915 ;
        RECT 110.945 66.825 112.155 67.915 ;
        RECT 109.585 66.355 109.915 66.605 ;
        RECT 108.765 65.875 109.020 66.075 ;
        RECT 108.300 65.365 108.585 65.825 ;
        RECT 108.765 65.705 109.105 65.875 ;
        RECT 108.765 65.545 109.020 65.705 ;
        RECT 109.605 65.365 109.835 66.185 ;
        RECT 110.085 66.165 110.335 66.765 ;
        RECT 110.005 65.535 110.335 66.165 ;
        RECT 110.505 65.365 110.715 66.185 ;
        RECT 110.945 66.115 111.465 66.655 ;
        RECT 111.635 66.285 112.155 66.825 ;
        RECT 112.325 66.825 113.535 67.915 ;
        RECT 112.325 66.285 112.845 66.825 ;
        RECT 113.015 66.115 113.535 66.655 ;
        RECT 110.945 65.365 112.155 66.115 ;
        RECT 112.325 65.365 113.535 66.115 ;
        RECT 5.520 65.195 113.620 65.365 ;
        RECT 5.605 64.445 6.815 65.195 ;
        RECT 7.075 64.645 7.245 64.935 ;
        RECT 7.415 64.815 7.745 65.195 ;
        RECT 7.075 64.475 7.740 64.645 ;
        RECT 5.605 63.905 6.125 64.445 ;
        RECT 6.295 63.735 6.815 64.275 ;
        RECT 5.605 62.645 6.815 63.735 ;
        RECT 6.990 63.655 7.340 64.305 ;
        RECT 7.510 63.485 7.740 64.475 ;
        RECT 7.075 63.315 7.740 63.485 ;
        RECT 7.075 62.815 7.245 63.315 ;
        RECT 7.415 62.645 7.745 63.145 ;
        RECT 7.915 62.815 8.140 64.935 ;
        RECT 8.355 64.815 8.685 65.195 ;
        RECT 8.855 64.645 9.025 64.975 ;
        RECT 9.325 64.815 10.340 65.015 ;
        RECT 8.330 64.455 9.025 64.645 ;
        RECT 8.330 63.485 8.500 64.455 ;
        RECT 8.670 63.655 9.080 64.275 ;
        RECT 9.250 63.705 9.470 64.575 ;
        RECT 9.650 64.265 10.000 64.635 ;
        RECT 10.170 64.085 10.340 64.815 ;
        RECT 10.510 64.755 10.920 65.195 ;
        RECT 11.210 64.555 11.460 64.985 ;
        RECT 11.660 64.735 11.980 65.195 ;
        RECT 12.540 64.805 13.390 64.975 ;
        RECT 10.510 64.215 10.920 64.545 ;
        RECT 11.210 64.215 11.630 64.555 ;
        RECT 9.920 64.045 10.340 64.085 ;
        RECT 9.920 63.875 11.270 64.045 ;
        RECT 8.330 63.315 9.025 63.485 ;
        RECT 9.250 63.325 9.750 63.705 ;
        RECT 8.355 62.645 8.685 63.145 ;
        RECT 8.855 62.815 9.025 63.315 ;
        RECT 9.920 63.030 10.090 63.875 ;
        RECT 11.020 63.715 11.270 63.875 ;
        RECT 10.260 63.445 10.510 63.705 ;
        RECT 11.440 63.445 11.630 64.215 ;
        RECT 10.260 63.195 11.630 63.445 ;
        RECT 11.800 64.385 13.050 64.555 ;
        RECT 11.800 63.625 11.970 64.385 ;
        RECT 12.720 64.265 13.050 64.385 ;
        RECT 12.140 63.805 12.320 64.215 ;
        RECT 13.220 64.045 13.390 64.805 ;
        RECT 13.590 64.715 14.250 65.195 ;
        RECT 14.430 64.600 14.750 64.930 ;
        RECT 13.580 64.275 14.240 64.545 ;
        RECT 13.580 64.215 13.910 64.275 ;
        RECT 14.060 64.045 14.390 64.105 ;
        RECT 12.490 63.875 14.390 64.045 ;
        RECT 11.800 63.315 12.320 63.625 ;
        RECT 12.490 63.365 12.660 63.875 ;
        RECT 14.560 63.705 14.750 64.600 ;
        RECT 12.830 63.535 14.750 63.705 ;
        RECT 14.430 63.515 14.750 63.535 ;
        RECT 14.950 64.285 15.200 64.935 ;
        RECT 15.380 64.735 15.665 65.195 ;
        RECT 15.845 64.855 16.100 65.015 ;
        RECT 15.845 64.685 16.185 64.855 ;
        RECT 15.845 64.485 16.100 64.685 ;
        RECT 14.950 63.955 15.750 64.285 ;
        RECT 12.490 63.195 13.700 63.365 ;
        RECT 9.260 62.860 10.090 63.030 ;
        RECT 10.330 62.645 10.710 63.025 ;
        RECT 10.890 62.905 11.060 63.195 ;
        RECT 12.490 63.115 12.660 63.195 ;
        RECT 11.230 62.645 11.560 63.025 ;
        RECT 12.030 62.865 12.660 63.115 ;
        RECT 12.840 62.645 13.260 63.025 ;
        RECT 13.460 62.905 13.700 63.195 ;
        RECT 13.930 62.645 14.260 63.335 ;
        RECT 14.430 62.905 14.600 63.515 ;
        RECT 14.950 63.365 15.200 63.955 ;
        RECT 15.920 63.625 16.100 64.485 ;
        RECT 16.705 64.375 16.915 65.195 ;
        RECT 17.085 64.395 17.415 65.025 ;
        RECT 17.085 63.795 17.335 64.395 ;
        RECT 17.585 64.375 17.815 65.195 ;
        RECT 18.025 64.425 20.615 65.195 ;
        RECT 17.505 63.955 17.835 64.205 ;
        RECT 18.025 63.905 19.235 64.425 ;
        RECT 20.785 64.395 21.125 65.025 ;
        RECT 21.295 64.395 21.545 65.195 ;
        RECT 21.735 64.545 22.065 65.025 ;
        RECT 22.235 64.735 22.460 65.195 ;
        RECT 22.630 64.545 22.960 65.025 ;
        RECT 14.870 62.855 15.200 63.365 ;
        RECT 15.380 62.645 15.665 63.445 ;
        RECT 15.845 62.955 16.100 63.625 ;
        RECT 16.705 62.645 16.915 63.785 ;
        RECT 17.085 62.815 17.415 63.795 ;
        RECT 17.585 62.645 17.815 63.785 ;
        RECT 19.405 63.735 20.615 64.255 ;
        RECT 18.025 62.645 20.615 63.735 ;
        RECT 20.785 63.785 20.960 64.395 ;
        RECT 21.735 64.375 22.960 64.545 ;
        RECT 23.590 64.415 24.090 65.025 ;
        RECT 24.670 64.415 25.170 65.025 ;
        RECT 21.130 64.035 21.825 64.205 ;
        RECT 21.655 63.785 21.825 64.035 ;
        RECT 22.000 64.005 22.420 64.205 ;
        RECT 22.590 64.005 22.920 64.205 ;
        RECT 23.090 64.005 23.420 64.205 ;
        RECT 23.590 63.785 23.760 64.415 ;
        RECT 23.945 63.955 24.295 64.205 ;
        RECT 24.465 63.955 24.815 64.205 ;
        RECT 25.000 63.785 25.170 64.415 ;
        RECT 25.800 64.545 26.130 65.025 ;
        RECT 26.300 64.735 26.525 65.195 ;
        RECT 26.695 64.545 27.025 65.025 ;
        RECT 25.800 64.375 27.025 64.545 ;
        RECT 27.215 64.395 27.465 65.195 ;
        RECT 27.635 64.395 27.975 65.025 ;
        RECT 25.340 64.005 25.670 64.205 ;
        RECT 25.840 64.005 26.170 64.205 ;
        RECT 26.340 64.005 26.760 64.205 ;
        RECT 26.935 64.035 27.630 64.205 ;
        RECT 26.935 63.785 27.105 64.035 ;
        RECT 27.800 63.785 27.975 64.395 ;
        RECT 28.145 64.425 30.735 65.195 ;
        RECT 31.365 64.470 31.655 65.195 ;
        RECT 28.145 63.905 29.355 64.425 ;
        RECT 31.825 64.395 32.165 65.025 ;
        RECT 32.335 64.395 32.585 65.195 ;
        RECT 32.775 64.545 33.105 65.025 ;
        RECT 33.275 64.735 33.500 65.195 ;
        RECT 33.670 64.545 34.000 65.025 ;
        RECT 20.785 62.815 21.125 63.785 ;
        RECT 21.295 62.645 21.465 63.785 ;
        RECT 21.655 63.615 24.090 63.785 ;
        RECT 21.735 62.645 21.985 63.445 ;
        RECT 22.630 62.815 22.960 63.615 ;
        RECT 23.260 62.645 23.590 63.445 ;
        RECT 23.760 62.815 24.090 63.615 ;
        RECT 24.670 63.615 27.105 63.785 ;
        RECT 24.670 62.815 25.000 63.615 ;
        RECT 25.170 62.645 25.500 63.445 ;
        RECT 25.800 62.815 26.130 63.615 ;
        RECT 26.775 62.645 27.025 63.445 ;
        RECT 27.295 62.645 27.465 63.785 ;
        RECT 27.635 62.815 27.975 63.785 ;
        RECT 29.525 63.735 30.735 64.255 ;
        RECT 28.145 62.645 30.735 63.735 ;
        RECT 31.365 62.645 31.655 63.810 ;
        RECT 31.825 63.785 32.000 64.395 ;
        RECT 32.775 64.375 34.000 64.545 ;
        RECT 34.630 64.415 35.130 65.025 ;
        RECT 35.505 64.425 39.015 65.195 ;
        RECT 32.170 64.035 32.865 64.205 ;
        RECT 32.695 63.785 32.865 64.035 ;
        RECT 33.040 64.005 33.460 64.205 ;
        RECT 33.630 64.005 33.960 64.205 ;
        RECT 34.130 64.005 34.460 64.205 ;
        RECT 34.630 63.785 34.800 64.415 ;
        RECT 34.985 63.955 35.335 64.205 ;
        RECT 35.505 63.905 37.155 64.425 ;
        RECT 39.225 64.375 39.455 65.195 ;
        RECT 39.625 64.395 39.955 65.025 ;
        RECT 31.825 62.815 32.165 63.785 ;
        RECT 32.335 62.645 32.505 63.785 ;
        RECT 32.695 63.615 35.130 63.785 ;
        RECT 37.325 63.735 39.015 64.255 ;
        RECT 39.205 63.955 39.535 64.205 ;
        RECT 39.705 63.795 39.955 64.395 ;
        RECT 40.125 64.375 40.335 65.195 ;
        RECT 40.565 64.650 45.910 65.195 ;
        RECT 42.150 63.820 42.490 64.650 ;
        RECT 46.085 64.425 49.595 65.195 ;
        RECT 32.775 62.645 33.025 63.445 ;
        RECT 33.670 62.815 34.000 63.615 ;
        RECT 34.300 62.645 34.630 63.445 ;
        RECT 34.800 62.815 35.130 63.615 ;
        RECT 35.505 62.645 39.015 63.735 ;
        RECT 39.225 62.645 39.455 63.785 ;
        RECT 39.625 62.815 39.955 63.795 ;
        RECT 40.125 62.645 40.335 63.785 ;
        RECT 43.970 63.080 44.320 64.330 ;
        RECT 46.085 63.905 47.735 64.425 ;
        RECT 50.685 64.395 51.025 65.025 ;
        RECT 51.195 64.395 51.445 65.195 ;
        RECT 51.635 64.545 51.965 65.025 ;
        RECT 52.135 64.735 52.360 65.195 ;
        RECT 52.530 64.545 52.860 65.025 ;
        RECT 47.905 63.735 49.595 64.255 ;
        RECT 40.565 62.645 45.910 63.080 ;
        RECT 46.085 62.645 49.595 63.735 ;
        RECT 50.685 63.785 50.860 64.395 ;
        RECT 51.635 64.375 52.860 64.545 ;
        RECT 53.490 64.415 53.990 65.025 ;
        RECT 51.030 64.035 51.725 64.205 ;
        RECT 51.555 63.785 51.725 64.035 ;
        RECT 51.900 64.005 52.320 64.205 ;
        RECT 52.490 64.005 52.820 64.205 ;
        RECT 52.990 64.005 53.320 64.205 ;
        RECT 53.490 63.785 53.660 64.415 ;
        RECT 55.290 64.355 55.550 65.195 ;
        RECT 55.725 64.450 55.980 65.025 ;
        RECT 56.150 64.815 56.480 65.195 ;
        RECT 56.695 64.645 56.865 65.025 ;
        RECT 56.150 64.475 56.865 64.645 ;
        RECT 53.845 63.955 54.195 64.205 ;
        RECT 50.685 62.815 51.025 63.785 ;
        RECT 51.195 62.645 51.365 63.785 ;
        RECT 51.555 63.615 53.990 63.785 ;
        RECT 51.635 62.645 51.885 63.445 ;
        RECT 52.530 62.815 52.860 63.615 ;
        RECT 53.160 62.645 53.490 63.445 ;
        RECT 53.660 62.815 53.990 63.615 ;
        RECT 55.290 62.645 55.550 63.795 ;
        RECT 55.725 63.720 55.895 64.450 ;
        RECT 56.150 64.285 56.320 64.475 ;
        RECT 57.125 64.470 57.415 65.195 ;
        RECT 58.050 64.355 58.310 65.195 ;
        RECT 58.485 64.450 58.740 65.025 ;
        RECT 58.910 64.815 59.240 65.195 ;
        RECT 59.455 64.645 59.625 65.025 ;
        RECT 58.910 64.475 59.625 64.645 ;
        RECT 59.975 64.645 60.145 65.025 ;
        RECT 60.360 64.815 60.690 65.195 ;
        RECT 59.975 64.475 60.690 64.645 ;
        RECT 56.065 63.955 56.320 64.285 ;
        RECT 56.150 63.745 56.320 63.955 ;
        RECT 56.600 63.925 56.955 64.295 ;
        RECT 55.725 62.815 55.980 63.720 ;
        RECT 56.150 63.575 56.865 63.745 ;
        RECT 56.150 62.645 56.480 63.405 ;
        RECT 56.695 62.815 56.865 63.575 ;
        RECT 57.125 62.645 57.415 63.810 ;
        RECT 58.050 62.645 58.310 63.795 ;
        RECT 58.485 63.720 58.655 64.450 ;
        RECT 58.910 64.285 59.080 64.475 ;
        RECT 58.825 63.955 59.080 64.285 ;
        RECT 58.910 63.745 59.080 63.955 ;
        RECT 59.360 63.925 59.715 64.295 ;
        RECT 59.885 63.925 60.240 64.295 ;
        RECT 60.520 64.285 60.690 64.475 ;
        RECT 60.860 64.450 61.115 65.025 ;
        RECT 60.520 63.955 60.775 64.285 ;
        RECT 60.520 63.745 60.690 63.955 ;
        RECT 58.485 62.815 58.740 63.720 ;
        RECT 58.910 63.575 59.625 63.745 ;
        RECT 58.910 62.645 59.240 63.405 ;
        RECT 59.455 62.815 59.625 63.575 ;
        RECT 59.975 63.575 60.690 63.745 ;
        RECT 60.945 63.720 61.115 64.450 ;
        RECT 61.290 64.355 61.550 65.195 ;
        RECT 61.815 64.645 61.985 65.025 ;
        RECT 62.200 64.815 62.530 65.195 ;
        RECT 61.815 64.475 62.530 64.645 ;
        RECT 61.725 63.925 62.080 64.295 ;
        RECT 62.360 64.285 62.530 64.475 ;
        RECT 62.700 64.450 62.955 65.025 ;
        RECT 62.360 63.955 62.615 64.285 ;
        RECT 59.975 62.815 60.145 63.575 ;
        RECT 60.360 62.645 60.690 63.405 ;
        RECT 60.860 62.815 61.115 63.720 ;
        RECT 61.290 62.645 61.550 63.795 ;
        RECT 62.360 63.745 62.530 63.955 ;
        RECT 61.815 63.575 62.530 63.745 ;
        RECT 62.785 63.720 62.955 64.450 ;
        RECT 63.130 64.355 63.390 65.195 ;
        RECT 63.655 64.645 63.825 65.025 ;
        RECT 64.040 64.815 64.370 65.195 ;
        RECT 63.655 64.475 64.370 64.645 ;
        RECT 63.565 63.925 63.920 64.295 ;
        RECT 64.200 64.285 64.370 64.475 ;
        RECT 64.540 64.450 64.795 65.025 ;
        RECT 64.200 63.955 64.455 64.285 ;
        RECT 61.815 62.815 61.985 63.575 ;
        RECT 62.200 62.645 62.530 63.405 ;
        RECT 62.700 62.815 62.955 63.720 ;
        RECT 63.130 62.645 63.390 63.795 ;
        RECT 64.200 63.745 64.370 63.955 ;
        RECT 63.655 63.575 64.370 63.745 ;
        RECT 64.625 63.720 64.795 64.450 ;
        RECT 64.970 64.355 65.230 65.195 ;
        RECT 65.405 64.520 65.665 65.025 ;
        RECT 65.845 64.815 66.175 65.195 ;
        RECT 66.355 64.645 66.525 65.025 ;
        RECT 63.655 62.815 63.825 63.575 ;
        RECT 64.040 62.645 64.370 63.405 ;
        RECT 64.540 62.815 64.795 63.720 ;
        RECT 64.970 62.645 65.230 63.795 ;
        RECT 65.405 63.720 65.575 64.520 ;
        RECT 65.860 64.475 66.525 64.645 ;
        RECT 65.860 64.220 66.030 64.475 ;
        RECT 66.785 64.425 70.295 65.195 ;
        RECT 65.745 63.890 66.030 64.220 ;
        RECT 66.265 63.925 66.595 64.295 ;
        RECT 66.785 63.905 68.435 64.425 ;
        RECT 70.670 64.415 71.170 65.025 ;
        RECT 65.860 63.745 66.030 63.890 ;
        RECT 65.405 62.815 65.675 63.720 ;
        RECT 65.860 63.575 66.525 63.745 ;
        RECT 68.605 63.735 70.295 64.255 ;
        RECT 70.465 63.955 70.815 64.205 ;
        RECT 71.000 63.785 71.170 64.415 ;
        RECT 71.800 64.545 72.130 65.025 ;
        RECT 72.300 64.735 72.525 65.195 ;
        RECT 72.695 64.545 73.025 65.025 ;
        RECT 71.800 64.375 73.025 64.545 ;
        RECT 73.215 64.395 73.465 65.195 ;
        RECT 73.635 64.395 73.975 65.025 ;
        RECT 74.145 64.650 79.490 65.195 ;
        RECT 71.340 64.005 71.670 64.205 ;
        RECT 71.840 64.005 72.170 64.205 ;
        RECT 72.340 64.005 72.760 64.205 ;
        RECT 72.935 64.035 73.630 64.205 ;
        RECT 72.935 63.785 73.105 64.035 ;
        RECT 73.800 63.785 73.975 64.395 ;
        RECT 75.730 63.820 76.070 64.650 ;
        RECT 79.665 64.425 82.255 65.195 ;
        RECT 82.885 64.470 83.175 65.195 ;
        RECT 65.845 62.645 66.175 63.405 ;
        RECT 66.355 62.815 66.525 63.575 ;
        RECT 66.785 62.645 70.295 63.735 ;
        RECT 70.670 63.615 73.105 63.785 ;
        RECT 70.670 62.815 71.000 63.615 ;
        RECT 71.170 62.645 71.500 63.445 ;
        RECT 71.800 62.815 72.130 63.615 ;
        RECT 72.775 62.645 73.025 63.445 ;
        RECT 73.295 62.645 73.465 63.785 ;
        RECT 73.635 62.815 73.975 63.785 ;
        RECT 77.550 63.080 77.900 64.330 ;
        RECT 79.665 63.905 80.875 64.425 ;
        RECT 83.345 64.395 83.685 65.025 ;
        RECT 83.855 64.395 84.105 65.195 ;
        RECT 84.295 64.545 84.625 65.025 ;
        RECT 84.795 64.735 85.020 65.195 ;
        RECT 85.190 64.545 85.520 65.025 ;
        RECT 81.045 63.735 82.255 64.255 ;
        RECT 74.145 62.645 79.490 63.080 ;
        RECT 79.665 62.645 82.255 63.735 ;
        RECT 82.885 62.645 83.175 63.810 ;
        RECT 83.345 63.785 83.520 64.395 ;
        RECT 84.295 64.375 85.520 64.545 ;
        RECT 86.150 64.415 86.650 65.025 ;
        RECT 87.025 64.445 88.235 65.195 ;
        RECT 88.495 64.645 88.665 65.025 ;
        RECT 88.845 64.815 89.175 65.195 ;
        RECT 88.495 64.475 89.160 64.645 ;
        RECT 89.355 64.520 89.615 65.025 ;
        RECT 83.690 64.035 84.385 64.205 ;
        RECT 84.215 63.785 84.385 64.035 ;
        RECT 84.560 64.005 84.980 64.205 ;
        RECT 85.150 64.005 85.480 64.205 ;
        RECT 85.650 64.005 85.980 64.205 ;
        RECT 86.150 63.785 86.320 64.415 ;
        RECT 86.505 63.955 86.855 64.205 ;
        RECT 87.025 63.905 87.545 64.445 ;
        RECT 83.345 62.815 83.685 63.785 ;
        RECT 83.855 62.645 84.025 63.785 ;
        RECT 84.215 63.615 86.650 63.785 ;
        RECT 87.715 63.735 88.235 64.275 ;
        RECT 88.425 63.925 88.755 64.295 ;
        RECT 88.990 64.220 89.160 64.475 ;
        RECT 88.990 63.890 89.275 64.220 ;
        RECT 88.990 63.745 89.160 63.890 ;
        RECT 84.295 62.645 84.545 63.445 ;
        RECT 85.190 62.815 85.520 63.615 ;
        RECT 85.820 62.645 86.150 63.445 ;
        RECT 86.320 62.815 86.650 63.615 ;
        RECT 87.025 62.645 88.235 63.735 ;
        RECT 88.495 63.575 89.160 63.745 ;
        RECT 89.445 63.720 89.615 64.520 ;
        RECT 89.875 64.645 90.045 64.935 ;
        RECT 90.215 64.815 90.545 65.195 ;
        RECT 89.875 64.475 90.540 64.645 ;
        RECT 88.495 62.815 88.665 63.575 ;
        RECT 88.845 62.645 89.175 63.405 ;
        RECT 89.345 62.815 89.615 63.720 ;
        RECT 89.790 63.655 90.140 64.305 ;
        RECT 90.310 63.485 90.540 64.475 ;
        RECT 89.875 63.315 90.540 63.485 ;
        RECT 89.875 62.815 90.045 63.315 ;
        RECT 90.215 62.645 90.545 63.145 ;
        RECT 90.715 62.815 90.940 64.935 ;
        RECT 91.155 64.815 91.485 65.195 ;
        RECT 91.655 64.645 91.825 64.975 ;
        RECT 92.125 64.815 93.140 65.015 ;
        RECT 91.130 64.455 91.825 64.645 ;
        RECT 91.130 63.485 91.300 64.455 ;
        RECT 91.470 63.655 91.880 64.275 ;
        RECT 92.050 63.705 92.270 64.575 ;
        RECT 92.450 64.265 92.800 64.635 ;
        RECT 92.970 64.085 93.140 64.815 ;
        RECT 93.310 64.755 93.720 65.195 ;
        RECT 94.010 64.555 94.260 64.985 ;
        RECT 94.460 64.735 94.780 65.195 ;
        RECT 95.340 64.805 96.190 64.975 ;
        RECT 93.310 64.215 93.720 64.545 ;
        RECT 94.010 64.215 94.430 64.555 ;
        RECT 92.720 64.045 93.140 64.085 ;
        RECT 92.720 63.875 94.070 64.045 ;
        RECT 91.130 63.315 91.825 63.485 ;
        RECT 92.050 63.325 92.550 63.705 ;
        RECT 91.155 62.645 91.485 63.145 ;
        RECT 91.655 62.815 91.825 63.315 ;
        RECT 92.720 63.030 92.890 63.875 ;
        RECT 93.820 63.715 94.070 63.875 ;
        RECT 93.060 63.445 93.310 63.705 ;
        RECT 94.240 63.445 94.430 64.215 ;
        RECT 93.060 63.195 94.430 63.445 ;
        RECT 94.600 64.385 95.850 64.555 ;
        RECT 94.600 63.625 94.770 64.385 ;
        RECT 95.520 64.265 95.850 64.385 ;
        RECT 94.940 63.805 95.120 64.215 ;
        RECT 96.020 64.045 96.190 64.805 ;
        RECT 96.390 64.715 97.050 65.195 ;
        RECT 97.230 64.600 97.550 64.930 ;
        RECT 96.380 64.275 97.040 64.545 ;
        RECT 96.380 64.215 96.710 64.275 ;
        RECT 96.860 64.045 97.190 64.105 ;
        RECT 95.290 63.875 97.190 64.045 ;
        RECT 94.600 63.315 95.120 63.625 ;
        RECT 95.290 63.365 95.460 63.875 ;
        RECT 97.360 63.705 97.550 64.600 ;
        RECT 95.630 63.535 97.550 63.705 ;
        RECT 97.230 63.515 97.550 63.535 ;
        RECT 97.750 64.285 98.000 64.935 ;
        RECT 98.180 64.735 98.465 65.195 ;
        RECT 98.645 64.485 98.900 65.015 ;
        RECT 97.750 63.955 98.550 64.285 ;
        RECT 95.290 63.195 96.500 63.365 ;
        RECT 92.060 62.860 92.890 63.030 ;
        RECT 93.130 62.645 93.510 63.025 ;
        RECT 93.690 62.905 93.860 63.195 ;
        RECT 95.290 63.115 95.460 63.195 ;
        RECT 94.030 62.645 94.360 63.025 ;
        RECT 94.830 62.865 95.460 63.115 ;
        RECT 95.640 62.645 96.060 63.025 ;
        RECT 96.260 62.905 96.500 63.195 ;
        RECT 96.730 62.645 97.060 63.335 ;
        RECT 97.230 62.905 97.400 63.515 ;
        RECT 97.750 63.365 98.000 63.955 ;
        RECT 98.720 63.835 98.900 64.485 ;
        RECT 99.450 64.455 99.705 65.025 ;
        RECT 99.875 64.795 100.205 65.195 ;
        RECT 100.630 64.660 101.160 65.025 ;
        RECT 100.630 64.625 100.805 64.660 ;
        RECT 99.875 64.455 100.805 64.625 ;
        RECT 98.720 63.665 98.985 63.835 ;
        RECT 99.450 63.785 99.620 64.455 ;
        RECT 99.875 64.285 100.045 64.455 ;
        RECT 99.790 63.955 100.045 64.285 ;
        RECT 100.270 63.955 100.465 64.285 ;
        RECT 98.720 63.625 98.900 63.665 ;
        RECT 97.670 62.855 98.000 63.365 ;
        RECT 98.180 62.645 98.465 63.445 ;
        RECT 98.645 62.955 98.900 63.625 ;
        RECT 99.450 62.815 99.785 63.785 ;
        RECT 99.955 62.645 100.125 63.785 ;
        RECT 100.295 62.985 100.465 63.955 ;
        RECT 100.635 63.325 100.805 64.455 ;
        RECT 100.975 63.665 101.145 64.465 ;
        RECT 101.350 64.175 101.625 65.025 ;
        RECT 101.345 64.005 101.625 64.175 ;
        RECT 101.350 63.865 101.625 64.005 ;
        RECT 101.795 63.665 101.985 65.025 ;
        RECT 102.165 64.660 102.675 65.195 ;
        RECT 102.895 64.385 103.140 64.990 ;
        RECT 103.590 64.455 103.845 65.025 ;
        RECT 104.015 64.795 104.345 65.195 ;
        RECT 104.770 64.660 105.300 65.025 ;
        RECT 104.770 64.625 104.945 64.660 ;
        RECT 104.015 64.455 104.945 64.625 ;
        RECT 105.490 64.515 105.765 65.025 ;
        RECT 102.185 64.215 103.415 64.385 ;
        RECT 100.975 63.495 101.985 63.665 ;
        RECT 102.155 63.650 102.905 63.840 ;
        RECT 100.635 63.155 101.760 63.325 ;
        RECT 102.155 62.985 102.325 63.650 ;
        RECT 103.075 63.405 103.415 64.215 ;
        RECT 100.295 62.815 102.325 62.985 ;
        RECT 102.495 62.645 102.665 63.405 ;
        RECT 102.900 62.995 103.415 63.405 ;
        RECT 103.590 63.785 103.760 64.455 ;
        RECT 104.015 64.285 104.185 64.455 ;
        RECT 103.930 63.955 104.185 64.285 ;
        RECT 104.410 63.955 104.605 64.285 ;
        RECT 103.590 62.815 103.925 63.785 ;
        RECT 104.095 62.645 104.265 63.785 ;
        RECT 104.435 62.985 104.605 63.955 ;
        RECT 104.775 63.325 104.945 64.455 ;
        RECT 105.115 63.665 105.285 64.465 ;
        RECT 105.485 64.345 105.765 64.515 ;
        RECT 105.490 63.865 105.765 64.345 ;
        RECT 105.935 63.665 106.125 65.025 ;
        RECT 106.305 64.660 106.815 65.195 ;
        RECT 107.035 64.385 107.280 64.990 ;
        RECT 108.645 64.470 108.935 65.195 ;
        RECT 109.105 64.425 111.695 65.195 ;
        RECT 112.325 64.445 113.535 65.195 ;
        RECT 106.325 64.215 107.555 64.385 ;
        RECT 105.115 63.495 106.125 63.665 ;
        RECT 106.295 63.650 107.045 63.840 ;
        RECT 104.775 63.155 105.900 63.325 ;
        RECT 106.295 62.985 106.465 63.650 ;
        RECT 107.215 63.405 107.555 64.215 ;
        RECT 109.105 63.905 110.315 64.425 ;
        RECT 104.435 62.815 106.465 62.985 ;
        RECT 106.635 62.645 106.805 63.405 ;
        RECT 107.040 62.995 107.555 63.405 ;
        RECT 108.645 62.645 108.935 63.810 ;
        RECT 110.485 63.735 111.695 64.255 ;
        RECT 109.105 62.645 111.695 63.735 ;
        RECT 112.325 63.735 112.845 64.275 ;
        RECT 113.015 63.905 113.535 64.445 ;
        RECT 112.325 62.645 113.535 63.735 ;
        RECT 5.520 62.475 113.620 62.645 ;
        RECT 5.605 61.385 6.815 62.475 ;
        RECT 7.910 61.805 8.165 62.305 ;
        RECT 8.335 61.975 8.665 62.475 ;
        RECT 7.910 61.635 8.660 61.805 ;
        RECT 5.605 60.675 6.125 61.215 ;
        RECT 6.295 60.845 6.815 61.385 ;
        RECT 7.910 60.815 8.260 61.465 ;
        RECT 5.605 59.925 6.815 60.675 ;
        RECT 8.430 60.645 8.660 61.635 ;
        RECT 7.910 60.475 8.660 60.645 ;
        RECT 7.910 60.185 8.165 60.475 ;
        RECT 8.335 59.925 8.665 60.305 ;
        RECT 8.835 60.185 9.005 62.305 ;
        RECT 9.175 61.505 9.500 62.290 ;
        RECT 9.670 62.015 9.920 62.475 ;
        RECT 10.090 61.975 10.340 62.305 ;
        RECT 10.555 61.975 11.235 62.305 ;
        RECT 10.090 61.845 10.260 61.975 ;
        RECT 9.865 61.675 10.260 61.845 ;
        RECT 9.235 60.455 9.695 61.505 ;
        RECT 9.865 60.315 10.035 61.675 ;
        RECT 10.430 61.415 10.895 61.805 ;
        RECT 10.205 60.605 10.555 61.225 ;
        RECT 10.725 60.825 10.895 61.415 ;
        RECT 11.065 61.195 11.235 61.975 ;
        RECT 11.405 61.875 11.575 62.215 ;
        RECT 11.810 62.045 12.140 62.475 ;
        RECT 12.310 61.875 12.480 62.215 ;
        RECT 12.775 62.015 13.145 62.475 ;
        RECT 11.405 61.705 12.480 61.875 ;
        RECT 13.315 61.845 13.485 62.305 ;
        RECT 13.720 61.965 14.590 62.305 ;
        RECT 14.760 62.015 15.010 62.475 ;
        RECT 12.925 61.675 13.485 61.845 ;
        RECT 12.925 61.535 13.095 61.675 ;
        RECT 11.595 61.365 13.095 61.535 ;
        RECT 13.790 61.505 14.250 61.795 ;
        RECT 11.065 61.025 12.755 61.195 ;
        RECT 10.725 60.605 11.080 60.825 ;
        RECT 11.250 60.315 11.420 61.025 ;
        RECT 11.625 60.605 12.415 60.855 ;
        RECT 12.585 60.845 12.755 61.025 ;
        RECT 12.925 60.675 13.095 61.365 ;
        RECT 9.365 59.925 9.695 60.285 ;
        RECT 9.865 60.145 10.360 60.315 ;
        RECT 10.565 60.145 11.420 60.315 ;
        RECT 12.295 59.925 12.625 60.385 ;
        RECT 12.835 60.285 13.095 60.675 ;
        RECT 13.285 61.495 14.250 61.505 ;
        RECT 14.420 61.585 14.590 61.965 ;
        RECT 15.180 61.925 15.350 62.215 ;
        RECT 15.530 62.095 15.860 62.475 ;
        RECT 15.180 61.755 15.980 61.925 ;
        RECT 13.285 61.335 13.960 61.495 ;
        RECT 14.420 61.415 15.640 61.585 ;
        RECT 13.285 60.545 13.495 61.335 ;
        RECT 14.420 61.325 14.590 61.415 ;
        RECT 13.665 60.545 14.015 61.165 ;
        RECT 14.185 61.155 14.590 61.325 ;
        RECT 14.185 60.375 14.355 61.155 ;
        RECT 14.525 60.705 14.745 60.985 ;
        RECT 14.925 60.875 15.465 61.245 ;
        RECT 15.810 61.165 15.980 61.755 ;
        RECT 16.200 61.335 16.505 62.475 ;
        RECT 16.675 61.285 16.930 62.165 ;
        RECT 17.105 61.385 18.315 62.475 ;
        RECT 15.810 61.135 16.550 61.165 ;
        RECT 14.525 60.535 15.055 60.705 ;
        RECT 12.835 60.115 13.185 60.285 ;
        RECT 13.405 60.095 14.355 60.375 ;
        RECT 14.525 59.925 14.715 60.365 ;
        RECT 14.885 60.305 15.055 60.535 ;
        RECT 15.225 60.475 15.465 60.875 ;
        RECT 15.635 60.835 16.550 61.135 ;
        RECT 15.635 60.660 15.960 60.835 ;
        RECT 15.635 60.305 15.955 60.660 ;
        RECT 16.720 60.635 16.930 61.285 ;
        RECT 14.885 60.135 15.955 60.305 ;
        RECT 16.200 59.925 16.505 60.385 ;
        RECT 16.675 60.105 16.930 60.635 ;
        RECT 17.105 60.675 17.625 61.215 ;
        RECT 17.795 60.845 18.315 61.385 ;
        RECT 18.485 61.310 18.775 62.475 ;
        RECT 18.945 61.385 20.615 62.475 ;
        RECT 18.945 60.695 19.695 61.215 ;
        RECT 19.865 60.865 20.615 61.385 ;
        RECT 21.450 61.505 21.780 62.305 ;
        RECT 21.950 61.675 22.280 62.475 ;
        RECT 22.580 61.505 22.910 62.305 ;
        RECT 23.555 61.675 23.805 62.475 ;
        RECT 21.450 61.335 23.885 61.505 ;
        RECT 24.075 61.335 24.245 62.475 ;
        RECT 24.415 61.335 24.755 62.305 ;
        RECT 24.925 62.040 30.270 62.475 ;
        RECT 30.445 62.040 35.790 62.475 ;
        RECT 35.965 62.040 41.310 62.475 ;
        RECT 21.245 60.915 21.595 61.165 ;
        RECT 21.780 60.705 21.950 61.335 ;
        RECT 22.120 60.915 22.450 61.115 ;
        RECT 22.620 60.915 22.950 61.115 ;
        RECT 23.120 60.915 23.540 61.115 ;
        RECT 23.715 61.085 23.885 61.335 ;
        RECT 23.715 60.915 24.410 61.085 ;
        RECT 17.105 59.925 18.315 60.675 ;
        RECT 18.485 59.925 18.775 60.650 ;
        RECT 18.945 59.925 20.615 60.695 ;
        RECT 21.450 60.095 21.950 60.705 ;
        RECT 22.580 60.575 23.805 60.745 ;
        RECT 24.580 60.725 24.755 61.335 ;
        RECT 22.580 60.095 22.910 60.575 ;
        RECT 23.080 59.925 23.305 60.385 ;
        RECT 23.475 60.095 23.805 60.575 ;
        RECT 23.995 59.925 24.245 60.725 ;
        RECT 24.415 60.095 24.755 60.725 ;
        RECT 26.510 60.470 26.850 61.300 ;
        RECT 28.330 60.790 28.680 62.040 ;
        RECT 32.030 60.470 32.370 61.300 ;
        RECT 33.850 60.790 34.200 62.040 ;
        RECT 37.550 60.470 37.890 61.300 ;
        RECT 39.370 60.790 39.720 62.040 ;
        RECT 41.485 61.385 44.075 62.475 ;
        RECT 41.485 60.695 42.695 61.215 ;
        RECT 42.865 60.865 44.075 61.385 ;
        RECT 44.245 61.310 44.535 62.475 ;
        RECT 44.795 61.805 44.965 62.305 ;
        RECT 45.135 61.975 45.465 62.475 ;
        RECT 44.795 61.635 45.460 61.805 ;
        RECT 44.710 60.815 45.060 61.465 ;
        RECT 24.925 59.925 30.270 60.470 ;
        RECT 30.445 59.925 35.790 60.470 ;
        RECT 35.965 59.925 41.310 60.470 ;
        RECT 41.485 59.925 44.075 60.695 ;
        RECT 44.245 59.925 44.535 60.650 ;
        RECT 45.230 60.645 45.460 61.635 ;
        RECT 44.795 60.475 45.460 60.645 ;
        RECT 44.795 60.185 44.965 60.475 ;
        RECT 45.135 59.925 45.465 60.305 ;
        RECT 45.635 60.185 45.860 62.305 ;
        RECT 46.075 61.975 46.405 62.475 ;
        RECT 46.575 61.805 46.745 62.305 ;
        RECT 46.980 62.090 47.810 62.260 ;
        RECT 48.050 62.095 48.430 62.475 ;
        RECT 46.050 61.635 46.745 61.805 ;
        RECT 46.050 60.665 46.220 61.635 ;
        RECT 46.390 60.845 46.800 61.465 ;
        RECT 46.970 61.415 47.470 61.795 ;
        RECT 46.050 60.475 46.745 60.665 ;
        RECT 46.970 60.545 47.190 61.415 ;
        RECT 47.640 61.245 47.810 62.090 ;
        RECT 48.610 61.925 48.780 62.215 ;
        RECT 48.950 62.095 49.280 62.475 ;
        RECT 49.750 62.005 50.380 62.255 ;
        RECT 50.560 62.095 50.980 62.475 ;
        RECT 50.210 61.925 50.380 62.005 ;
        RECT 51.180 61.925 51.420 62.215 ;
        RECT 47.980 61.675 49.350 61.925 ;
        RECT 47.980 61.415 48.230 61.675 ;
        RECT 48.740 61.245 48.990 61.405 ;
        RECT 47.640 61.075 48.990 61.245 ;
        RECT 47.640 61.035 48.060 61.075 ;
        RECT 47.370 60.485 47.720 60.855 ;
        RECT 46.075 59.925 46.405 60.305 ;
        RECT 46.575 60.145 46.745 60.475 ;
        RECT 47.890 60.305 48.060 61.035 ;
        RECT 49.160 60.905 49.350 61.675 ;
        RECT 48.230 60.575 48.640 60.905 ;
        RECT 48.930 60.565 49.350 60.905 ;
        RECT 49.520 61.495 50.040 61.805 ;
        RECT 50.210 61.755 51.420 61.925 ;
        RECT 51.650 61.785 51.980 62.475 ;
        RECT 49.520 60.735 49.690 61.495 ;
        RECT 49.860 60.905 50.040 61.315 ;
        RECT 50.210 61.245 50.380 61.755 ;
        RECT 52.150 61.605 52.320 62.215 ;
        RECT 52.590 61.755 52.920 62.265 ;
        RECT 52.150 61.585 52.470 61.605 ;
        RECT 50.550 61.415 52.470 61.585 ;
        RECT 50.210 61.075 52.110 61.245 ;
        RECT 50.440 60.735 50.770 60.855 ;
        RECT 49.520 60.565 50.770 60.735 ;
        RECT 47.045 60.105 48.060 60.305 ;
        RECT 48.230 59.925 48.640 60.365 ;
        RECT 48.930 60.135 49.180 60.565 ;
        RECT 49.380 59.925 49.700 60.385 ;
        RECT 50.940 60.315 51.110 61.075 ;
        RECT 51.780 61.015 52.110 61.075 ;
        RECT 51.300 60.845 51.630 60.905 ;
        RECT 51.300 60.575 51.960 60.845 ;
        RECT 52.280 60.520 52.470 61.415 ;
        RECT 50.260 60.145 51.110 60.315 ;
        RECT 51.310 59.925 51.970 60.405 ;
        RECT 52.150 60.190 52.470 60.520 ;
        RECT 52.670 61.165 52.920 61.755 ;
        RECT 53.100 61.675 53.385 62.475 ;
        RECT 53.565 61.495 53.820 62.165 ;
        RECT 52.670 60.835 53.470 61.165 ;
        RECT 52.670 60.185 52.920 60.835 ;
        RECT 53.640 60.635 53.820 61.495 ;
        RECT 53.565 60.435 53.820 60.635 ;
        RECT 54.365 61.335 54.705 62.305 ;
        RECT 54.875 61.335 55.045 62.475 ;
        RECT 55.315 61.675 55.565 62.475 ;
        RECT 56.210 61.505 56.540 62.305 ;
        RECT 56.840 61.675 57.170 62.475 ;
        RECT 57.340 61.505 57.670 62.305 ;
        RECT 55.235 61.335 57.670 61.505 ;
        RECT 58.045 61.385 59.715 62.475 ;
        RECT 54.365 60.725 54.540 61.335 ;
        RECT 55.235 61.085 55.405 61.335 ;
        RECT 54.710 60.915 55.405 61.085 ;
        RECT 55.580 60.915 56.000 61.115 ;
        RECT 56.170 60.915 56.500 61.115 ;
        RECT 56.670 60.915 57.000 61.115 ;
        RECT 53.100 59.925 53.385 60.385 ;
        RECT 53.565 60.265 53.905 60.435 ;
        RECT 53.565 60.105 53.820 60.265 ;
        RECT 54.365 60.095 54.705 60.725 ;
        RECT 54.875 59.925 55.125 60.725 ;
        RECT 55.315 60.575 56.540 60.745 ;
        RECT 55.315 60.095 55.645 60.575 ;
        RECT 55.815 59.925 56.040 60.385 ;
        RECT 56.210 60.095 56.540 60.575 ;
        RECT 57.170 60.705 57.340 61.335 ;
        RECT 57.525 60.915 57.875 61.165 ;
        RECT 57.170 60.095 57.670 60.705 ;
        RECT 58.045 60.695 58.795 61.215 ;
        RECT 58.965 60.865 59.715 61.385 ;
        RECT 59.975 61.545 60.145 62.305 ;
        RECT 60.360 61.715 60.690 62.475 ;
        RECT 59.975 61.375 60.690 61.545 ;
        RECT 60.860 61.400 61.115 62.305 ;
        RECT 59.885 60.825 60.240 61.195 ;
        RECT 60.520 61.165 60.690 61.375 ;
        RECT 60.520 60.835 60.775 61.165 ;
        RECT 58.045 59.925 59.715 60.695 ;
        RECT 60.520 60.645 60.690 60.835 ;
        RECT 60.945 60.670 61.115 61.400 ;
        RECT 61.290 61.325 61.550 62.475 ;
        RECT 61.815 61.545 61.985 62.305 ;
        RECT 62.200 61.715 62.530 62.475 ;
        RECT 61.815 61.375 62.530 61.545 ;
        RECT 62.700 61.400 62.955 62.305 ;
        RECT 61.725 60.825 62.080 61.195 ;
        RECT 62.360 61.165 62.530 61.375 ;
        RECT 62.360 60.835 62.615 61.165 ;
        RECT 59.975 60.475 60.690 60.645 ;
        RECT 59.975 60.095 60.145 60.475 ;
        RECT 60.360 59.925 60.690 60.305 ;
        RECT 60.860 60.095 61.115 60.670 ;
        RECT 61.290 59.925 61.550 60.765 ;
        RECT 62.360 60.645 62.530 60.835 ;
        RECT 62.785 60.670 62.955 61.400 ;
        RECT 63.130 61.325 63.390 62.475 ;
        RECT 64.490 61.335 64.825 62.305 ;
        RECT 64.995 61.335 65.165 62.475 ;
        RECT 65.335 62.135 67.365 62.305 ;
        RECT 61.815 60.475 62.530 60.645 ;
        RECT 61.815 60.095 61.985 60.475 ;
        RECT 62.200 59.925 62.530 60.305 ;
        RECT 62.700 60.095 62.955 60.670 ;
        RECT 63.130 59.925 63.390 60.765 ;
        RECT 64.490 60.665 64.660 61.335 ;
        RECT 65.335 61.165 65.505 62.135 ;
        RECT 64.830 60.835 65.085 61.165 ;
        RECT 65.310 60.835 65.505 61.165 ;
        RECT 65.675 61.795 66.800 61.965 ;
        RECT 64.915 60.665 65.085 60.835 ;
        RECT 65.675 60.665 65.845 61.795 ;
        RECT 64.490 60.095 64.745 60.665 ;
        RECT 64.915 60.495 65.845 60.665 ;
        RECT 66.015 61.455 67.025 61.625 ;
        RECT 66.015 60.655 66.185 61.455 ;
        RECT 65.670 60.460 65.845 60.495 ;
        RECT 64.915 59.925 65.245 60.325 ;
        RECT 65.670 60.095 66.200 60.460 ;
        RECT 66.390 60.435 66.665 61.255 ;
        RECT 66.385 60.265 66.665 60.435 ;
        RECT 66.390 60.095 66.665 60.265 ;
        RECT 66.835 60.095 67.025 61.455 ;
        RECT 67.195 61.470 67.365 62.135 ;
        RECT 67.535 61.715 67.705 62.475 ;
        RECT 67.940 61.715 68.455 62.125 ;
        RECT 67.195 61.280 67.945 61.470 ;
        RECT 68.115 60.905 68.455 61.715 ;
        RECT 68.715 61.545 68.885 62.305 ;
        RECT 69.065 61.715 69.395 62.475 ;
        RECT 68.715 61.375 69.380 61.545 ;
        RECT 69.565 61.400 69.835 62.305 ;
        RECT 69.210 61.230 69.380 61.375 ;
        RECT 67.225 60.735 68.455 60.905 ;
        RECT 68.645 60.825 68.975 61.195 ;
        RECT 69.210 60.900 69.495 61.230 ;
        RECT 67.205 59.925 67.715 60.460 ;
        RECT 67.935 60.130 68.180 60.735 ;
        RECT 69.210 60.645 69.380 60.900 ;
        RECT 68.715 60.475 69.380 60.645 ;
        RECT 69.665 60.600 69.835 61.400 ;
        RECT 70.005 61.310 70.295 62.475 ;
        RECT 70.465 62.040 75.810 62.475 ;
        RECT 68.715 60.095 68.885 60.475 ;
        RECT 69.065 59.925 69.395 60.305 ;
        RECT 69.575 60.095 69.835 60.600 ;
        RECT 70.005 59.925 70.295 60.650 ;
        RECT 72.050 60.470 72.390 61.300 ;
        RECT 73.870 60.790 74.220 62.040 ;
        RECT 76.190 61.505 76.520 62.305 ;
        RECT 76.690 61.675 77.020 62.475 ;
        RECT 77.320 61.505 77.650 62.305 ;
        RECT 78.295 61.675 78.545 62.475 ;
        RECT 76.190 61.335 78.625 61.505 ;
        RECT 78.815 61.335 78.985 62.475 ;
        RECT 79.155 61.335 79.495 62.305 ;
        RECT 75.985 60.915 76.335 61.165 ;
        RECT 76.520 60.705 76.690 61.335 ;
        RECT 76.860 60.915 77.190 61.115 ;
        RECT 77.360 60.915 77.690 61.115 ;
        RECT 77.860 60.915 78.280 61.115 ;
        RECT 78.455 61.085 78.625 61.335 ;
        RECT 78.455 60.915 79.150 61.085 ;
        RECT 70.465 59.925 75.810 60.470 ;
        RECT 76.190 60.095 76.690 60.705 ;
        RECT 77.320 60.575 78.545 60.745 ;
        RECT 79.320 60.725 79.495 61.335 ;
        RECT 77.320 60.095 77.650 60.575 ;
        RECT 77.820 59.925 78.045 60.385 ;
        RECT 78.215 60.095 78.545 60.575 ;
        RECT 78.735 59.925 78.985 60.725 ;
        RECT 79.155 60.095 79.495 60.725 ;
        RECT 79.665 61.335 80.005 62.305 ;
        RECT 80.175 61.335 80.345 62.475 ;
        RECT 80.615 61.675 80.865 62.475 ;
        RECT 81.510 61.505 81.840 62.305 ;
        RECT 82.140 61.675 82.470 62.475 ;
        RECT 82.640 61.505 82.970 62.305 ;
        RECT 80.535 61.335 82.970 61.505 ;
        RECT 83.345 61.335 83.685 62.305 ;
        RECT 83.855 61.335 84.025 62.475 ;
        RECT 84.295 61.675 84.545 62.475 ;
        RECT 85.190 61.505 85.520 62.305 ;
        RECT 85.820 61.675 86.150 62.475 ;
        RECT 86.320 61.505 86.650 62.305 ;
        RECT 84.215 61.335 86.650 61.505 ;
        RECT 87.025 61.385 90.535 62.475 ;
        RECT 79.665 61.285 79.895 61.335 ;
        RECT 79.665 60.725 79.840 61.285 ;
        RECT 80.535 61.085 80.705 61.335 ;
        RECT 80.010 60.915 80.705 61.085 ;
        RECT 80.880 60.915 81.300 61.115 ;
        RECT 81.470 60.915 81.800 61.115 ;
        RECT 81.970 60.915 82.300 61.115 ;
        RECT 79.665 60.095 80.005 60.725 ;
        RECT 80.175 59.925 80.425 60.725 ;
        RECT 80.615 60.575 81.840 60.745 ;
        RECT 80.615 60.095 80.945 60.575 ;
        RECT 81.115 59.925 81.340 60.385 ;
        RECT 81.510 60.095 81.840 60.575 ;
        RECT 82.470 60.705 82.640 61.335 ;
        RECT 83.345 61.285 83.575 61.335 ;
        RECT 82.825 60.915 83.175 61.165 ;
        RECT 83.345 60.725 83.520 61.285 ;
        RECT 84.215 61.085 84.385 61.335 ;
        RECT 83.690 60.915 84.385 61.085 ;
        RECT 84.555 60.945 84.980 61.115 ;
        RECT 84.560 60.915 84.980 60.945 ;
        RECT 85.150 60.915 85.480 61.115 ;
        RECT 85.650 60.915 85.980 61.115 ;
        RECT 82.470 60.095 82.970 60.705 ;
        RECT 83.345 60.095 83.685 60.725 ;
        RECT 83.855 59.925 84.105 60.725 ;
        RECT 84.295 60.575 85.520 60.745 ;
        RECT 84.295 60.095 84.625 60.575 ;
        RECT 84.795 59.925 85.020 60.385 ;
        RECT 85.190 60.095 85.520 60.575 ;
        RECT 86.150 60.705 86.320 61.335 ;
        RECT 86.505 60.915 86.855 61.165 ;
        RECT 86.150 60.095 86.650 60.705 ;
        RECT 87.025 60.695 88.675 61.215 ;
        RECT 88.845 60.865 90.535 61.385 ;
        RECT 90.710 61.335 91.045 62.305 ;
        RECT 91.215 61.335 91.385 62.475 ;
        RECT 91.555 62.135 93.585 62.305 ;
        RECT 87.025 59.925 90.535 60.695 ;
        RECT 90.710 60.665 90.880 61.335 ;
        RECT 91.555 61.165 91.725 62.135 ;
        RECT 91.050 60.835 91.305 61.165 ;
        RECT 91.530 60.835 91.725 61.165 ;
        RECT 91.895 61.795 93.020 61.965 ;
        RECT 91.135 60.665 91.305 60.835 ;
        RECT 91.895 60.665 92.065 61.795 ;
        RECT 90.710 60.095 90.965 60.665 ;
        RECT 91.135 60.495 92.065 60.665 ;
        RECT 92.235 61.455 93.245 61.625 ;
        RECT 92.235 60.655 92.405 61.455 ;
        RECT 91.890 60.460 92.065 60.495 ;
        RECT 91.135 59.925 91.465 60.325 ;
        RECT 91.890 60.095 92.420 60.460 ;
        RECT 92.610 60.435 92.885 61.255 ;
        RECT 92.605 60.265 92.885 60.435 ;
        RECT 92.610 60.095 92.885 60.265 ;
        RECT 93.055 60.095 93.245 61.455 ;
        RECT 93.415 61.470 93.585 62.135 ;
        RECT 93.755 61.715 93.925 62.475 ;
        RECT 94.160 61.715 94.675 62.125 ;
        RECT 93.415 61.280 94.165 61.470 ;
        RECT 94.335 60.905 94.675 61.715 ;
        RECT 95.765 61.310 96.055 62.475 ;
        RECT 96.225 62.040 101.570 62.475 ;
        RECT 93.445 60.735 94.675 60.905 ;
        RECT 93.425 59.925 93.935 60.460 ;
        RECT 94.155 60.130 94.400 60.735 ;
        RECT 95.765 59.925 96.055 60.650 ;
        RECT 97.810 60.470 98.150 61.300 ;
        RECT 99.630 60.790 99.980 62.040 ;
        RECT 102.295 61.805 102.465 62.305 ;
        RECT 102.635 61.975 102.965 62.475 ;
        RECT 102.295 61.635 102.960 61.805 ;
        RECT 102.210 60.815 102.560 61.465 ;
        RECT 102.730 60.645 102.960 61.635 ;
        RECT 102.295 60.475 102.960 60.645 ;
        RECT 96.225 59.925 101.570 60.470 ;
        RECT 102.295 60.185 102.465 60.475 ;
        RECT 102.635 59.925 102.965 60.305 ;
        RECT 103.135 60.185 103.360 62.305 ;
        RECT 103.575 61.975 103.905 62.475 ;
        RECT 104.075 61.805 104.245 62.305 ;
        RECT 104.480 62.090 105.310 62.260 ;
        RECT 105.550 62.095 105.930 62.475 ;
        RECT 103.550 61.635 104.245 61.805 ;
        RECT 103.550 60.665 103.720 61.635 ;
        RECT 103.890 60.845 104.300 61.465 ;
        RECT 104.470 61.415 104.970 61.795 ;
        RECT 103.550 60.475 104.245 60.665 ;
        RECT 104.470 60.545 104.690 61.415 ;
        RECT 105.140 61.245 105.310 62.090 ;
        RECT 106.110 61.925 106.280 62.215 ;
        RECT 106.450 62.095 106.780 62.475 ;
        RECT 107.250 62.005 107.880 62.255 ;
        RECT 108.060 62.095 108.480 62.475 ;
        RECT 107.710 61.925 107.880 62.005 ;
        RECT 108.680 61.925 108.920 62.215 ;
        RECT 105.480 61.675 106.850 61.925 ;
        RECT 105.480 61.415 105.730 61.675 ;
        RECT 106.240 61.245 106.490 61.405 ;
        RECT 105.140 61.075 106.490 61.245 ;
        RECT 105.140 61.035 105.560 61.075 ;
        RECT 104.870 60.485 105.220 60.855 ;
        RECT 103.575 59.925 103.905 60.305 ;
        RECT 104.075 60.145 104.245 60.475 ;
        RECT 105.390 60.305 105.560 61.035 ;
        RECT 106.660 60.905 106.850 61.675 ;
        RECT 105.730 60.575 106.140 60.905 ;
        RECT 106.430 60.565 106.850 60.905 ;
        RECT 107.020 61.495 107.540 61.805 ;
        RECT 107.710 61.755 108.920 61.925 ;
        RECT 109.150 61.785 109.480 62.475 ;
        RECT 107.020 60.735 107.190 61.495 ;
        RECT 107.360 60.905 107.540 61.315 ;
        RECT 107.710 61.245 107.880 61.755 ;
        RECT 109.650 61.605 109.820 62.215 ;
        RECT 110.090 61.755 110.420 62.265 ;
        RECT 109.650 61.585 109.970 61.605 ;
        RECT 108.050 61.415 109.970 61.585 ;
        RECT 107.710 61.075 109.610 61.245 ;
        RECT 107.940 60.735 108.270 60.855 ;
        RECT 107.020 60.565 108.270 60.735 ;
        RECT 104.545 60.105 105.560 60.305 ;
        RECT 105.730 59.925 106.140 60.365 ;
        RECT 106.430 60.135 106.680 60.565 ;
        RECT 106.880 59.925 107.200 60.385 ;
        RECT 108.440 60.315 108.610 61.075 ;
        RECT 109.280 61.015 109.610 61.075 ;
        RECT 108.800 60.845 109.130 60.905 ;
        RECT 108.800 60.575 109.460 60.845 ;
        RECT 109.780 60.520 109.970 61.415 ;
        RECT 107.760 60.145 108.610 60.315 ;
        RECT 108.810 59.925 109.470 60.405 ;
        RECT 109.650 60.190 109.970 60.520 ;
        RECT 110.170 61.165 110.420 61.755 ;
        RECT 110.600 61.675 110.885 62.475 ;
        RECT 111.065 62.135 111.320 62.165 ;
        RECT 111.065 61.965 111.405 62.135 ;
        RECT 111.065 61.495 111.320 61.965 ;
        RECT 110.170 60.835 110.970 61.165 ;
        RECT 110.170 60.185 110.420 60.835 ;
        RECT 111.140 60.635 111.320 61.495 ;
        RECT 112.325 61.385 113.535 62.475 ;
        RECT 112.325 60.845 112.845 61.385 ;
        RECT 113.015 60.675 113.535 61.215 ;
        RECT 110.600 59.925 110.885 60.385 ;
        RECT 111.065 60.105 111.320 60.635 ;
        RECT 112.325 59.925 113.535 60.675 ;
        RECT 5.520 59.755 113.620 59.925 ;
        RECT 5.605 59.005 6.815 59.755 ;
        RECT 6.985 59.210 12.330 59.755 ;
        RECT 5.605 58.465 6.125 59.005 ;
        RECT 6.295 58.295 6.815 58.835 ;
        RECT 8.570 58.380 8.910 59.210 ;
        RECT 12.505 59.005 13.715 59.755 ;
        RECT 5.605 57.205 6.815 58.295 ;
        RECT 10.390 57.640 10.740 58.890 ;
        RECT 12.505 58.465 13.025 59.005 ;
        RECT 14.035 58.955 14.365 59.755 ;
        RECT 14.535 59.105 14.705 59.585 ;
        RECT 14.875 59.275 15.205 59.755 ;
        RECT 15.375 59.105 15.545 59.585 ;
        RECT 15.795 59.275 16.035 59.755 ;
        RECT 16.215 59.105 16.385 59.585 ;
        RECT 16.645 59.210 21.990 59.755 ;
        RECT 14.535 58.935 15.545 59.105 ;
        RECT 15.750 58.935 16.385 59.105 ;
        RECT 14.535 58.905 15.035 58.935 ;
        RECT 13.195 58.295 13.715 58.835 ;
        RECT 14.535 58.395 15.030 58.905 ;
        RECT 15.750 58.765 15.920 58.935 ;
        RECT 15.420 58.595 15.920 58.765 ;
        RECT 6.985 57.205 12.330 57.640 ;
        RECT 12.505 57.205 13.715 58.295 ;
        RECT 14.035 57.205 14.365 58.355 ;
        RECT 14.535 58.225 15.545 58.395 ;
        RECT 14.535 57.375 14.705 58.225 ;
        RECT 14.875 57.205 15.205 58.005 ;
        RECT 15.375 57.375 15.545 58.225 ;
        RECT 15.750 58.355 15.920 58.595 ;
        RECT 16.090 58.525 16.470 58.765 ;
        RECT 18.230 58.380 18.570 59.210 ;
        RECT 22.165 58.985 25.675 59.755 ;
        RECT 26.310 59.015 26.565 59.585 ;
        RECT 26.735 59.355 27.065 59.755 ;
        RECT 27.490 59.220 28.020 59.585 ;
        RECT 28.210 59.415 28.485 59.585 ;
        RECT 28.205 59.245 28.485 59.415 ;
        RECT 27.490 59.185 27.665 59.220 ;
        RECT 26.735 59.015 27.665 59.185 ;
        RECT 15.750 58.185 16.465 58.355 ;
        RECT 15.725 57.205 15.965 58.005 ;
        RECT 16.135 57.375 16.465 58.185 ;
        RECT 20.050 57.640 20.400 58.890 ;
        RECT 22.165 58.465 23.815 58.985 ;
        RECT 23.985 58.295 25.675 58.815 ;
        RECT 16.645 57.205 21.990 57.640 ;
        RECT 22.165 57.205 25.675 58.295 ;
        RECT 26.310 58.345 26.480 59.015 ;
        RECT 26.735 58.845 26.905 59.015 ;
        RECT 26.650 58.515 26.905 58.845 ;
        RECT 27.130 58.515 27.325 58.845 ;
        RECT 26.310 57.375 26.645 58.345 ;
        RECT 26.815 57.205 26.985 58.345 ;
        RECT 27.155 57.545 27.325 58.515 ;
        RECT 27.495 57.885 27.665 59.015 ;
        RECT 27.835 58.225 28.005 59.025 ;
        RECT 28.210 58.425 28.485 59.245 ;
        RECT 28.655 58.225 28.845 59.585 ;
        RECT 29.025 59.220 29.535 59.755 ;
        RECT 29.755 58.945 30.000 59.550 ;
        RECT 31.365 59.030 31.655 59.755 ;
        RECT 31.825 58.985 34.415 59.755 ;
        RECT 34.590 59.015 34.845 59.585 ;
        RECT 35.015 59.355 35.345 59.755 ;
        RECT 35.770 59.220 36.300 59.585 ;
        RECT 36.490 59.415 36.765 59.585 ;
        RECT 36.485 59.245 36.765 59.415 ;
        RECT 35.770 59.185 35.945 59.220 ;
        RECT 35.015 59.015 35.945 59.185 ;
        RECT 29.045 58.775 30.275 58.945 ;
        RECT 27.835 58.055 28.845 58.225 ;
        RECT 29.015 58.210 29.765 58.400 ;
        RECT 27.495 57.715 28.620 57.885 ;
        RECT 29.015 57.545 29.185 58.210 ;
        RECT 29.935 57.965 30.275 58.775 ;
        RECT 31.825 58.465 33.035 58.985 ;
        RECT 27.155 57.375 29.185 57.545 ;
        RECT 29.355 57.205 29.525 57.965 ;
        RECT 29.760 57.555 30.275 57.965 ;
        RECT 31.365 57.205 31.655 58.370 ;
        RECT 33.205 58.295 34.415 58.815 ;
        RECT 31.825 57.205 34.415 58.295 ;
        RECT 34.590 58.345 34.760 59.015 ;
        RECT 35.015 58.845 35.185 59.015 ;
        RECT 34.930 58.515 35.185 58.845 ;
        RECT 35.410 58.515 35.605 58.845 ;
        RECT 34.590 57.375 34.925 58.345 ;
        RECT 35.095 57.205 35.265 58.345 ;
        RECT 35.435 57.545 35.605 58.515 ;
        RECT 35.775 57.885 35.945 59.015 ;
        RECT 36.115 58.225 36.285 59.025 ;
        RECT 36.490 58.425 36.765 59.245 ;
        RECT 36.935 58.225 37.125 59.585 ;
        RECT 37.305 59.220 37.815 59.755 ;
        RECT 38.035 58.945 38.280 59.550 ;
        RECT 38.725 58.985 42.235 59.755 ;
        RECT 42.495 59.205 42.665 59.585 ;
        RECT 42.845 59.375 43.175 59.755 ;
        RECT 42.495 59.035 43.160 59.205 ;
        RECT 43.355 59.080 43.615 59.585 ;
        RECT 37.325 58.775 38.555 58.945 ;
        RECT 36.115 58.055 37.125 58.225 ;
        RECT 37.295 58.210 38.045 58.400 ;
        RECT 35.775 57.715 36.900 57.885 ;
        RECT 37.295 57.545 37.465 58.210 ;
        RECT 38.215 57.965 38.555 58.775 ;
        RECT 38.725 58.465 40.375 58.985 ;
        RECT 40.545 58.295 42.235 58.815 ;
        RECT 42.425 58.485 42.755 58.855 ;
        RECT 42.990 58.780 43.160 59.035 ;
        RECT 42.990 58.450 43.275 58.780 ;
        RECT 42.990 58.305 43.160 58.450 ;
        RECT 35.435 57.375 37.465 57.545 ;
        RECT 37.635 57.205 37.805 57.965 ;
        RECT 38.040 57.555 38.555 57.965 ;
        RECT 38.725 57.205 42.235 58.295 ;
        RECT 42.495 58.135 43.160 58.305 ;
        RECT 43.445 58.280 43.615 59.080 ;
        RECT 43.825 58.935 44.055 59.755 ;
        RECT 44.225 58.955 44.555 59.585 ;
        RECT 43.805 58.515 44.135 58.765 ;
        RECT 44.305 58.355 44.555 58.955 ;
        RECT 44.725 58.935 44.935 59.755 ;
        RECT 45.170 59.015 45.425 59.585 ;
        RECT 45.595 59.355 45.925 59.755 ;
        RECT 46.350 59.220 46.880 59.585 ;
        RECT 46.350 59.185 46.525 59.220 ;
        RECT 45.595 59.015 46.525 59.185 ;
        RECT 42.495 57.375 42.665 58.135 ;
        RECT 42.845 57.205 43.175 57.965 ;
        RECT 43.345 57.375 43.615 58.280 ;
        RECT 43.825 57.205 44.055 58.345 ;
        RECT 44.225 57.375 44.555 58.355 ;
        RECT 45.170 58.345 45.340 59.015 ;
        RECT 45.595 58.845 45.765 59.015 ;
        RECT 45.510 58.515 45.765 58.845 ;
        RECT 45.990 58.515 46.185 58.845 ;
        RECT 44.725 57.205 44.935 58.345 ;
        RECT 45.170 57.375 45.505 58.345 ;
        RECT 45.675 57.205 45.845 58.345 ;
        RECT 46.015 57.545 46.185 58.515 ;
        RECT 46.355 57.885 46.525 59.015 ;
        RECT 46.695 58.225 46.865 59.025 ;
        RECT 47.070 58.735 47.345 59.585 ;
        RECT 47.065 58.565 47.345 58.735 ;
        RECT 47.070 58.425 47.345 58.565 ;
        RECT 47.515 58.225 47.705 59.585 ;
        RECT 47.885 59.220 48.395 59.755 ;
        RECT 48.615 58.945 48.860 59.550 ;
        RECT 49.765 58.955 50.105 59.585 ;
        RECT 50.275 58.955 50.525 59.755 ;
        RECT 50.715 59.105 51.045 59.585 ;
        RECT 51.215 59.295 51.440 59.755 ;
        RECT 51.610 59.105 51.940 59.585 ;
        RECT 47.905 58.775 49.135 58.945 ;
        RECT 46.695 58.055 47.705 58.225 ;
        RECT 47.875 58.210 48.625 58.400 ;
        RECT 46.355 57.715 47.480 57.885 ;
        RECT 47.875 57.545 48.045 58.210 ;
        RECT 48.795 57.965 49.135 58.775 ;
        RECT 46.015 57.375 48.045 57.545 ;
        RECT 48.215 57.205 48.385 57.965 ;
        RECT 48.620 57.555 49.135 57.965 ;
        RECT 49.765 58.345 49.940 58.955 ;
        RECT 50.715 58.935 51.940 59.105 ;
        RECT 52.570 58.975 53.070 59.585 ;
        RECT 53.445 58.985 56.955 59.755 ;
        RECT 57.125 59.030 57.415 59.755 ;
        RECT 50.110 58.595 50.805 58.765 ;
        RECT 50.635 58.345 50.805 58.595 ;
        RECT 50.980 58.565 51.400 58.765 ;
        RECT 51.570 58.565 51.900 58.765 ;
        RECT 52.070 58.565 52.400 58.765 ;
        RECT 52.570 58.345 52.740 58.975 ;
        RECT 52.925 58.515 53.275 58.765 ;
        RECT 53.445 58.465 55.095 58.985 ;
        RECT 58.510 58.915 58.770 59.755 ;
        RECT 58.945 59.010 59.200 59.585 ;
        RECT 59.370 59.375 59.700 59.755 ;
        RECT 59.915 59.205 60.085 59.585 ;
        RECT 59.370 59.035 60.085 59.205 ;
        RECT 60.350 59.205 60.605 59.495 ;
        RECT 60.775 59.375 61.105 59.755 ;
        RECT 60.350 59.035 61.100 59.205 ;
        RECT 49.765 57.375 50.105 58.345 ;
        RECT 50.275 57.205 50.445 58.345 ;
        RECT 50.635 58.175 53.070 58.345 ;
        RECT 55.265 58.295 56.955 58.815 ;
        RECT 50.715 57.205 50.965 58.005 ;
        RECT 51.610 57.375 51.940 58.175 ;
        RECT 52.240 57.205 52.570 58.005 ;
        RECT 52.740 57.375 53.070 58.175 ;
        RECT 53.445 57.205 56.955 58.295 ;
        RECT 57.125 57.205 57.415 58.370 ;
        RECT 58.510 57.205 58.770 58.355 ;
        RECT 58.945 58.280 59.115 59.010 ;
        RECT 59.370 58.845 59.540 59.035 ;
        RECT 59.285 58.515 59.540 58.845 ;
        RECT 59.370 58.305 59.540 58.515 ;
        RECT 59.820 58.485 60.175 58.855 ;
        RECT 58.945 57.375 59.200 58.280 ;
        RECT 59.370 58.135 60.085 58.305 ;
        RECT 60.350 58.215 60.700 58.865 ;
        RECT 59.370 57.205 59.700 57.965 ;
        RECT 59.915 57.375 60.085 58.135 ;
        RECT 60.870 58.045 61.100 59.035 ;
        RECT 60.350 57.875 61.100 58.045 ;
        RECT 60.350 57.375 60.605 57.875 ;
        RECT 60.775 57.205 61.105 57.705 ;
        RECT 61.275 57.375 61.445 59.495 ;
        RECT 61.805 59.395 62.135 59.755 ;
        RECT 62.305 59.365 62.800 59.535 ;
        RECT 63.005 59.365 63.860 59.535 ;
        RECT 61.675 58.175 62.135 59.225 ;
        RECT 61.615 57.390 61.940 58.175 ;
        RECT 62.305 58.005 62.475 59.365 ;
        RECT 62.645 58.455 62.995 59.075 ;
        RECT 63.165 58.855 63.520 59.075 ;
        RECT 63.165 58.265 63.335 58.855 ;
        RECT 63.690 58.655 63.860 59.365 ;
        RECT 64.735 59.295 65.065 59.755 ;
        RECT 65.275 59.395 65.625 59.565 ;
        RECT 64.065 58.825 64.855 59.075 ;
        RECT 65.275 59.005 65.535 59.395 ;
        RECT 65.845 59.305 66.795 59.585 ;
        RECT 66.965 59.315 67.155 59.755 ;
        RECT 67.325 59.375 68.395 59.545 ;
        RECT 65.025 58.655 65.195 58.835 ;
        RECT 62.305 57.835 62.700 58.005 ;
        RECT 62.870 57.875 63.335 58.265 ;
        RECT 63.505 58.485 65.195 58.655 ;
        RECT 62.530 57.705 62.700 57.835 ;
        RECT 63.505 57.705 63.675 58.485 ;
        RECT 65.365 58.315 65.535 59.005 ;
        RECT 64.035 58.145 65.535 58.315 ;
        RECT 65.725 58.345 65.935 59.135 ;
        RECT 66.105 58.515 66.455 59.135 ;
        RECT 66.625 58.525 66.795 59.305 ;
        RECT 67.325 59.145 67.495 59.375 ;
        RECT 66.965 58.975 67.495 59.145 ;
        RECT 66.965 58.695 67.185 58.975 ;
        RECT 67.665 58.805 67.905 59.205 ;
        RECT 66.625 58.355 67.030 58.525 ;
        RECT 67.365 58.435 67.905 58.805 ;
        RECT 68.075 59.020 68.395 59.375 ;
        RECT 68.640 59.295 68.945 59.755 ;
        RECT 69.115 59.045 69.370 59.575 ;
        RECT 68.075 58.845 68.400 59.020 ;
        RECT 68.075 58.545 68.990 58.845 ;
        RECT 68.250 58.515 68.990 58.545 ;
        RECT 65.725 58.185 66.400 58.345 ;
        RECT 66.860 58.265 67.030 58.355 ;
        RECT 65.725 58.175 66.690 58.185 ;
        RECT 65.365 58.005 65.535 58.145 ;
        RECT 62.110 57.205 62.360 57.665 ;
        RECT 62.530 57.375 62.780 57.705 ;
        RECT 62.995 57.375 63.675 57.705 ;
        RECT 63.845 57.805 64.920 57.975 ;
        RECT 65.365 57.835 65.925 58.005 ;
        RECT 66.230 57.885 66.690 58.175 ;
        RECT 66.860 58.095 68.080 58.265 ;
        RECT 63.845 57.465 64.015 57.805 ;
        RECT 64.250 57.205 64.580 57.635 ;
        RECT 64.750 57.465 64.920 57.805 ;
        RECT 65.215 57.205 65.585 57.665 ;
        RECT 65.755 57.375 65.925 57.835 ;
        RECT 66.860 57.715 67.030 58.095 ;
        RECT 68.250 57.925 68.420 58.515 ;
        RECT 69.160 58.395 69.370 59.045 ;
        RECT 66.160 57.375 67.030 57.715 ;
        RECT 67.620 57.755 68.420 57.925 ;
        RECT 67.200 57.205 67.450 57.665 ;
        RECT 67.620 57.465 67.790 57.755 ;
        RECT 67.970 57.205 68.300 57.585 ;
        RECT 68.640 57.205 68.945 58.345 ;
        RECT 69.115 57.515 69.370 58.395 ;
        RECT 69.550 59.015 69.805 59.585 ;
        RECT 69.975 59.355 70.305 59.755 ;
        RECT 70.730 59.220 71.260 59.585 ;
        RECT 71.450 59.415 71.725 59.585 ;
        RECT 71.445 59.245 71.725 59.415 ;
        RECT 70.730 59.185 70.905 59.220 ;
        RECT 69.975 59.015 70.905 59.185 ;
        RECT 69.550 58.345 69.720 59.015 ;
        RECT 69.975 58.845 70.145 59.015 ;
        RECT 69.890 58.515 70.145 58.845 ;
        RECT 70.370 58.515 70.565 58.845 ;
        RECT 69.550 57.375 69.885 58.345 ;
        RECT 70.055 57.205 70.225 58.345 ;
        RECT 70.395 57.545 70.565 58.515 ;
        RECT 70.735 57.885 70.905 59.015 ;
        RECT 71.075 58.225 71.245 59.025 ;
        RECT 71.450 58.425 71.725 59.245 ;
        RECT 71.895 58.225 72.085 59.585 ;
        RECT 72.265 59.220 72.775 59.755 ;
        RECT 72.995 58.945 73.240 59.550 ;
        RECT 74.420 58.945 74.665 59.550 ;
        RECT 74.885 59.220 75.395 59.755 ;
        RECT 72.285 58.775 73.515 58.945 ;
        RECT 71.075 58.055 72.085 58.225 ;
        RECT 72.255 58.210 73.005 58.400 ;
        RECT 70.735 57.715 71.860 57.885 ;
        RECT 72.255 57.545 72.425 58.210 ;
        RECT 73.175 57.965 73.515 58.775 ;
        RECT 70.395 57.375 72.425 57.545 ;
        RECT 72.595 57.205 72.765 57.965 ;
        RECT 73.000 57.555 73.515 57.965 ;
        RECT 74.145 58.775 75.375 58.945 ;
        RECT 74.145 57.965 74.485 58.775 ;
        RECT 74.655 58.210 75.405 58.400 ;
        RECT 74.145 57.555 74.660 57.965 ;
        RECT 74.895 57.205 75.065 57.965 ;
        RECT 75.235 57.545 75.405 58.210 ;
        RECT 75.575 58.225 75.765 59.585 ;
        RECT 75.935 58.735 76.210 59.585 ;
        RECT 76.400 59.220 76.930 59.585 ;
        RECT 77.355 59.355 77.685 59.755 ;
        RECT 76.755 59.185 76.930 59.220 ;
        RECT 75.935 58.565 76.215 58.735 ;
        RECT 75.935 58.425 76.210 58.565 ;
        RECT 76.415 58.225 76.585 59.025 ;
        RECT 75.575 58.055 76.585 58.225 ;
        RECT 76.755 59.015 77.685 59.185 ;
        RECT 77.855 59.015 78.110 59.585 ;
        RECT 76.755 57.885 76.925 59.015 ;
        RECT 77.515 58.845 77.685 59.015 ;
        RECT 75.800 57.715 76.925 57.885 ;
        RECT 77.095 58.515 77.290 58.845 ;
        RECT 77.515 58.515 77.770 58.845 ;
        RECT 77.095 57.545 77.265 58.515 ;
        RECT 77.940 58.345 78.110 59.015 ;
        RECT 78.285 58.985 81.795 59.755 ;
        RECT 82.885 59.030 83.175 59.755 ;
        RECT 78.285 58.465 79.935 58.985 ;
        RECT 83.550 58.975 84.050 59.585 ;
        RECT 75.235 57.375 77.265 57.545 ;
        RECT 77.435 57.205 77.605 58.345 ;
        RECT 77.775 57.375 78.110 58.345 ;
        RECT 80.105 58.295 81.795 58.815 ;
        RECT 83.345 58.515 83.695 58.765 ;
        RECT 78.285 57.205 81.795 58.295 ;
        RECT 82.885 57.205 83.175 58.370 ;
        RECT 83.880 58.345 84.050 58.975 ;
        RECT 84.680 59.105 85.010 59.585 ;
        RECT 85.180 59.295 85.405 59.755 ;
        RECT 85.575 59.105 85.905 59.585 ;
        RECT 84.680 58.935 85.905 59.105 ;
        RECT 86.095 58.955 86.345 59.755 ;
        RECT 86.515 58.955 86.855 59.585 ;
        RECT 87.025 59.210 92.370 59.755 ;
        RECT 92.545 59.210 97.890 59.755 ;
        RECT 84.220 58.565 84.550 58.765 ;
        RECT 84.720 58.565 85.050 58.765 ;
        RECT 85.220 58.565 85.640 58.765 ;
        RECT 85.815 58.595 86.510 58.765 ;
        RECT 85.815 58.345 85.985 58.595 ;
        RECT 86.680 58.345 86.855 58.955 ;
        RECT 88.610 58.380 88.950 59.210 ;
        RECT 83.550 58.175 85.985 58.345 ;
        RECT 83.550 57.375 83.880 58.175 ;
        RECT 84.050 57.205 84.380 58.005 ;
        RECT 84.680 57.375 85.010 58.175 ;
        RECT 85.655 57.205 85.905 58.005 ;
        RECT 86.175 57.205 86.345 58.345 ;
        RECT 86.515 57.375 86.855 58.345 ;
        RECT 90.430 57.640 90.780 58.890 ;
        RECT 94.130 58.380 94.470 59.210 ;
        RECT 98.065 58.985 100.655 59.755 ;
        RECT 100.830 59.015 101.085 59.585 ;
        RECT 101.255 59.355 101.585 59.755 ;
        RECT 102.010 59.220 102.540 59.585 ;
        RECT 102.730 59.415 103.005 59.585 ;
        RECT 102.725 59.245 103.005 59.415 ;
        RECT 102.010 59.185 102.185 59.220 ;
        RECT 101.255 59.015 102.185 59.185 ;
        RECT 95.950 57.640 96.300 58.890 ;
        RECT 98.065 58.465 99.275 58.985 ;
        RECT 99.445 58.295 100.655 58.815 ;
        RECT 87.025 57.205 92.370 57.640 ;
        RECT 92.545 57.205 97.890 57.640 ;
        RECT 98.065 57.205 100.655 58.295 ;
        RECT 100.830 58.345 101.000 59.015 ;
        RECT 101.255 58.845 101.425 59.015 ;
        RECT 101.170 58.515 101.425 58.845 ;
        RECT 101.650 58.515 101.845 58.845 ;
        RECT 100.830 57.375 101.165 58.345 ;
        RECT 101.335 57.205 101.505 58.345 ;
        RECT 101.675 57.545 101.845 58.515 ;
        RECT 102.015 57.885 102.185 59.015 ;
        RECT 102.355 58.225 102.525 59.025 ;
        RECT 102.730 58.425 103.005 59.245 ;
        RECT 103.175 58.225 103.365 59.585 ;
        RECT 103.545 59.220 104.055 59.755 ;
        RECT 104.275 58.945 104.520 59.550 ;
        RECT 103.565 58.775 104.795 58.945 ;
        RECT 105.025 58.935 105.235 59.755 ;
        RECT 105.405 58.955 105.735 59.585 ;
        RECT 102.355 58.055 103.365 58.225 ;
        RECT 103.535 58.210 104.285 58.400 ;
        RECT 102.015 57.715 103.140 57.885 ;
        RECT 103.535 57.545 103.705 58.210 ;
        RECT 104.455 57.965 104.795 58.775 ;
        RECT 105.405 58.355 105.655 58.955 ;
        RECT 105.905 58.935 106.135 59.755 ;
        RECT 106.345 58.985 108.015 59.755 ;
        RECT 108.645 59.030 108.935 59.755 ;
        RECT 109.105 58.985 111.695 59.755 ;
        RECT 112.325 59.005 113.535 59.755 ;
        RECT 105.825 58.515 106.155 58.765 ;
        RECT 106.345 58.465 107.095 58.985 ;
        RECT 101.675 57.375 103.705 57.545 ;
        RECT 103.875 57.205 104.045 57.965 ;
        RECT 104.280 57.555 104.795 57.965 ;
        RECT 105.025 57.205 105.235 58.345 ;
        RECT 105.405 57.375 105.735 58.355 ;
        RECT 105.905 57.205 106.135 58.345 ;
        RECT 107.265 58.295 108.015 58.815 ;
        RECT 109.105 58.465 110.315 58.985 ;
        RECT 106.345 57.205 108.015 58.295 ;
        RECT 108.645 57.205 108.935 58.370 ;
        RECT 110.485 58.295 111.695 58.815 ;
        RECT 109.105 57.205 111.695 58.295 ;
        RECT 112.325 58.295 112.845 58.835 ;
        RECT 113.015 58.465 113.535 59.005 ;
        RECT 112.325 57.205 113.535 58.295 ;
        RECT 5.520 57.035 113.620 57.205 ;
        RECT 5.605 55.945 6.815 57.035 ;
        RECT 6.985 55.945 10.495 57.035 ;
        RECT 5.605 55.235 6.125 55.775 ;
        RECT 6.295 55.405 6.815 55.945 ;
        RECT 6.985 55.255 8.635 55.775 ;
        RECT 8.805 55.425 10.495 55.945 ;
        RECT 11.125 55.960 11.395 56.865 ;
        RECT 11.565 56.275 11.895 57.035 ;
        RECT 12.075 56.105 12.245 56.865 ;
        RECT 5.605 54.485 6.815 55.235 ;
        RECT 6.985 54.485 10.495 55.255 ;
        RECT 11.125 55.160 11.295 55.960 ;
        RECT 11.580 55.935 12.245 56.105 ;
        RECT 12.975 56.055 13.305 56.865 ;
        RECT 13.475 56.235 13.715 57.035 ;
        RECT 11.580 55.790 11.750 55.935 ;
        RECT 12.975 55.885 13.690 56.055 ;
        RECT 11.465 55.460 11.750 55.790 ;
        RECT 11.580 55.205 11.750 55.460 ;
        RECT 11.985 55.385 12.315 55.755 ;
        RECT 12.970 55.475 13.350 55.715 ;
        RECT 13.520 55.645 13.690 55.885 ;
        RECT 13.895 56.015 14.065 56.865 ;
        RECT 14.235 56.235 14.565 57.035 ;
        RECT 14.735 56.015 14.905 56.865 ;
        RECT 13.895 55.845 14.905 56.015 ;
        RECT 15.075 55.885 15.405 57.035 ;
        RECT 15.725 55.945 16.935 57.035 ;
        RECT 13.520 55.475 14.020 55.645 ;
        RECT 13.520 55.305 13.690 55.475 ;
        RECT 14.410 55.305 14.905 55.845 ;
        RECT 11.125 54.655 11.385 55.160 ;
        RECT 11.580 55.035 12.245 55.205 ;
        RECT 11.565 54.485 11.895 54.865 ;
        RECT 12.075 54.655 12.245 55.035 ;
        RECT 13.055 55.135 13.690 55.305 ;
        RECT 13.895 55.135 14.905 55.305 ;
        RECT 13.055 54.655 13.225 55.135 ;
        RECT 13.405 54.485 13.645 54.965 ;
        RECT 13.895 54.655 14.065 55.135 ;
        RECT 14.235 54.485 14.565 54.965 ;
        RECT 14.735 54.655 14.905 55.135 ;
        RECT 15.075 54.485 15.405 55.285 ;
        RECT 15.725 55.235 16.245 55.775 ;
        RECT 16.415 55.405 16.935 55.945 ;
        RECT 17.195 56.105 17.365 56.865 ;
        RECT 17.545 56.275 17.875 57.035 ;
        RECT 17.195 55.935 17.860 56.105 ;
        RECT 18.045 55.960 18.315 56.865 ;
        RECT 17.690 55.790 17.860 55.935 ;
        RECT 17.125 55.385 17.455 55.755 ;
        RECT 17.690 55.460 17.975 55.790 ;
        RECT 15.725 54.485 16.935 55.235 ;
        RECT 17.690 55.205 17.860 55.460 ;
        RECT 17.195 55.035 17.860 55.205 ;
        RECT 18.145 55.160 18.315 55.960 ;
        RECT 18.485 55.870 18.775 57.035 ;
        RECT 18.950 55.895 19.285 56.865 ;
        RECT 19.455 55.895 19.625 57.035 ;
        RECT 19.795 56.695 21.825 56.865 ;
        RECT 18.950 55.225 19.120 55.895 ;
        RECT 19.795 55.725 19.965 56.695 ;
        RECT 19.290 55.395 19.545 55.725 ;
        RECT 19.770 55.395 19.965 55.725 ;
        RECT 20.135 56.355 21.260 56.525 ;
        RECT 19.375 55.225 19.545 55.395 ;
        RECT 20.135 55.225 20.305 56.355 ;
        RECT 17.195 54.655 17.365 55.035 ;
        RECT 17.545 54.485 17.875 54.865 ;
        RECT 18.055 54.655 18.315 55.160 ;
        RECT 18.485 54.485 18.775 55.210 ;
        RECT 18.950 54.655 19.205 55.225 ;
        RECT 19.375 55.055 20.305 55.225 ;
        RECT 20.475 56.015 21.485 56.185 ;
        RECT 20.475 55.215 20.645 56.015 ;
        RECT 20.130 55.020 20.305 55.055 ;
        RECT 19.375 54.485 19.705 54.885 ;
        RECT 20.130 54.655 20.660 55.020 ;
        RECT 20.850 54.995 21.125 55.815 ;
        RECT 20.845 54.825 21.125 54.995 ;
        RECT 20.850 54.655 21.125 54.825 ;
        RECT 21.295 54.655 21.485 56.015 ;
        RECT 21.655 56.030 21.825 56.695 ;
        RECT 21.995 56.275 22.165 57.035 ;
        RECT 22.400 56.275 22.915 56.685 ;
        RECT 21.655 55.840 22.405 56.030 ;
        RECT 22.575 55.465 22.915 56.275 ;
        RECT 23.175 56.365 23.345 56.865 ;
        RECT 23.515 56.535 23.845 57.035 ;
        RECT 23.175 56.195 23.840 56.365 ;
        RECT 21.685 55.295 22.915 55.465 ;
        RECT 23.090 55.375 23.440 56.025 ;
        RECT 21.665 54.485 22.175 55.020 ;
        RECT 22.395 54.690 22.640 55.295 ;
        RECT 23.610 55.205 23.840 56.195 ;
        RECT 23.175 55.035 23.840 55.205 ;
        RECT 23.175 54.745 23.345 55.035 ;
        RECT 23.515 54.485 23.845 54.865 ;
        RECT 24.015 54.745 24.240 56.865 ;
        RECT 24.455 56.535 24.785 57.035 ;
        RECT 24.955 56.365 25.125 56.865 ;
        RECT 25.360 56.650 26.190 56.820 ;
        RECT 26.430 56.655 26.810 57.035 ;
        RECT 24.430 56.195 25.125 56.365 ;
        RECT 24.430 55.225 24.600 56.195 ;
        RECT 24.770 55.405 25.180 56.025 ;
        RECT 25.350 55.975 25.850 56.355 ;
        RECT 24.430 55.035 25.125 55.225 ;
        RECT 25.350 55.105 25.570 55.975 ;
        RECT 26.020 55.805 26.190 56.650 ;
        RECT 26.990 56.485 27.160 56.775 ;
        RECT 27.330 56.655 27.660 57.035 ;
        RECT 28.130 56.565 28.760 56.815 ;
        RECT 28.940 56.655 29.360 57.035 ;
        RECT 28.590 56.485 28.760 56.565 ;
        RECT 29.560 56.485 29.800 56.775 ;
        RECT 26.360 56.235 27.730 56.485 ;
        RECT 26.360 55.975 26.610 56.235 ;
        RECT 27.120 55.805 27.370 55.965 ;
        RECT 26.020 55.635 27.370 55.805 ;
        RECT 26.020 55.595 26.440 55.635 ;
        RECT 25.750 55.045 26.100 55.415 ;
        RECT 24.455 54.485 24.785 54.865 ;
        RECT 24.955 54.705 25.125 55.035 ;
        RECT 26.270 54.865 26.440 55.595 ;
        RECT 27.540 55.465 27.730 56.235 ;
        RECT 26.610 55.135 27.020 55.465 ;
        RECT 27.310 55.125 27.730 55.465 ;
        RECT 27.900 56.055 28.420 56.365 ;
        RECT 28.590 56.315 29.800 56.485 ;
        RECT 30.030 56.345 30.360 57.035 ;
        RECT 27.900 55.295 28.070 56.055 ;
        RECT 28.240 55.465 28.420 55.875 ;
        RECT 28.590 55.805 28.760 56.315 ;
        RECT 30.530 56.165 30.700 56.775 ;
        RECT 30.970 56.315 31.300 56.825 ;
        RECT 30.530 56.145 30.850 56.165 ;
        RECT 28.930 55.975 30.850 56.145 ;
        RECT 28.590 55.635 30.490 55.805 ;
        RECT 28.820 55.295 29.150 55.415 ;
        RECT 27.900 55.125 29.150 55.295 ;
        RECT 25.425 54.665 26.440 54.865 ;
        RECT 26.610 54.485 27.020 54.925 ;
        RECT 27.310 54.695 27.560 55.125 ;
        RECT 27.760 54.485 28.080 54.945 ;
        RECT 29.320 54.875 29.490 55.635 ;
        RECT 30.160 55.575 30.490 55.635 ;
        RECT 29.680 55.405 30.010 55.465 ;
        RECT 29.680 55.135 30.340 55.405 ;
        RECT 30.660 55.080 30.850 55.975 ;
        RECT 28.640 54.705 29.490 54.875 ;
        RECT 29.690 54.485 30.350 54.965 ;
        RECT 30.530 54.750 30.850 55.080 ;
        RECT 31.050 55.725 31.300 56.315 ;
        RECT 31.480 56.235 31.765 57.035 ;
        RECT 31.945 56.695 32.200 56.725 ;
        RECT 31.945 56.525 32.285 56.695 ;
        RECT 31.945 56.055 32.200 56.525 ;
        RECT 32.835 56.365 33.005 56.865 ;
        RECT 33.175 56.535 33.505 57.035 ;
        RECT 32.835 56.195 33.500 56.365 ;
        RECT 31.050 55.395 31.850 55.725 ;
        RECT 31.050 54.745 31.300 55.395 ;
        RECT 32.020 55.195 32.200 56.055 ;
        RECT 32.750 55.375 33.100 56.025 ;
        RECT 33.270 55.205 33.500 56.195 ;
        RECT 31.480 54.485 31.765 54.945 ;
        RECT 31.945 54.665 32.200 55.195 ;
        RECT 32.835 55.035 33.500 55.205 ;
        RECT 32.835 54.745 33.005 55.035 ;
        RECT 33.175 54.485 33.505 54.865 ;
        RECT 33.675 54.745 33.900 56.865 ;
        RECT 34.115 56.535 34.445 57.035 ;
        RECT 34.615 56.365 34.785 56.865 ;
        RECT 35.020 56.650 35.850 56.820 ;
        RECT 36.090 56.655 36.470 57.035 ;
        RECT 34.090 56.195 34.785 56.365 ;
        RECT 34.090 55.225 34.260 56.195 ;
        RECT 34.430 55.405 34.840 56.025 ;
        RECT 35.010 55.975 35.510 56.355 ;
        RECT 34.090 55.035 34.785 55.225 ;
        RECT 35.010 55.105 35.230 55.975 ;
        RECT 35.680 55.805 35.850 56.650 ;
        RECT 36.650 56.485 36.820 56.775 ;
        RECT 36.990 56.655 37.320 57.035 ;
        RECT 37.790 56.565 38.420 56.815 ;
        RECT 38.600 56.655 39.020 57.035 ;
        RECT 38.250 56.485 38.420 56.565 ;
        RECT 39.220 56.485 39.460 56.775 ;
        RECT 36.020 56.235 37.390 56.485 ;
        RECT 36.020 55.975 36.270 56.235 ;
        RECT 36.780 55.805 37.030 55.965 ;
        RECT 35.680 55.635 37.030 55.805 ;
        RECT 35.680 55.595 36.100 55.635 ;
        RECT 35.410 55.045 35.760 55.415 ;
        RECT 34.115 54.485 34.445 54.865 ;
        RECT 34.615 54.705 34.785 55.035 ;
        RECT 35.930 54.865 36.100 55.595 ;
        RECT 37.200 55.465 37.390 56.235 ;
        RECT 36.270 55.135 36.680 55.465 ;
        RECT 36.970 55.125 37.390 55.465 ;
        RECT 37.560 56.055 38.080 56.365 ;
        RECT 38.250 56.315 39.460 56.485 ;
        RECT 39.690 56.345 40.020 57.035 ;
        RECT 37.560 55.295 37.730 56.055 ;
        RECT 37.900 55.465 38.080 55.875 ;
        RECT 38.250 55.805 38.420 56.315 ;
        RECT 40.190 56.165 40.360 56.775 ;
        RECT 40.630 56.315 40.960 56.825 ;
        RECT 40.190 56.145 40.510 56.165 ;
        RECT 38.590 55.975 40.510 56.145 ;
        RECT 38.250 55.635 40.150 55.805 ;
        RECT 38.480 55.295 38.810 55.415 ;
        RECT 37.560 55.125 38.810 55.295 ;
        RECT 35.085 54.665 36.100 54.865 ;
        RECT 36.270 54.485 36.680 54.925 ;
        RECT 36.970 54.695 37.220 55.125 ;
        RECT 37.420 54.485 37.740 54.945 ;
        RECT 38.980 54.875 39.150 55.635 ;
        RECT 39.820 55.575 40.150 55.635 ;
        RECT 39.340 55.405 39.670 55.465 ;
        RECT 39.340 55.135 40.000 55.405 ;
        RECT 40.320 55.080 40.510 55.975 ;
        RECT 38.300 54.705 39.150 54.875 ;
        RECT 39.350 54.485 40.010 54.965 ;
        RECT 40.190 54.750 40.510 55.080 ;
        RECT 40.710 55.725 40.960 56.315 ;
        RECT 41.140 56.235 41.425 57.035 ;
        RECT 41.605 56.695 41.860 56.725 ;
        RECT 41.605 56.525 41.945 56.695 ;
        RECT 41.605 56.055 41.860 56.525 ;
        RECT 40.710 55.395 41.510 55.725 ;
        RECT 40.710 54.745 40.960 55.395 ;
        RECT 41.680 55.195 41.860 56.055 ;
        RECT 42.405 55.945 44.075 57.035 ;
        RECT 41.140 54.485 41.425 54.945 ;
        RECT 41.605 54.665 41.860 55.195 ;
        RECT 42.405 55.255 43.155 55.775 ;
        RECT 43.325 55.425 44.075 55.945 ;
        RECT 44.245 55.870 44.535 57.035 ;
        RECT 44.705 55.945 46.375 57.035 ;
        RECT 44.705 55.255 45.455 55.775 ;
        RECT 45.625 55.425 46.375 55.945 ;
        RECT 47.005 55.960 47.275 56.865 ;
        RECT 47.445 56.275 47.775 57.035 ;
        RECT 47.955 56.105 48.125 56.865 ;
        RECT 42.405 54.485 44.075 55.255 ;
        RECT 44.245 54.485 44.535 55.210 ;
        RECT 44.705 54.485 46.375 55.255 ;
        RECT 47.005 55.160 47.175 55.960 ;
        RECT 47.460 55.935 48.125 56.105 ;
        RECT 47.460 55.790 47.630 55.935 ;
        RECT 47.345 55.460 47.630 55.790 ;
        RECT 48.390 55.895 48.725 56.865 ;
        RECT 48.895 55.895 49.065 57.035 ;
        RECT 49.235 56.695 51.265 56.865 ;
        RECT 47.460 55.205 47.630 55.460 ;
        RECT 47.865 55.385 48.195 55.755 ;
        RECT 48.390 55.225 48.560 55.895 ;
        RECT 49.235 55.725 49.405 56.695 ;
        RECT 48.730 55.395 48.985 55.725 ;
        RECT 49.210 55.395 49.405 55.725 ;
        RECT 49.575 56.355 50.700 56.525 ;
        RECT 48.815 55.225 48.985 55.395 ;
        RECT 49.575 55.225 49.745 56.355 ;
        RECT 47.005 54.655 47.265 55.160 ;
        RECT 47.460 55.035 48.125 55.205 ;
        RECT 47.445 54.485 47.775 54.865 ;
        RECT 47.955 54.655 48.125 55.035 ;
        RECT 48.390 54.655 48.645 55.225 ;
        RECT 48.815 55.055 49.745 55.225 ;
        RECT 49.915 56.015 50.925 56.185 ;
        RECT 49.915 55.215 50.085 56.015 ;
        RECT 50.290 55.675 50.565 55.815 ;
        RECT 50.285 55.505 50.565 55.675 ;
        RECT 49.570 55.020 49.745 55.055 ;
        RECT 48.815 54.485 49.145 54.885 ;
        RECT 49.570 54.655 50.100 55.020 ;
        RECT 50.290 54.655 50.565 55.505 ;
        RECT 50.735 54.655 50.925 56.015 ;
        RECT 51.095 56.030 51.265 56.695 ;
        RECT 51.435 56.275 51.605 57.035 ;
        RECT 51.840 56.275 52.355 56.685 ;
        RECT 51.095 55.840 51.845 56.030 ;
        RECT 52.015 55.465 52.355 56.275 ;
        RECT 51.125 55.295 52.355 55.465 ;
        RECT 52.530 55.895 52.865 56.865 ;
        RECT 53.035 55.895 53.205 57.035 ;
        RECT 53.375 56.695 55.405 56.865 ;
        RECT 51.105 54.485 51.615 55.020 ;
        RECT 51.835 54.690 52.080 55.295 ;
        RECT 52.530 55.225 52.700 55.895 ;
        RECT 53.375 55.725 53.545 56.695 ;
        RECT 52.870 55.395 53.125 55.725 ;
        RECT 53.350 55.395 53.545 55.725 ;
        RECT 53.715 56.355 54.840 56.525 ;
        RECT 52.955 55.225 53.125 55.395 ;
        RECT 53.715 55.225 53.885 56.355 ;
        RECT 52.530 54.655 52.785 55.225 ;
        RECT 52.955 55.055 53.885 55.225 ;
        RECT 54.055 56.015 55.065 56.185 ;
        RECT 54.055 55.215 54.225 56.015 ;
        RECT 54.430 55.675 54.705 55.815 ;
        RECT 54.425 55.505 54.705 55.675 ;
        RECT 53.710 55.020 53.885 55.055 ;
        RECT 52.955 54.485 53.285 54.885 ;
        RECT 53.710 54.655 54.240 55.020 ;
        RECT 54.430 54.655 54.705 55.505 ;
        RECT 54.875 54.655 55.065 56.015 ;
        RECT 55.235 56.030 55.405 56.695 ;
        RECT 55.575 56.275 55.745 57.035 ;
        RECT 55.980 56.275 56.495 56.685 ;
        RECT 55.235 55.840 55.985 56.030 ;
        RECT 56.155 55.465 56.495 56.275 ;
        RECT 56.665 55.945 60.175 57.035 ;
        RECT 55.265 55.295 56.495 55.465 ;
        RECT 55.245 54.485 55.755 55.020 ;
        RECT 55.975 54.690 56.220 55.295 ;
        RECT 56.665 55.255 58.315 55.775 ;
        RECT 58.485 55.425 60.175 55.945 ;
        RECT 60.350 55.885 60.610 57.035 ;
        RECT 60.785 55.960 61.040 56.865 ;
        RECT 61.210 56.275 61.540 57.035 ;
        RECT 61.755 56.105 61.925 56.865 ;
        RECT 56.665 54.485 60.175 55.255 ;
        RECT 60.350 54.485 60.610 55.325 ;
        RECT 60.785 55.230 60.955 55.960 ;
        RECT 61.210 55.935 61.925 56.105 ;
        RECT 62.185 55.945 64.775 57.035 ;
        RECT 61.210 55.725 61.380 55.935 ;
        RECT 61.125 55.395 61.380 55.725 ;
        RECT 60.785 54.655 61.040 55.230 ;
        RECT 61.210 55.205 61.380 55.395 ;
        RECT 61.660 55.385 62.015 55.755 ;
        RECT 62.185 55.255 63.395 55.775 ;
        RECT 63.565 55.425 64.775 55.945 ;
        RECT 65.005 55.895 65.215 57.035 ;
        RECT 65.385 55.885 65.715 56.865 ;
        RECT 65.885 55.895 66.115 57.035 ;
        RECT 66.335 56.055 66.665 56.865 ;
        RECT 66.835 56.235 67.075 57.035 ;
        RECT 66.335 55.885 67.050 56.055 ;
        RECT 61.210 55.035 61.925 55.205 ;
        RECT 61.210 54.485 61.540 54.865 ;
        RECT 61.755 54.655 61.925 55.035 ;
        RECT 62.185 54.485 64.775 55.255 ;
        RECT 65.005 54.485 65.215 55.305 ;
        RECT 65.385 55.285 65.635 55.885 ;
        RECT 65.805 55.475 66.135 55.725 ;
        RECT 66.330 55.475 66.710 55.715 ;
        RECT 66.880 55.645 67.050 55.885 ;
        RECT 67.255 56.015 67.425 56.865 ;
        RECT 67.595 56.235 67.925 57.035 ;
        RECT 68.095 56.015 68.265 56.865 ;
        RECT 67.255 55.845 68.265 56.015 ;
        RECT 68.435 55.885 68.765 57.035 ;
        RECT 70.005 55.870 70.295 57.035 ;
        RECT 70.470 56.365 70.725 56.865 ;
        RECT 70.895 56.535 71.225 57.035 ;
        RECT 70.470 56.195 71.220 56.365 ;
        RECT 66.880 55.475 67.380 55.645 ;
        RECT 66.880 55.305 67.050 55.475 ;
        RECT 67.770 55.305 68.265 55.845 ;
        RECT 70.470 55.375 70.820 56.025 ;
        RECT 65.385 54.655 65.715 55.285 ;
        RECT 65.885 54.485 66.115 55.305 ;
        RECT 66.415 55.135 67.050 55.305 ;
        RECT 67.255 55.135 68.265 55.305 ;
        RECT 66.415 54.655 66.585 55.135 ;
        RECT 66.765 54.485 67.005 54.965 ;
        RECT 67.255 54.655 67.425 55.135 ;
        RECT 67.595 54.485 67.925 54.965 ;
        RECT 68.095 54.655 68.265 55.135 ;
        RECT 68.435 54.485 68.765 55.285 ;
        RECT 70.005 54.485 70.295 55.210 ;
        RECT 70.990 55.205 71.220 56.195 ;
        RECT 70.470 55.035 71.220 55.205 ;
        RECT 70.470 54.745 70.725 55.035 ;
        RECT 70.895 54.485 71.225 54.865 ;
        RECT 71.395 54.745 71.565 56.865 ;
        RECT 71.735 56.065 72.060 56.850 ;
        RECT 72.230 56.575 72.480 57.035 ;
        RECT 72.650 56.535 72.900 56.865 ;
        RECT 73.115 56.535 73.795 56.865 ;
        RECT 72.650 56.405 72.820 56.535 ;
        RECT 72.425 56.235 72.820 56.405 ;
        RECT 71.795 55.015 72.255 56.065 ;
        RECT 72.425 54.875 72.595 56.235 ;
        RECT 72.990 55.975 73.455 56.365 ;
        RECT 72.765 55.165 73.115 55.785 ;
        RECT 73.285 55.385 73.455 55.975 ;
        RECT 73.625 55.755 73.795 56.535 ;
        RECT 73.965 56.435 74.135 56.775 ;
        RECT 74.370 56.605 74.700 57.035 ;
        RECT 74.870 56.435 75.040 56.775 ;
        RECT 75.335 56.575 75.705 57.035 ;
        RECT 73.965 56.265 75.040 56.435 ;
        RECT 75.875 56.405 76.045 56.865 ;
        RECT 76.280 56.525 77.150 56.865 ;
        RECT 77.320 56.575 77.570 57.035 ;
        RECT 75.485 56.235 76.045 56.405 ;
        RECT 75.485 56.095 75.655 56.235 ;
        RECT 74.155 55.925 75.655 56.095 ;
        RECT 76.350 56.065 76.810 56.355 ;
        RECT 73.625 55.585 75.315 55.755 ;
        RECT 73.285 55.165 73.640 55.385 ;
        RECT 73.810 54.875 73.980 55.585 ;
        RECT 74.185 55.165 74.975 55.415 ;
        RECT 75.145 55.405 75.315 55.585 ;
        RECT 75.485 55.235 75.655 55.925 ;
        RECT 71.925 54.485 72.255 54.845 ;
        RECT 72.425 54.705 72.920 54.875 ;
        RECT 73.125 54.705 73.980 54.875 ;
        RECT 74.855 54.485 75.185 54.945 ;
        RECT 75.395 54.845 75.655 55.235 ;
        RECT 75.845 56.055 76.810 56.065 ;
        RECT 76.980 56.145 77.150 56.525 ;
        RECT 77.740 56.485 77.910 56.775 ;
        RECT 78.090 56.655 78.420 57.035 ;
        RECT 77.740 56.315 78.540 56.485 ;
        RECT 75.845 55.895 76.520 56.055 ;
        RECT 76.980 55.975 78.200 56.145 ;
        RECT 75.845 55.105 76.055 55.895 ;
        RECT 76.980 55.885 77.150 55.975 ;
        RECT 76.225 55.105 76.575 55.725 ;
        RECT 76.745 55.715 77.150 55.885 ;
        RECT 76.745 54.935 76.915 55.715 ;
        RECT 77.085 55.265 77.305 55.545 ;
        RECT 77.485 55.435 78.025 55.805 ;
        RECT 78.370 55.725 78.540 56.315 ;
        RECT 78.760 55.895 79.065 57.035 ;
        RECT 79.235 55.845 79.490 56.725 ;
        RECT 78.370 55.695 79.110 55.725 ;
        RECT 77.085 55.095 77.615 55.265 ;
        RECT 75.395 54.675 75.745 54.845 ;
        RECT 75.965 54.655 76.915 54.935 ;
        RECT 77.085 54.485 77.275 54.925 ;
        RECT 77.445 54.865 77.615 55.095 ;
        RECT 77.785 55.035 78.025 55.435 ;
        RECT 78.195 55.395 79.110 55.695 ;
        RECT 78.195 55.220 78.520 55.395 ;
        RECT 78.195 54.865 78.515 55.220 ;
        RECT 79.280 55.195 79.490 55.845 ;
        RECT 77.445 54.695 78.515 54.865 ;
        RECT 78.760 54.485 79.065 54.945 ;
        RECT 79.235 54.665 79.490 55.195 ;
        RECT 79.665 55.960 79.935 56.865 ;
        RECT 80.105 56.275 80.435 57.035 ;
        RECT 80.615 56.105 80.785 56.865 ;
        RECT 79.665 55.160 79.835 55.960 ;
        RECT 80.120 55.935 80.785 56.105 ;
        RECT 81.045 56.275 81.560 56.685 ;
        RECT 81.795 56.275 81.965 57.035 ;
        RECT 82.135 56.695 84.165 56.865 ;
        RECT 80.120 55.790 80.290 55.935 ;
        RECT 80.005 55.460 80.290 55.790 ;
        RECT 80.120 55.205 80.290 55.460 ;
        RECT 80.525 55.385 80.855 55.755 ;
        RECT 81.045 55.465 81.385 56.275 ;
        RECT 82.135 56.030 82.305 56.695 ;
        RECT 82.700 56.355 83.825 56.525 ;
        RECT 81.555 55.840 82.305 56.030 ;
        RECT 82.475 56.015 83.485 56.185 ;
        RECT 81.045 55.295 82.275 55.465 ;
        RECT 79.665 54.655 79.925 55.160 ;
        RECT 80.120 55.035 80.785 55.205 ;
        RECT 80.105 54.485 80.435 54.865 ;
        RECT 80.615 54.655 80.785 55.035 ;
        RECT 81.320 54.690 81.565 55.295 ;
        RECT 81.785 54.485 82.295 55.020 ;
        RECT 82.475 54.655 82.665 56.015 ;
        RECT 82.835 55.335 83.110 55.815 ;
        RECT 82.835 55.165 83.115 55.335 ;
        RECT 83.315 55.215 83.485 56.015 ;
        RECT 83.655 55.225 83.825 56.355 ;
        RECT 83.995 55.725 84.165 56.695 ;
        RECT 84.335 55.895 84.505 57.035 ;
        RECT 84.675 55.895 85.010 56.865 ;
        RECT 83.995 55.395 84.190 55.725 ;
        RECT 84.415 55.395 84.670 55.725 ;
        RECT 84.415 55.225 84.585 55.395 ;
        RECT 84.840 55.225 85.010 55.895 ;
        RECT 82.835 54.655 83.110 55.165 ;
        RECT 83.655 55.055 84.585 55.225 ;
        RECT 83.655 55.020 83.830 55.055 ;
        RECT 83.300 54.655 83.830 55.020 ;
        RECT 84.255 54.485 84.585 54.885 ;
        RECT 84.755 54.655 85.010 55.225 ;
        RECT 85.185 55.960 85.455 56.865 ;
        RECT 85.625 56.275 85.955 57.035 ;
        RECT 86.135 56.105 86.305 56.865 ;
        RECT 85.185 55.160 85.355 55.960 ;
        RECT 85.640 55.935 86.305 56.105 ;
        RECT 86.565 55.945 87.775 57.035 ;
        RECT 85.640 55.790 85.810 55.935 ;
        RECT 85.525 55.460 85.810 55.790 ;
        RECT 85.640 55.205 85.810 55.460 ;
        RECT 86.045 55.385 86.375 55.755 ;
        RECT 86.565 55.235 87.085 55.775 ;
        RECT 87.255 55.405 87.775 55.945 ;
        RECT 87.945 55.960 88.215 56.865 ;
        RECT 88.385 56.275 88.715 57.035 ;
        RECT 88.895 56.105 89.065 56.865 ;
        RECT 85.185 54.655 85.445 55.160 ;
        RECT 85.640 55.035 86.305 55.205 ;
        RECT 85.625 54.485 85.955 54.865 ;
        RECT 86.135 54.655 86.305 55.035 ;
        RECT 86.565 54.485 87.775 55.235 ;
        RECT 87.945 55.160 88.115 55.960 ;
        RECT 88.400 55.935 89.065 56.105 ;
        RECT 88.400 55.790 88.570 55.935 ;
        RECT 88.285 55.460 88.570 55.790 ;
        RECT 89.330 55.895 89.665 56.865 ;
        RECT 89.835 55.895 90.005 57.035 ;
        RECT 90.175 56.695 92.205 56.865 ;
        RECT 88.400 55.205 88.570 55.460 ;
        RECT 88.805 55.385 89.135 55.755 ;
        RECT 89.330 55.225 89.500 55.895 ;
        RECT 90.175 55.725 90.345 56.695 ;
        RECT 89.670 55.395 89.925 55.725 ;
        RECT 90.150 55.395 90.345 55.725 ;
        RECT 90.515 56.355 91.640 56.525 ;
        RECT 89.755 55.225 89.925 55.395 ;
        RECT 90.515 55.225 90.685 56.355 ;
        RECT 87.945 54.655 88.205 55.160 ;
        RECT 88.400 55.035 89.065 55.205 ;
        RECT 88.385 54.485 88.715 54.865 ;
        RECT 88.895 54.655 89.065 55.035 ;
        RECT 89.330 54.655 89.585 55.225 ;
        RECT 89.755 55.055 90.685 55.225 ;
        RECT 90.855 56.015 91.865 56.185 ;
        RECT 90.855 55.215 91.025 56.015 ;
        RECT 90.510 55.020 90.685 55.055 ;
        RECT 89.755 54.485 90.085 54.885 ;
        RECT 90.510 54.655 91.040 55.020 ;
        RECT 91.230 54.995 91.505 55.815 ;
        RECT 91.225 54.825 91.505 54.995 ;
        RECT 91.230 54.655 91.505 54.825 ;
        RECT 91.675 54.655 91.865 56.015 ;
        RECT 92.035 56.030 92.205 56.695 ;
        RECT 92.375 56.275 92.545 57.035 ;
        RECT 92.780 56.275 93.295 56.685 ;
        RECT 92.035 55.840 92.785 56.030 ;
        RECT 92.955 55.465 93.295 56.275 ;
        RECT 93.465 55.945 95.135 57.035 ;
        RECT 92.065 55.295 93.295 55.465 ;
        RECT 92.045 54.485 92.555 55.020 ;
        RECT 92.775 54.690 93.020 55.295 ;
        RECT 93.465 55.255 94.215 55.775 ;
        RECT 94.385 55.425 95.135 55.945 ;
        RECT 95.765 55.870 96.055 57.035 ;
        RECT 97.235 56.105 97.405 56.865 ;
        RECT 97.585 56.275 97.915 57.035 ;
        RECT 97.235 55.935 97.900 56.105 ;
        RECT 98.085 55.960 98.355 56.865 ;
        RECT 97.730 55.790 97.900 55.935 ;
        RECT 97.165 55.385 97.495 55.755 ;
        RECT 97.730 55.460 98.015 55.790 ;
        RECT 93.465 54.485 95.135 55.255 ;
        RECT 95.765 54.485 96.055 55.210 ;
        RECT 97.730 55.205 97.900 55.460 ;
        RECT 97.235 55.035 97.900 55.205 ;
        RECT 98.185 55.160 98.355 55.960 ;
        RECT 98.615 56.105 98.785 56.865 ;
        RECT 98.965 56.275 99.295 57.035 ;
        RECT 98.615 55.935 99.280 56.105 ;
        RECT 99.465 55.960 99.735 56.865 ;
        RECT 99.995 56.365 100.165 56.865 ;
        RECT 100.335 56.535 100.665 57.035 ;
        RECT 99.995 56.195 100.660 56.365 ;
        RECT 99.110 55.790 99.280 55.935 ;
        RECT 98.545 55.385 98.875 55.755 ;
        RECT 99.110 55.460 99.395 55.790 ;
        RECT 99.110 55.205 99.280 55.460 ;
        RECT 97.235 54.655 97.405 55.035 ;
        RECT 97.585 54.485 97.915 54.865 ;
        RECT 98.095 54.655 98.355 55.160 ;
        RECT 98.615 55.035 99.280 55.205 ;
        RECT 99.565 55.160 99.735 55.960 ;
        RECT 99.910 55.375 100.260 56.025 ;
        RECT 100.430 55.205 100.660 56.195 ;
        RECT 98.615 54.655 98.785 55.035 ;
        RECT 98.965 54.485 99.295 54.865 ;
        RECT 99.475 54.655 99.735 55.160 ;
        RECT 99.995 55.035 100.660 55.205 ;
        RECT 99.995 54.745 100.165 55.035 ;
        RECT 100.335 54.485 100.665 54.865 ;
        RECT 100.835 54.745 101.060 56.865 ;
        RECT 101.275 56.535 101.605 57.035 ;
        RECT 101.775 56.365 101.945 56.865 ;
        RECT 102.180 56.650 103.010 56.820 ;
        RECT 103.250 56.655 103.630 57.035 ;
        RECT 101.250 56.195 101.945 56.365 ;
        RECT 101.250 55.225 101.420 56.195 ;
        RECT 101.590 55.405 102.000 56.025 ;
        RECT 102.170 55.975 102.670 56.355 ;
        RECT 101.250 55.035 101.945 55.225 ;
        RECT 102.170 55.105 102.390 55.975 ;
        RECT 102.840 55.805 103.010 56.650 ;
        RECT 103.810 56.485 103.980 56.775 ;
        RECT 104.150 56.655 104.480 57.035 ;
        RECT 104.950 56.565 105.580 56.815 ;
        RECT 105.760 56.655 106.180 57.035 ;
        RECT 105.410 56.485 105.580 56.565 ;
        RECT 106.380 56.485 106.620 56.775 ;
        RECT 103.180 56.235 104.550 56.485 ;
        RECT 103.180 55.975 103.430 56.235 ;
        RECT 103.940 55.805 104.190 55.965 ;
        RECT 102.840 55.635 104.190 55.805 ;
        RECT 102.840 55.595 103.260 55.635 ;
        RECT 102.570 55.045 102.920 55.415 ;
        RECT 101.275 54.485 101.605 54.865 ;
        RECT 101.775 54.705 101.945 55.035 ;
        RECT 103.090 54.865 103.260 55.595 ;
        RECT 104.360 55.465 104.550 56.235 ;
        RECT 103.430 55.135 103.840 55.465 ;
        RECT 104.130 55.125 104.550 55.465 ;
        RECT 104.720 56.055 105.240 56.365 ;
        RECT 105.410 56.315 106.620 56.485 ;
        RECT 106.850 56.345 107.180 57.035 ;
        RECT 104.720 55.295 104.890 56.055 ;
        RECT 105.060 55.465 105.240 55.875 ;
        RECT 105.410 55.805 105.580 56.315 ;
        RECT 107.350 56.165 107.520 56.775 ;
        RECT 107.790 56.315 108.120 56.825 ;
        RECT 107.350 56.145 107.670 56.165 ;
        RECT 105.750 55.975 107.670 56.145 ;
        RECT 105.410 55.635 107.310 55.805 ;
        RECT 105.640 55.295 105.970 55.415 ;
        RECT 104.720 55.125 105.970 55.295 ;
        RECT 102.245 54.665 103.260 54.865 ;
        RECT 103.430 54.485 103.840 54.925 ;
        RECT 104.130 54.695 104.380 55.125 ;
        RECT 104.580 54.485 104.900 54.945 ;
        RECT 106.140 54.875 106.310 55.635 ;
        RECT 106.980 55.575 107.310 55.635 ;
        RECT 106.500 55.405 106.830 55.465 ;
        RECT 106.500 55.135 107.160 55.405 ;
        RECT 107.480 55.080 107.670 55.975 ;
        RECT 105.460 54.705 106.310 54.875 ;
        RECT 106.510 54.485 107.170 54.965 ;
        RECT 107.350 54.750 107.670 55.080 ;
        RECT 107.870 55.725 108.120 56.315 ;
        RECT 108.300 56.235 108.585 57.035 ;
        RECT 108.765 56.695 109.020 56.725 ;
        RECT 108.765 56.525 109.105 56.695 ;
        RECT 108.765 56.055 109.020 56.525 ;
        RECT 107.870 55.395 108.670 55.725 ;
        RECT 107.870 54.745 108.120 55.395 ;
        RECT 108.840 55.195 109.020 56.055 ;
        RECT 109.605 55.895 109.835 57.035 ;
        RECT 110.005 55.885 110.335 56.865 ;
        RECT 110.505 55.895 110.715 57.035 ;
        RECT 110.945 55.945 112.155 57.035 ;
        RECT 109.585 55.475 109.915 55.725 ;
        RECT 108.300 54.485 108.585 54.945 ;
        RECT 108.765 54.665 109.020 55.195 ;
        RECT 109.605 54.485 109.835 55.305 ;
        RECT 110.085 55.285 110.335 55.885 ;
        RECT 110.005 54.655 110.335 55.285 ;
        RECT 110.505 54.485 110.715 55.305 ;
        RECT 110.945 55.235 111.465 55.775 ;
        RECT 111.635 55.405 112.155 55.945 ;
        RECT 112.325 55.945 113.535 57.035 ;
        RECT 112.325 55.405 112.845 55.945 ;
        RECT 113.015 55.235 113.535 55.775 ;
        RECT 110.945 54.485 112.155 55.235 ;
        RECT 112.325 54.485 113.535 55.235 ;
        RECT 5.520 54.315 113.620 54.485 ;
        RECT 5.605 53.565 6.815 54.315 ;
        RECT 6.985 53.565 8.195 54.315 ;
        RECT 8.370 53.765 8.625 54.055 ;
        RECT 8.795 53.935 9.125 54.315 ;
        RECT 8.370 53.595 9.120 53.765 ;
        RECT 5.605 53.025 6.125 53.565 ;
        RECT 6.295 52.855 6.815 53.395 ;
        RECT 6.985 53.025 7.505 53.565 ;
        RECT 7.675 52.855 8.195 53.395 ;
        RECT 5.605 51.765 6.815 52.855 ;
        RECT 6.985 51.765 8.195 52.855 ;
        RECT 8.370 52.775 8.720 53.425 ;
        RECT 8.890 52.605 9.120 53.595 ;
        RECT 8.370 52.435 9.120 52.605 ;
        RECT 8.370 51.935 8.625 52.435 ;
        RECT 8.795 51.765 9.125 52.265 ;
        RECT 9.295 51.935 9.465 54.055 ;
        RECT 9.825 53.955 10.155 54.315 ;
        RECT 10.325 53.925 10.820 54.095 ;
        RECT 11.025 53.925 11.880 54.095 ;
        RECT 9.695 52.735 10.155 53.785 ;
        RECT 9.635 51.950 9.960 52.735 ;
        RECT 10.325 52.565 10.495 53.925 ;
        RECT 10.665 53.015 11.015 53.635 ;
        RECT 11.185 53.415 11.540 53.635 ;
        RECT 11.185 52.825 11.355 53.415 ;
        RECT 11.710 53.215 11.880 53.925 ;
        RECT 12.755 53.855 13.085 54.315 ;
        RECT 13.295 53.955 13.645 54.125 ;
        RECT 12.085 53.385 12.875 53.635 ;
        RECT 13.295 53.565 13.555 53.955 ;
        RECT 13.865 53.865 14.815 54.145 ;
        RECT 14.985 53.875 15.175 54.315 ;
        RECT 15.345 53.935 16.415 54.105 ;
        RECT 13.045 53.215 13.215 53.395 ;
        RECT 10.325 52.395 10.720 52.565 ;
        RECT 10.890 52.435 11.355 52.825 ;
        RECT 11.525 53.045 13.215 53.215 ;
        RECT 10.550 52.265 10.720 52.395 ;
        RECT 11.525 52.265 11.695 53.045 ;
        RECT 13.385 52.875 13.555 53.565 ;
        RECT 12.055 52.705 13.555 52.875 ;
        RECT 13.745 52.905 13.955 53.695 ;
        RECT 14.125 53.075 14.475 53.695 ;
        RECT 14.645 53.085 14.815 53.865 ;
        RECT 15.345 53.705 15.515 53.935 ;
        RECT 14.985 53.535 15.515 53.705 ;
        RECT 14.985 53.255 15.205 53.535 ;
        RECT 15.685 53.365 15.925 53.765 ;
        RECT 14.645 52.915 15.050 53.085 ;
        RECT 15.385 52.995 15.925 53.365 ;
        RECT 16.095 53.580 16.415 53.935 ;
        RECT 16.660 53.855 16.965 54.315 ;
        RECT 17.135 53.605 17.390 54.135 ;
        RECT 16.095 53.405 16.420 53.580 ;
        RECT 16.095 53.105 17.010 53.405 ;
        RECT 16.270 53.075 17.010 53.105 ;
        RECT 13.745 52.745 14.420 52.905 ;
        RECT 14.880 52.825 15.050 52.915 ;
        RECT 13.745 52.735 14.710 52.745 ;
        RECT 13.385 52.565 13.555 52.705 ;
        RECT 10.130 51.765 10.380 52.225 ;
        RECT 10.550 51.935 10.800 52.265 ;
        RECT 11.015 51.935 11.695 52.265 ;
        RECT 11.865 52.365 12.940 52.535 ;
        RECT 13.385 52.395 13.945 52.565 ;
        RECT 14.250 52.445 14.710 52.735 ;
        RECT 14.880 52.655 16.100 52.825 ;
        RECT 11.865 52.025 12.035 52.365 ;
        RECT 12.270 51.765 12.600 52.195 ;
        RECT 12.770 52.025 12.940 52.365 ;
        RECT 13.235 51.765 13.605 52.225 ;
        RECT 13.775 51.935 13.945 52.395 ;
        RECT 14.880 52.275 15.050 52.655 ;
        RECT 16.270 52.485 16.440 53.075 ;
        RECT 17.180 52.955 17.390 53.605 ;
        RECT 18.030 53.765 18.285 54.055 ;
        RECT 18.455 53.935 18.785 54.315 ;
        RECT 18.030 53.595 18.780 53.765 ;
        RECT 14.180 51.935 15.050 52.275 ;
        RECT 15.640 52.315 16.440 52.485 ;
        RECT 15.220 51.765 15.470 52.225 ;
        RECT 15.640 52.025 15.810 52.315 ;
        RECT 15.990 51.765 16.320 52.145 ;
        RECT 16.660 51.765 16.965 52.905 ;
        RECT 17.135 52.075 17.390 52.955 ;
        RECT 18.030 52.775 18.380 53.425 ;
        RECT 18.550 52.605 18.780 53.595 ;
        RECT 18.030 52.435 18.780 52.605 ;
        RECT 18.030 51.935 18.285 52.435 ;
        RECT 18.455 51.765 18.785 52.265 ;
        RECT 18.955 51.935 19.125 54.055 ;
        RECT 19.485 53.955 19.815 54.315 ;
        RECT 19.985 53.925 20.480 54.095 ;
        RECT 20.685 53.925 21.540 54.095 ;
        RECT 19.355 52.735 19.815 53.785 ;
        RECT 19.295 51.950 19.620 52.735 ;
        RECT 19.985 52.565 20.155 53.925 ;
        RECT 20.325 53.015 20.675 53.635 ;
        RECT 20.845 53.415 21.200 53.635 ;
        RECT 20.845 52.825 21.015 53.415 ;
        RECT 21.370 53.215 21.540 53.925 ;
        RECT 22.415 53.855 22.745 54.315 ;
        RECT 22.955 53.955 23.305 54.125 ;
        RECT 21.745 53.385 22.535 53.635 ;
        RECT 22.955 53.565 23.215 53.955 ;
        RECT 23.525 53.865 24.475 54.145 ;
        RECT 24.645 53.875 24.835 54.315 ;
        RECT 25.005 53.935 26.075 54.105 ;
        RECT 22.705 53.215 22.875 53.395 ;
        RECT 19.985 52.395 20.380 52.565 ;
        RECT 20.550 52.435 21.015 52.825 ;
        RECT 21.185 53.045 22.875 53.215 ;
        RECT 20.210 52.265 20.380 52.395 ;
        RECT 21.185 52.265 21.355 53.045 ;
        RECT 23.045 52.875 23.215 53.565 ;
        RECT 21.715 52.705 23.215 52.875 ;
        RECT 23.405 52.905 23.615 53.695 ;
        RECT 23.785 53.075 24.135 53.695 ;
        RECT 24.305 53.085 24.475 53.865 ;
        RECT 25.005 53.705 25.175 53.935 ;
        RECT 24.645 53.535 25.175 53.705 ;
        RECT 24.645 53.255 24.865 53.535 ;
        RECT 25.345 53.365 25.585 53.765 ;
        RECT 24.305 52.915 24.710 53.085 ;
        RECT 25.045 52.995 25.585 53.365 ;
        RECT 25.755 53.580 26.075 53.935 ;
        RECT 26.320 53.855 26.625 54.315 ;
        RECT 26.795 53.605 27.050 54.135 ;
        RECT 25.755 53.405 26.080 53.580 ;
        RECT 25.755 53.105 26.670 53.405 ;
        RECT 25.930 53.075 26.670 53.105 ;
        RECT 23.405 52.745 24.080 52.905 ;
        RECT 24.540 52.825 24.710 52.915 ;
        RECT 23.405 52.735 24.370 52.745 ;
        RECT 23.045 52.565 23.215 52.705 ;
        RECT 19.790 51.765 20.040 52.225 ;
        RECT 20.210 51.935 20.460 52.265 ;
        RECT 20.675 51.935 21.355 52.265 ;
        RECT 21.525 52.365 22.600 52.535 ;
        RECT 23.045 52.395 23.605 52.565 ;
        RECT 23.910 52.445 24.370 52.735 ;
        RECT 24.540 52.655 25.760 52.825 ;
        RECT 21.525 52.025 21.695 52.365 ;
        RECT 21.930 51.765 22.260 52.195 ;
        RECT 22.430 52.025 22.600 52.365 ;
        RECT 22.895 51.765 23.265 52.225 ;
        RECT 23.435 51.935 23.605 52.395 ;
        RECT 24.540 52.275 24.710 52.655 ;
        RECT 25.930 52.485 26.100 53.075 ;
        RECT 26.840 52.955 27.050 53.605 ;
        RECT 23.840 51.935 24.710 52.275 ;
        RECT 25.300 52.315 26.100 52.485 ;
        RECT 24.880 51.765 25.130 52.225 ;
        RECT 25.300 52.025 25.470 52.315 ;
        RECT 25.650 51.765 25.980 52.145 ;
        RECT 26.320 51.765 26.625 52.905 ;
        RECT 26.795 52.075 27.050 52.955 ;
        RECT 27.225 53.640 27.485 54.145 ;
        RECT 27.665 53.935 27.995 54.315 ;
        RECT 28.175 53.765 28.345 54.145 ;
        RECT 27.225 52.840 27.395 53.640 ;
        RECT 27.680 53.595 28.345 53.765 ;
        RECT 27.680 53.340 27.850 53.595 ;
        RECT 28.665 53.495 28.875 54.315 ;
        RECT 29.045 53.515 29.375 54.145 ;
        RECT 27.565 53.010 27.850 53.340 ;
        RECT 28.085 53.045 28.415 53.415 ;
        RECT 27.680 52.865 27.850 53.010 ;
        RECT 29.045 52.915 29.295 53.515 ;
        RECT 29.545 53.495 29.775 54.315 ;
        RECT 29.985 53.565 31.195 54.315 ;
        RECT 31.365 53.590 31.655 54.315 ;
        RECT 29.465 53.075 29.795 53.325 ;
        RECT 29.985 53.025 30.505 53.565 ;
        RECT 31.885 53.495 32.095 54.315 ;
        RECT 32.265 53.515 32.595 54.145 ;
        RECT 27.225 51.935 27.495 52.840 ;
        RECT 27.680 52.695 28.345 52.865 ;
        RECT 27.665 51.765 27.995 52.525 ;
        RECT 28.175 51.935 28.345 52.695 ;
        RECT 28.665 51.765 28.875 52.905 ;
        RECT 29.045 51.935 29.375 52.915 ;
        RECT 29.545 51.765 29.775 52.905 ;
        RECT 30.675 52.855 31.195 53.395 ;
        RECT 29.985 51.765 31.195 52.855 ;
        RECT 31.365 51.765 31.655 52.930 ;
        RECT 32.265 52.915 32.515 53.515 ;
        RECT 32.765 53.495 32.995 54.315 ;
        RECT 33.205 53.565 34.415 54.315 ;
        RECT 34.585 53.640 34.845 54.145 ;
        RECT 35.025 53.935 35.355 54.315 ;
        RECT 35.535 53.765 35.705 54.145 ;
        RECT 32.685 53.075 33.015 53.325 ;
        RECT 33.205 53.025 33.725 53.565 ;
        RECT 31.885 51.765 32.095 52.905 ;
        RECT 32.265 51.935 32.595 52.915 ;
        RECT 32.765 51.765 32.995 52.905 ;
        RECT 33.895 52.855 34.415 53.395 ;
        RECT 33.205 51.765 34.415 52.855 ;
        RECT 34.585 52.840 34.755 53.640 ;
        RECT 35.040 53.595 35.705 53.765 ;
        RECT 35.040 53.340 35.210 53.595 ;
        RECT 35.965 53.565 37.175 54.315 ;
        RECT 34.925 53.010 35.210 53.340 ;
        RECT 35.445 53.045 35.775 53.415 ;
        RECT 35.965 53.025 36.485 53.565 ;
        RECT 37.385 53.495 37.615 54.315 ;
        RECT 37.785 53.515 38.115 54.145 ;
        RECT 35.040 52.865 35.210 53.010 ;
        RECT 34.585 51.935 34.855 52.840 ;
        RECT 35.040 52.695 35.705 52.865 ;
        RECT 36.655 52.855 37.175 53.395 ;
        RECT 37.365 53.075 37.695 53.325 ;
        RECT 37.865 52.915 38.115 53.515 ;
        RECT 38.285 53.495 38.495 54.315 ;
        RECT 38.725 53.545 42.235 54.315 ;
        RECT 38.725 53.025 40.375 53.545 ;
        RECT 43.365 53.495 43.595 54.315 ;
        RECT 43.765 53.515 44.095 54.145 ;
        RECT 35.025 51.765 35.355 52.525 ;
        RECT 35.535 51.935 35.705 52.695 ;
        RECT 35.965 51.765 37.175 52.855 ;
        RECT 37.385 51.765 37.615 52.905 ;
        RECT 37.785 51.935 38.115 52.915 ;
        RECT 38.285 51.765 38.495 52.905 ;
        RECT 40.545 52.855 42.235 53.375 ;
        RECT 43.345 53.075 43.675 53.325 ;
        RECT 43.845 52.915 44.095 53.515 ;
        RECT 44.265 53.495 44.475 54.315 ;
        RECT 44.795 53.765 44.965 54.055 ;
        RECT 45.135 53.935 45.465 54.315 ;
        RECT 44.795 53.595 45.460 53.765 ;
        RECT 38.725 51.765 42.235 52.855 ;
        RECT 43.365 51.765 43.595 52.905 ;
        RECT 43.765 51.935 44.095 52.915 ;
        RECT 44.265 51.765 44.475 52.905 ;
        RECT 44.710 52.775 45.060 53.425 ;
        RECT 45.230 52.605 45.460 53.595 ;
        RECT 44.795 52.435 45.460 52.605 ;
        RECT 44.795 51.935 44.965 52.435 ;
        RECT 45.135 51.765 45.465 52.265 ;
        RECT 45.635 51.935 45.860 54.055 ;
        RECT 46.075 53.935 46.405 54.315 ;
        RECT 46.575 53.765 46.745 54.095 ;
        RECT 47.045 53.935 48.060 54.135 ;
        RECT 46.050 53.575 46.745 53.765 ;
        RECT 46.050 52.605 46.220 53.575 ;
        RECT 46.390 52.775 46.800 53.395 ;
        RECT 46.970 52.825 47.190 53.695 ;
        RECT 47.370 53.385 47.720 53.755 ;
        RECT 47.890 53.205 48.060 53.935 ;
        RECT 48.230 53.875 48.640 54.315 ;
        RECT 48.930 53.675 49.180 54.105 ;
        RECT 49.380 53.855 49.700 54.315 ;
        RECT 50.260 53.925 51.110 54.095 ;
        RECT 48.230 53.335 48.640 53.665 ;
        RECT 48.930 53.335 49.350 53.675 ;
        RECT 47.640 53.165 48.060 53.205 ;
        RECT 47.640 52.995 48.990 53.165 ;
        RECT 46.050 52.435 46.745 52.605 ;
        RECT 46.970 52.445 47.470 52.825 ;
        RECT 46.075 51.765 46.405 52.265 ;
        RECT 46.575 51.935 46.745 52.435 ;
        RECT 47.640 52.150 47.810 52.995 ;
        RECT 48.740 52.835 48.990 52.995 ;
        RECT 47.980 52.565 48.230 52.825 ;
        RECT 49.160 52.565 49.350 53.335 ;
        RECT 47.980 52.315 49.350 52.565 ;
        RECT 49.520 53.505 50.770 53.675 ;
        RECT 49.520 52.745 49.690 53.505 ;
        RECT 50.440 53.385 50.770 53.505 ;
        RECT 49.860 52.925 50.040 53.335 ;
        RECT 50.940 53.165 51.110 53.925 ;
        RECT 51.310 53.835 51.970 54.315 ;
        RECT 52.150 53.720 52.470 54.050 ;
        RECT 51.300 53.395 51.960 53.665 ;
        RECT 51.300 53.335 51.630 53.395 ;
        RECT 51.780 53.165 52.110 53.225 ;
        RECT 50.210 52.995 52.110 53.165 ;
        RECT 49.520 52.435 50.040 52.745 ;
        RECT 50.210 52.485 50.380 52.995 ;
        RECT 52.280 52.825 52.470 53.720 ;
        RECT 50.550 52.655 52.470 52.825 ;
        RECT 52.150 52.635 52.470 52.655 ;
        RECT 52.670 53.405 52.920 54.055 ;
        RECT 53.100 53.855 53.385 54.315 ;
        RECT 53.565 53.975 53.820 54.135 ;
        RECT 53.565 53.805 53.905 53.975 ;
        RECT 54.425 53.835 54.705 54.315 ;
        RECT 53.565 53.605 53.820 53.805 ;
        RECT 54.875 53.665 55.135 54.055 ;
        RECT 55.310 53.835 55.565 54.315 ;
        RECT 55.735 53.665 56.030 54.055 ;
        RECT 56.210 53.835 56.485 54.315 ;
        RECT 56.655 53.815 56.955 54.145 ;
        RECT 52.670 53.075 53.470 53.405 ;
        RECT 50.210 52.315 51.420 52.485 ;
        RECT 46.980 51.980 47.810 52.150 ;
        RECT 48.050 51.765 48.430 52.145 ;
        RECT 48.610 52.025 48.780 52.315 ;
        RECT 50.210 52.235 50.380 52.315 ;
        RECT 48.950 51.765 49.280 52.145 ;
        RECT 49.750 51.985 50.380 52.235 ;
        RECT 50.560 51.765 50.980 52.145 ;
        RECT 51.180 52.025 51.420 52.315 ;
        RECT 51.650 51.765 51.980 52.455 ;
        RECT 52.150 52.025 52.320 52.635 ;
        RECT 52.670 52.485 52.920 53.075 ;
        RECT 53.640 52.745 53.820 53.605 ;
        RECT 54.380 53.495 56.030 53.665 ;
        RECT 54.380 52.985 54.785 53.495 ;
        RECT 54.955 53.155 56.095 53.325 ;
        RECT 54.380 52.815 55.135 52.985 ;
        RECT 52.590 51.975 52.920 52.485 ;
        RECT 53.100 51.765 53.385 52.565 ;
        RECT 53.565 52.075 53.820 52.745 ;
        RECT 54.420 51.765 54.705 52.635 ;
        RECT 54.875 52.565 55.135 52.815 ;
        RECT 55.925 52.905 56.095 53.155 ;
        RECT 56.265 53.075 56.615 53.645 ;
        RECT 56.785 52.905 56.955 53.815 ;
        RECT 57.125 53.590 57.415 54.315 ;
        RECT 57.585 53.545 59.255 54.315 ;
        RECT 59.515 53.665 59.685 54.145 ;
        RECT 59.865 53.835 60.105 54.315 ;
        RECT 60.355 53.665 60.525 54.145 ;
        RECT 60.695 53.835 61.025 54.315 ;
        RECT 61.195 53.665 61.365 54.145 ;
        RECT 57.585 53.025 58.335 53.545 ;
        RECT 59.515 53.495 60.150 53.665 ;
        RECT 60.355 53.495 61.365 53.665 ;
        RECT 61.535 53.515 61.865 54.315 ;
        RECT 62.185 53.815 62.485 54.145 ;
        RECT 62.655 53.835 62.930 54.315 ;
        RECT 55.925 52.735 56.955 52.905 ;
        RECT 54.875 52.395 55.995 52.565 ;
        RECT 54.875 51.935 55.135 52.395 ;
        RECT 55.310 51.765 55.565 52.225 ;
        RECT 55.735 51.935 55.995 52.395 ;
        RECT 56.165 51.765 56.475 52.565 ;
        RECT 56.645 51.935 56.955 52.735 ;
        RECT 57.125 51.765 57.415 52.930 ;
        RECT 58.505 52.855 59.255 53.375 ;
        RECT 59.980 53.325 60.150 53.495 ;
        RECT 59.430 53.085 59.810 53.325 ;
        RECT 59.980 53.155 60.480 53.325 ;
        RECT 59.980 52.915 60.150 53.155 ;
        RECT 60.870 52.955 61.365 53.495 ;
        RECT 57.585 51.765 59.255 52.855 ;
        RECT 59.435 52.745 60.150 52.915 ;
        RECT 60.355 52.785 61.365 52.955 ;
        RECT 59.435 51.935 59.765 52.745 ;
        RECT 59.935 51.765 60.175 52.565 ;
        RECT 60.355 51.935 60.525 52.785 ;
        RECT 60.695 51.765 61.025 52.565 ;
        RECT 61.195 51.935 61.365 52.785 ;
        RECT 61.535 51.765 61.865 52.915 ;
        RECT 62.185 52.905 62.355 53.815 ;
        RECT 63.110 53.665 63.405 54.055 ;
        RECT 63.575 53.835 63.830 54.315 ;
        RECT 64.005 53.665 64.265 54.055 ;
        RECT 64.435 53.835 64.715 54.315 ;
        RECT 65.495 53.665 65.665 54.145 ;
        RECT 65.845 53.835 66.085 54.315 ;
        RECT 66.335 53.665 66.505 54.145 ;
        RECT 66.675 53.835 67.005 54.315 ;
        RECT 67.175 53.665 67.345 54.145 ;
        RECT 62.525 53.075 62.875 53.645 ;
        RECT 63.110 53.495 64.760 53.665 ;
        RECT 65.495 53.495 66.130 53.665 ;
        RECT 66.335 53.495 67.345 53.665 ;
        RECT 67.515 53.515 67.845 54.315 ;
        RECT 68.165 53.545 70.755 54.315 ;
        RECT 63.045 53.155 64.185 53.325 ;
        RECT 63.045 52.905 63.215 53.155 ;
        RECT 64.355 52.985 64.760 53.495 ;
        RECT 65.960 53.325 66.130 53.495 ;
        RECT 65.410 53.085 65.790 53.325 ;
        RECT 65.960 53.155 66.460 53.325 ;
        RECT 62.185 52.735 63.215 52.905 ;
        RECT 64.005 52.815 64.760 52.985 ;
        RECT 65.960 52.915 66.130 53.155 ;
        RECT 66.850 52.955 67.345 53.495 ;
        RECT 68.165 53.025 69.375 53.545 ;
        RECT 70.965 53.495 71.195 54.315 ;
        RECT 71.365 53.515 71.695 54.145 ;
        RECT 62.185 51.935 62.495 52.735 ;
        RECT 64.005 52.565 64.265 52.815 ;
        RECT 65.415 52.745 66.130 52.915 ;
        RECT 66.335 52.785 67.345 52.955 ;
        RECT 62.665 51.765 62.975 52.565 ;
        RECT 63.145 52.395 64.265 52.565 ;
        RECT 63.145 51.935 63.405 52.395 ;
        RECT 63.575 51.765 63.830 52.225 ;
        RECT 64.005 51.935 64.265 52.395 ;
        RECT 64.435 51.765 64.720 52.635 ;
        RECT 65.415 51.935 65.745 52.745 ;
        RECT 65.915 51.765 66.155 52.565 ;
        RECT 66.335 51.935 66.505 52.785 ;
        RECT 66.675 51.765 67.005 52.565 ;
        RECT 67.175 51.935 67.345 52.785 ;
        RECT 67.515 51.765 67.845 52.915 ;
        RECT 69.545 52.855 70.755 53.375 ;
        RECT 70.945 53.075 71.275 53.325 ;
        RECT 71.445 52.915 71.695 53.515 ;
        RECT 71.865 53.495 72.075 54.315 ;
        RECT 72.310 53.605 72.565 54.135 ;
        RECT 72.735 53.855 73.040 54.315 ;
        RECT 73.285 53.935 74.355 54.105 ;
        RECT 68.165 51.765 70.755 52.855 ;
        RECT 70.965 51.765 71.195 52.905 ;
        RECT 71.365 51.935 71.695 52.915 ;
        RECT 72.310 52.955 72.520 53.605 ;
        RECT 73.285 53.580 73.605 53.935 ;
        RECT 73.280 53.405 73.605 53.580 ;
        RECT 72.690 53.105 73.605 53.405 ;
        RECT 73.775 53.365 74.015 53.765 ;
        RECT 74.185 53.705 74.355 53.935 ;
        RECT 74.525 53.875 74.715 54.315 ;
        RECT 74.885 53.865 75.835 54.145 ;
        RECT 76.055 53.955 76.405 54.125 ;
        RECT 74.185 53.535 74.715 53.705 ;
        RECT 72.690 53.075 73.430 53.105 ;
        RECT 71.865 51.765 72.075 52.905 ;
        RECT 72.310 52.075 72.565 52.955 ;
        RECT 72.735 51.765 73.040 52.905 ;
        RECT 73.260 52.485 73.430 53.075 ;
        RECT 73.775 52.995 74.315 53.365 ;
        RECT 74.495 53.255 74.715 53.535 ;
        RECT 74.885 53.085 75.055 53.865 ;
        RECT 74.650 52.915 75.055 53.085 ;
        RECT 75.225 53.075 75.575 53.695 ;
        RECT 74.650 52.825 74.820 52.915 ;
        RECT 75.745 52.905 75.955 53.695 ;
        RECT 73.600 52.655 74.820 52.825 ;
        RECT 75.280 52.745 75.955 52.905 ;
        RECT 73.260 52.315 74.060 52.485 ;
        RECT 73.380 51.765 73.710 52.145 ;
        RECT 73.890 52.025 74.060 52.315 ;
        RECT 74.650 52.275 74.820 52.655 ;
        RECT 74.990 52.735 75.955 52.745 ;
        RECT 76.145 53.565 76.405 53.955 ;
        RECT 76.615 53.855 76.945 54.315 ;
        RECT 77.820 53.925 78.675 54.095 ;
        RECT 78.880 53.925 79.375 54.095 ;
        RECT 79.545 53.955 79.875 54.315 ;
        RECT 76.145 52.875 76.315 53.565 ;
        RECT 76.485 53.215 76.655 53.395 ;
        RECT 76.825 53.385 77.615 53.635 ;
        RECT 77.820 53.215 77.990 53.925 ;
        RECT 78.160 53.415 78.515 53.635 ;
        RECT 76.485 53.045 78.175 53.215 ;
        RECT 74.990 52.445 75.450 52.735 ;
        RECT 76.145 52.705 77.645 52.875 ;
        RECT 76.145 52.565 76.315 52.705 ;
        RECT 75.755 52.395 76.315 52.565 ;
        RECT 74.230 51.765 74.480 52.225 ;
        RECT 74.650 51.935 75.520 52.275 ;
        RECT 75.755 51.935 75.925 52.395 ;
        RECT 76.760 52.365 77.835 52.535 ;
        RECT 76.095 51.765 76.465 52.225 ;
        RECT 76.760 52.025 76.930 52.365 ;
        RECT 77.100 51.765 77.430 52.195 ;
        RECT 77.665 52.025 77.835 52.365 ;
        RECT 78.005 52.265 78.175 53.045 ;
        RECT 78.345 52.825 78.515 53.415 ;
        RECT 78.685 53.015 79.035 53.635 ;
        RECT 78.345 52.435 78.810 52.825 ;
        RECT 79.205 52.565 79.375 53.925 ;
        RECT 79.545 52.735 80.005 53.785 ;
        RECT 78.980 52.395 79.375 52.565 ;
        RECT 78.980 52.265 79.150 52.395 ;
        RECT 78.005 51.935 78.685 52.265 ;
        RECT 78.900 51.935 79.150 52.265 ;
        RECT 79.320 51.765 79.570 52.225 ;
        RECT 79.740 51.950 80.065 52.735 ;
        RECT 80.235 51.935 80.405 54.055 ;
        RECT 80.575 53.935 80.905 54.315 ;
        RECT 81.075 53.765 81.330 54.055 ;
        RECT 80.580 53.595 81.330 53.765 ;
        RECT 80.580 52.605 80.810 53.595 ;
        RECT 81.505 53.565 82.715 54.315 ;
        RECT 82.885 53.590 83.175 54.315 ;
        RECT 83.350 53.765 83.605 54.055 ;
        RECT 83.775 53.935 84.105 54.315 ;
        RECT 83.350 53.595 84.100 53.765 ;
        RECT 80.980 52.775 81.330 53.425 ;
        RECT 81.505 53.025 82.025 53.565 ;
        RECT 82.195 52.855 82.715 53.395 ;
        RECT 80.580 52.435 81.330 52.605 ;
        RECT 80.575 51.765 80.905 52.265 ;
        RECT 81.075 51.935 81.330 52.435 ;
        RECT 81.505 51.765 82.715 52.855 ;
        RECT 82.885 51.765 83.175 52.930 ;
        RECT 83.350 52.775 83.700 53.425 ;
        RECT 83.870 52.605 84.100 53.595 ;
        RECT 83.350 52.435 84.100 52.605 ;
        RECT 83.350 51.935 83.605 52.435 ;
        RECT 83.775 51.765 84.105 52.265 ;
        RECT 84.275 51.935 84.445 54.055 ;
        RECT 84.805 53.955 85.135 54.315 ;
        RECT 85.305 53.925 85.800 54.095 ;
        RECT 86.005 53.925 86.860 54.095 ;
        RECT 84.675 52.735 85.135 53.785 ;
        RECT 84.615 51.950 84.940 52.735 ;
        RECT 85.305 52.565 85.475 53.925 ;
        RECT 85.645 53.015 85.995 53.635 ;
        RECT 86.165 53.415 86.520 53.635 ;
        RECT 86.165 52.825 86.335 53.415 ;
        RECT 86.690 53.215 86.860 53.925 ;
        RECT 87.735 53.855 88.065 54.315 ;
        RECT 88.275 53.955 88.625 54.125 ;
        RECT 87.065 53.385 87.855 53.635 ;
        RECT 88.275 53.565 88.535 53.955 ;
        RECT 88.845 53.865 89.795 54.145 ;
        RECT 89.965 53.875 90.155 54.315 ;
        RECT 90.325 53.935 91.395 54.105 ;
        RECT 88.025 53.215 88.195 53.395 ;
        RECT 85.305 52.395 85.700 52.565 ;
        RECT 85.870 52.435 86.335 52.825 ;
        RECT 86.505 53.045 88.195 53.215 ;
        RECT 85.530 52.265 85.700 52.395 ;
        RECT 86.505 52.265 86.675 53.045 ;
        RECT 88.365 52.875 88.535 53.565 ;
        RECT 87.035 52.705 88.535 52.875 ;
        RECT 88.725 52.905 88.935 53.695 ;
        RECT 89.105 53.075 89.455 53.695 ;
        RECT 89.625 53.085 89.795 53.865 ;
        RECT 90.325 53.705 90.495 53.935 ;
        RECT 89.965 53.535 90.495 53.705 ;
        RECT 89.965 53.255 90.185 53.535 ;
        RECT 90.665 53.365 90.905 53.765 ;
        RECT 89.625 52.915 90.030 53.085 ;
        RECT 90.365 52.995 90.905 53.365 ;
        RECT 91.075 53.580 91.395 53.935 ;
        RECT 91.640 53.855 91.945 54.315 ;
        RECT 92.115 53.605 92.370 54.135 ;
        RECT 91.075 53.405 91.400 53.580 ;
        RECT 91.075 53.105 91.990 53.405 ;
        RECT 91.250 53.075 91.990 53.105 ;
        RECT 88.725 52.745 89.400 52.905 ;
        RECT 89.860 52.825 90.030 52.915 ;
        RECT 88.725 52.735 89.690 52.745 ;
        RECT 88.365 52.565 88.535 52.705 ;
        RECT 85.110 51.765 85.360 52.225 ;
        RECT 85.530 51.935 85.780 52.265 ;
        RECT 85.995 51.935 86.675 52.265 ;
        RECT 86.845 52.365 87.920 52.535 ;
        RECT 88.365 52.395 88.925 52.565 ;
        RECT 89.230 52.445 89.690 52.735 ;
        RECT 89.860 52.655 91.080 52.825 ;
        RECT 86.845 52.025 87.015 52.365 ;
        RECT 87.250 51.765 87.580 52.195 ;
        RECT 87.750 52.025 87.920 52.365 ;
        RECT 88.215 51.765 88.585 52.225 ;
        RECT 88.755 51.935 88.925 52.395 ;
        RECT 89.860 52.275 90.030 52.655 ;
        RECT 91.250 52.485 91.420 53.075 ;
        RECT 92.160 52.955 92.370 53.605 ;
        RECT 92.605 53.495 92.815 54.315 ;
        RECT 92.985 53.515 93.315 54.145 ;
        RECT 89.160 51.935 90.030 52.275 ;
        RECT 90.620 52.315 91.420 52.485 ;
        RECT 90.200 51.765 90.450 52.225 ;
        RECT 90.620 52.025 90.790 52.315 ;
        RECT 90.970 51.765 91.300 52.145 ;
        RECT 91.640 51.765 91.945 52.905 ;
        RECT 92.115 52.075 92.370 52.955 ;
        RECT 92.985 52.915 93.235 53.515 ;
        RECT 93.485 53.495 93.715 54.315 ;
        RECT 94.445 53.495 94.655 54.315 ;
        RECT 94.825 53.515 95.155 54.145 ;
        RECT 93.405 53.075 93.735 53.325 ;
        RECT 94.825 52.915 95.075 53.515 ;
        RECT 95.325 53.495 95.555 54.315 ;
        RECT 95.765 53.545 98.355 54.315 ;
        RECT 99.075 53.765 99.245 54.055 ;
        RECT 99.415 53.935 99.745 54.315 ;
        RECT 99.075 53.595 99.740 53.765 ;
        RECT 95.245 53.075 95.575 53.325 ;
        RECT 95.765 53.025 96.975 53.545 ;
        RECT 92.605 51.765 92.815 52.905 ;
        RECT 92.985 51.935 93.315 52.915 ;
        RECT 93.485 51.765 93.715 52.905 ;
        RECT 94.445 51.765 94.655 52.905 ;
        RECT 94.825 51.935 95.155 52.915 ;
        RECT 95.325 51.765 95.555 52.905 ;
        RECT 97.145 52.855 98.355 53.375 ;
        RECT 95.765 51.765 98.355 52.855 ;
        RECT 98.990 52.775 99.340 53.425 ;
        RECT 99.510 52.605 99.740 53.595 ;
        RECT 99.075 52.435 99.740 52.605 ;
        RECT 99.075 51.935 99.245 52.435 ;
        RECT 99.415 51.765 99.745 52.265 ;
        RECT 99.915 51.935 100.140 54.055 ;
        RECT 100.355 53.935 100.685 54.315 ;
        RECT 100.855 53.765 101.025 54.095 ;
        RECT 101.325 53.935 102.340 54.135 ;
        RECT 100.330 53.575 101.025 53.765 ;
        RECT 100.330 52.605 100.500 53.575 ;
        RECT 100.670 52.775 101.080 53.395 ;
        RECT 101.250 52.825 101.470 53.695 ;
        RECT 101.650 53.385 102.000 53.755 ;
        RECT 102.170 53.205 102.340 53.935 ;
        RECT 102.510 53.875 102.920 54.315 ;
        RECT 103.210 53.675 103.460 54.105 ;
        RECT 103.660 53.855 103.980 54.315 ;
        RECT 104.540 53.925 105.390 54.095 ;
        RECT 102.510 53.335 102.920 53.665 ;
        RECT 103.210 53.335 103.630 53.675 ;
        RECT 101.920 53.165 102.340 53.205 ;
        RECT 101.920 52.995 103.270 53.165 ;
        RECT 100.330 52.435 101.025 52.605 ;
        RECT 101.250 52.445 101.750 52.825 ;
        RECT 100.355 51.765 100.685 52.265 ;
        RECT 100.855 51.935 101.025 52.435 ;
        RECT 101.920 52.150 102.090 52.995 ;
        RECT 103.020 52.835 103.270 52.995 ;
        RECT 102.260 52.565 102.510 52.825 ;
        RECT 103.440 52.565 103.630 53.335 ;
        RECT 102.260 52.315 103.630 52.565 ;
        RECT 103.800 53.505 105.050 53.675 ;
        RECT 103.800 52.745 103.970 53.505 ;
        RECT 104.720 53.385 105.050 53.505 ;
        RECT 104.140 52.925 104.320 53.335 ;
        RECT 105.220 53.165 105.390 53.925 ;
        RECT 105.590 53.835 106.250 54.315 ;
        RECT 106.430 53.720 106.750 54.050 ;
        RECT 105.580 53.395 106.240 53.665 ;
        RECT 105.580 53.335 105.910 53.395 ;
        RECT 106.060 53.165 106.390 53.225 ;
        RECT 104.490 52.995 106.390 53.165 ;
        RECT 103.800 52.435 104.320 52.745 ;
        RECT 104.490 52.485 104.660 52.995 ;
        RECT 106.560 52.825 106.750 53.720 ;
        RECT 104.830 52.655 106.750 52.825 ;
        RECT 106.430 52.635 106.750 52.655 ;
        RECT 106.950 53.405 107.200 54.055 ;
        RECT 107.380 53.855 107.665 54.315 ;
        RECT 107.845 53.605 108.100 54.135 ;
        RECT 106.950 53.075 107.750 53.405 ;
        RECT 104.490 52.315 105.700 52.485 ;
        RECT 101.260 51.980 102.090 52.150 ;
        RECT 102.330 51.765 102.710 52.145 ;
        RECT 102.890 52.025 103.060 52.315 ;
        RECT 104.490 52.235 104.660 52.315 ;
        RECT 103.230 51.765 103.560 52.145 ;
        RECT 104.030 51.985 104.660 52.235 ;
        RECT 104.840 51.765 105.260 52.145 ;
        RECT 105.460 52.025 105.700 52.315 ;
        RECT 105.930 51.765 106.260 52.455 ;
        RECT 106.430 52.025 106.600 52.635 ;
        RECT 106.950 52.485 107.200 53.075 ;
        RECT 107.920 52.745 108.100 53.605 ;
        RECT 108.645 53.590 108.935 54.315 ;
        RECT 109.105 53.545 111.695 54.315 ;
        RECT 112.325 53.565 113.535 54.315 ;
        RECT 109.105 53.025 110.315 53.545 ;
        RECT 106.870 51.975 107.200 52.485 ;
        RECT 107.380 51.765 107.665 52.565 ;
        RECT 107.845 52.275 108.100 52.745 ;
        RECT 107.845 52.105 108.185 52.275 ;
        RECT 107.845 52.075 108.100 52.105 ;
        RECT 108.645 51.765 108.935 52.930 ;
        RECT 110.485 52.855 111.695 53.375 ;
        RECT 109.105 51.765 111.695 52.855 ;
        RECT 112.325 52.855 112.845 53.395 ;
        RECT 113.015 53.025 113.535 53.565 ;
        RECT 112.325 51.765 113.535 52.855 ;
        RECT 5.520 51.595 113.620 51.765 ;
        RECT 5.605 50.505 6.815 51.595 ;
        RECT 5.605 49.795 6.125 50.335 ;
        RECT 6.295 49.965 6.815 50.505 ;
        RECT 7.905 50.625 8.175 51.395 ;
        RECT 8.345 50.815 8.675 51.595 ;
        RECT 8.880 50.990 9.065 51.395 ;
        RECT 9.235 51.170 9.570 51.595 ;
        RECT 8.880 50.815 9.545 50.990 ;
        RECT 7.905 50.455 9.035 50.625 ;
        RECT 5.605 49.045 6.815 49.795 ;
        RECT 7.905 49.545 8.075 50.455 ;
        RECT 8.245 49.705 8.605 50.285 ;
        RECT 8.785 49.955 9.035 50.455 ;
        RECT 9.205 49.785 9.545 50.815 ;
        RECT 9.745 50.835 10.260 51.245 ;
        RECT 10.495 50.835 10.665 51.595 ;
        RECT 10.835 51.255 12.865 51.425 ;
        RECT 9.745 50.025 10.085 50.835 ;
        RECT 10.835 50.590 11.005 51.255 ;
        RECT 11.400 50.915 12.525 51.085 ;
        RECT 10.255 50.400 11.005 50.590 ;
        RECT 11.175 50.575 12.185 50.745 ;
        RECT 9.745 49.855 10.975 50.025 ;
        RECT 8.860 49.615 9.545 49.785 ;
        RECT 7.905 49.215 8.165 49.545 ;
        RECT 8.375 49.045 8.650 49.525 ;
        RECT 8.860 49.215 9.065 49.615 ;
        RECT 9.235 49.045 9.570 49.445 ;
        RECT 10.020 49.250 10.265 49.855 ;
        RECT 10.485 49.045 10.995 49.580 ;
        RECT 11.175 49.215 11.365 50.575 ;
        RECT 11.535 49.555 11.810 50.375 ;
        RECT 12.015 49.775 12.185 50.575 ;
        RECT 12.355 49.785 12.525 50.915 ;
        RECT 12.695 50.285 12.865 51.255 ;
        RECT 13.035 50.455 13.205 51.595 ;
        RECT 13.375 50.455 13.710 51.425 ;
        RECT 12.695 49.955 12.890 50.285 ;
        RECT 13.115 49.955 13.370 50.285 ;
        RECT 13.115 49.785 13.285 49.955 ;
        RECT 13.540 49.785 13.710 50.455 ;
        RECT 12.355 49.615 13.285 49.785 ;
        RECT 12.355 49.580 12.530 49.615 ;
        RECT 11.535 49.385 11.815 49.555 ;
        RECT 11.535 49.215 11.810 49.385 ;
        RECT 12.000 49.215 12.530 49.580 ;
        RECT 12.955 49.045 13.285 49.445 ;
        RECT 13.455 49.215 13.710 49.785 ;
        RECT 13.890 50.455 14.225 51.425 ;
        RECT 14.395 50.455 14.565 51.595 ;
        RECT 14.735 51.255 16.765 51.425 ;
        RECT 13.890 49.785 14.060 50.455 ;
        RECT 14.735 50.285 14.905 51.255 ;
        RECT 14.230 49.955 14.485 50.285 ;
        RECT 14.710 49.955 14.905 50.285 ;
        RECT 15.075 50.915 16.200 51.085 ;
        RECT 14.315 49.785 14.485 49.955 ;
        RECT 15.075 49.785 15.245 50.915 ;
        RECT 13.890 49.215 14.145 49.785 ;
        RECT 14.315 49.615 15.245 49.785 ;
        RECT 15.415 50.575 16.425 50.745 ;
        RECT 15.415 49.775 15.585 50.575 ;
        RECT 15.790 49.895 16.065 50.375 ;
        RECT 15.785 49.725 16.065 49.895 ;
        RECT 15.070 49.580 15.245 49.615 ;
        RECT 14.315 49.045 14.645 49.445 ;
        RECT 15.070 49.215 15.600 49.580 ;
        RECT 15.790 49.215 16.065 49.725 ;
        RECT 16.235 49.215 16.425 50.575 ;
        RECT 16.595 50.590 16.765 51.255 ;
        RECT 16.935 50.835 17.105 51.595 ;
        RECT 17.340 50.835 17.855 51.245 ;
        RECT 16.595 50.400 17.345 50.590 ;
        RECT 17.515 50.025 17.855 50.835 ;
        RECT 18.485 50.430 18.775 51.595 ;
        RECT 19.495 50.850 19.765 51.595 ;
        RECT 20.395 51.590 26.670 51.595 ;
        RECT 19.935 50.680 20.225 51.420 ;
        RECT 20.395 50.865 20.650 51.590 ;
        RECT 20.835 50.695 21.095 51.420 ;
        RECT 21.265 50.865 21.510 51.590 ;
        RECT 21.695 50.695 21.955 51.420 ;
        RECT 22.125 50.865 22.370 51.590 ;
        RECT 22.555 50.695 22.815 51.420 ;
        RECT 22.985 50.865 23.230 51.590 ;
        RECT 23.400 50.695 23.660 51.420 ;
        RECT 23.830 50.865 24.090 51.590 ;
        RECT 24.260 50.695 24.520 51.420 ;
        RECT 24.690 50.865 24.950 51.590 ;
        RECT 25.120 50.695 25.380 51.420 ;
        RECT 25.550 50.865 25.810 51.590 ;
        RECT 25.980 50.695 26.240 51.420 ;
        RECT 26.410 50.795 26.670 51.590 ;
        RECT 20.835 50.680 26.240 50.695 ;
        RECT 19.495 50.455 26.240 50.680 ;
        RECT 16.625 49.855 17.855 50.025 ;
        RECT 19.495 49.865 20.660 50.455 ;
        RECT 26.840 50.285 27.090 51.420 ;
        RECT 27.270 50.785 27.530 51.595 ;
        RECT 27.705 50.285 27.950 51.425 ;
        RECT 28.130 50.785 28.425 51.595 ;
        RECT 28.610 50.455 28.945 51.425 ;
        RECT 29.115 50.455 29.285 51.595 ;
        RECT 29.455 51.255 31.485 51.425 ;
        RECT 20.830 50.035 27.950 50.285 ;
        RECT 16.605 49.045 17.115 49.580 ;
        RECT 17.335 49.250 17.580 49.855 ;
        RECT 18.485 49.045 18.775 49.770 ;
        RECT 19.495 49.695 26.240 49.865 ;
        RECT 19.495 49.045 19.795 49.525 ;
        RECT 19.965 49.240 20.225 49.695 ;
        RECT 20.395 49.045 20.655 49.525 ;
        RECT 20.835 49.240 21.095 49.695 ;
        RECT 21.265 49.045 21.515 49.525 ;
        RECT 21.695 49.240 21.955 49.695 ;
        RECT 22.125 49.045 22.375 49.525 ;
        RECT 22.555 49.240 22.815 49.695 ;
        RECT 22.985 49.045 23.230 49.525 ;
        RECT 23.400 49.240 23.675 49.695 ;
        RECT 23.845 49.045 24.090 49.525 ;
        RECT 24.260 49.240 24.520 49.695 ;
        RECT 24.690 49.045 24.950 49.525 ;
        RECT 25.120 49.240 25.380 49.695 ;
        RECT 25.550 49.045 25.810 49.525 ;
        RECT 25.980 49.240 26.240 49.695 ;
        RECT 26.410 49.045 26.670 49.605 ;
        RECT 26.840 49.225 27.090 50.035 ;
        RECT 27.270 49.045 27.530 49.570 ;
        RECT 27.700 49.225 27.950 50.035 ;
        RECT 28.120 49.725 28.435 50.285 ;
        RECT 28.610 49.785 28.780 50.455 ;
        RECT 29.455 50.285 29.625 51.255 ;
        RECT 28.950 49.955 29.205 50.285 ;
        RECT 29.430 49.955 29.625 50.285 ;
        RECT 29.795 50.915 30.920 51.085 ;
        RECT 29.035 49.785 29.205 49.955 ;
        RECT 29.795 49.785 29.965 50.915 ;
        RECT 28.130 49.045 28.435 49.555 ;
        RECT 28.610 49.215 28.865 49.785 ;
        RECT 29.035 49.615 29.965 49.785 ;
        RECT 30.135 50.575 31.145 50.745 ;
        RECT 30.135 49.775 30.305 50.575 ;
        RECT 30.510 50.235 30.785 50.375 ;
        RECT 30.505 50.065 30.785 50.235 ;
        RECT 29.790 49.580 29.965 49.615 ;
        RECT 29.035 49.045 29.365 49.445 ;
        RECT 29.790 49.215 30.320 49.580 ;
        RECT 30.510 49.215 30.785 50.065 ;
        RECT 30.955 49.215 31.145 50.575 ;
        RECT 31.315 50.590 31.485 51.255 ;
        RECT 31.655 50.835 31.825 51.595 ;
        RECT 32.060 50.835 32.575 51.245 ;
        RECT 31.315 50.400 32.065 50.590 ;
        RECT 32.235 50.025 32.575 50.835 ;
        RECT 32.745 50.505 35.335 51.595 ;
        RECT 31.345 49.855 32.575 50.025 ;
        RECT 31.325 49.045 31.835 49.580 ;
        RECT 32.055 49.250 32.300 49.855 ;
        RECT 32.745 49.815 33.955 50.335 ;
        RECT 34.125 49.985 35.335 50.505 ;
        RECT 35.505 50.520 35.775 51.425 ;
        RECT 35.945 50.835 36.275 51.595 ;
        RECT 36.455 50.665 36.625 51.425 ;
        RECT 32.745 49.045 35.335 49.815 ;
        RECT 35.505 49.720 35.675 50.520 ;
        RECT 35.960 50.495 36.625 50.665 ;
        RECT 35.960 50.350 36.130 50.495 ;
        RECT 35.845 50.020 36.130 50.350 ;
        RECT 36.890 50.455 37.225 51.425 ;
        RECT 37.395 50.455 37.565 51.595 ;
        RECT 37.735 51.255 39.765 51.425 ;
        RECT 35.960 49.765 36.130 50.020 ;
        RECT 36.365 49.945 36.695 50.315 ;
        RECT 36.890 49.785 37.060 50.455 ;
        RECT 37.735 50.285 37.905 51.255 ;
        RECT 37.230 49.955 37.485 50.285 ;
        RECT 37.710 49.955 37.905 50.285 ;
        RECT 38.075 50.915 39.200 51.085 ;
        RECT 37.315 49.785 37.485 49.955 ;
        RECT 38.075 49.785 38.245 50.915 ;
        RECT 35.505 49.215 35.765 49.720 ;
        RECT 35.960 49.595 36.625 49.765 ;
        RECT 35.945 49.045 36.275 49.425 ;
        RECT 36.455 49.215 36.625 49.595 ;
        RECT 36.890 49.215 37.145 49.785 ;
        RECT 37.315 49.615 38.245 49.785 ;
        RECT 38.415 50.575 39.425 50.745 ;
        RECT 38.415 49.775 38.585 50.575 ;
        RECT 38.070 49.580 38.245 49.615 ;
        RECT 37.315 49.045 37.645 49.445 ;
        RECT 38.070 49.215 38.600 49.580 ;
        RECT 38.790 49.555 39.065 50.375 ;
        RECT 38.785 49.385 39.065 49.555 ;
        RECT 38.790 49.215 39.065 49.385 ;
        RECT 39.235 49.215 39.425 50.575 ;
        RECT 39.595 50.590 39.765 51.255 ;
        RECT 39.935 50.835 40.105 51.595 ;
        RECT 40.340 50.835 40.855 51.245 ;
        RECT 39.595 50.400 40.345 50.590 ;
        RECT 40.515 50.025 40.855 50.835 ;
        RECT 41.025 50.505 42.695 51.595 ;
        RECT 39.625 49.855 40.855 50.025 ;
        RECT 39.605 49.045 40.115 49.580 ;
        RECT 40.335 49.250 40.580 49.855 ;
        RECT 41.025 49.815 41.775 50.335 ;
        RECT 41.945 49.985 42.695 50.505 ;
        RECT 42.955 50.665 43.125 51.425 ;
        RECT 43.305 50.835 43.635 51.595 ;
        RECT 42.955 50.495 43.620 50.665 ;
        RECT 43.805 50.520 44.075 51.425 ;
        RECT 43.450 50.350 43.620 50.495 ;
        RECT 42.885 49.945 43.215 50.315 ;
        RECT 43.450 50.020 43.735 50.350 ;
        RECT 41.025 49.045 42.695 49.815 ;
        RECT 43.450 49.765 43.620 50.020 ;
        RECT 42.955 49.595 43.620 49.765 ;
        RECT 43.905 49.720 44.075 50.520 ;
        RECT 44.245 50.430 44.535 51.595 ;
        RECT 44.795 50.925 44.965 51.425 ;
        RECT 45.135 51.095 45.465 51.595 ;
        RECT 44.795 50.755 45.460 50.925 ;
        RECT 44.710 49.935 45.060 50.585 ;
        RECT 42.955 49.215 43.125 49.595 ;
        RECT 43.305 49.045 43.635 49.425 ;
        RECT 43.815 49.215 44.075 49.720 ;
        RECT 44.245 49.045 44.535 49.770 ;
        RECT 45.230 49.765 45.460 50.755 ;
        RECT 44.795 49.595 45.460 49.765 ;
        RECT 44.795 49.305 44.965 49.595 ;
        RECT 45.135 49.045 45.465 49.425 ;
        RECT 45.635 49.305 45.860 51.425 ;
        RECT 46.075 51.095 46.405 51.595 ;
        RECT 46.575 50.925 46.745 51.425 ;
        RECT 46.980 51.210 47.810 51.380 ;
        RECT 48.050 51.215 48.430 51.595 ;
        RECT 46.050 50.755 46.745 50.925 ;
        RECT 46.050 49.785 46.220 50.755 ;
        RECT 46.390 49.965 46.800 50.585 ;
        RECT 46.970 50.535 47.470 50.915 ;
        RECT 46.050 49.595 46.745 49.785 ;
        RECT 46.970 49.665 47.190 50.535 ;
        RECT 47.640 50.365 47.810 51.210 ;
        RECT 48.610 51.045 48.780 51.335 ;
        RECT 48.950 51.215 49.280 51.595 ;
        RECT 49.750 51.125 50.380 51.375 ;
        RECT 50.560 51.215 50.980 51.595 ;
        RECT 50.210 51.045 50.380 51.125 ;
        RECT 51.180 51.045 51.420 51.335 ;
        RECT 47.980 50.795 49.350 51.045 ;
        RECT 47.980 50.535 48.230 50.795 ;
        RECT 48.740 50.365 48.990 50.525 ;
        RECT 47.640 50.195 48.990 50.365 ;
        RECT 47.640 50.155 48.060 50.195 ;
        RECT 47.370 49.605 47.720 49.975 ;
        RECT 46.075 49.045 46.405 49.425 ;
        RECT 46.575 49.265 46.745 49.595 ;
        RECT 47.890 49.425 48.060 50.155 ;
        RECT 49.160 50.025 49.350 50.795 ;
        RECT 48.230 49.695 48.640 50.025 ;
        RECT 48.930 49.685 49.350 50.025 ;
        RECT 49.520 50.615 50.040 50.925 ;
        RECT 50.210 50.875 51.420 51.045 ;
        RECT 51.650 50.905 51.980 51.595 ;
        RECT 49.520 49.855 49.690 50.615 ;
        RECT 49.860 50.025 50.040 50.435 ;
        RECT 50.210 50.365 50.380 50.875 ;
        RECT 52.150 50.725 52.320 51.335 ;
        RECT 52.590 50.875 52.920 51.385 ;
        RECT 52.150 50.705 52.470 50.725 ;
        RECT 50.550 50.535 52.470 50.705 ;
        RECT 50.210 50.195 52.110 50.365 ;
        RECT 50.440 49.855 50.770 49.975 ;
        RECT 49.520 49.685 50.770 49.855 ;
        RECT 47.045 49.225 48.060 49.425 ;
        RECT 48.230 49.045 48.640 49.485 ;
        RECT 48.930 49.255 49.180 49.685 ;
        RECT 49.380 49.045 49.700 49.505 ;
        RECT 50.940 49.435 51.110 50.195 ;
        RECT 51.780 50.135 52.110 50.195 ;
        RECT 51.300 49.965 51.630 50.025 ;
        RECT 51.300 49.695 51.960 49.965 ;
        RECT 52.280 49.640 52.470 50.535 ;
        RECT 50.260 49.265 51.110 49.435 ;
        RECT 51.310 49.045 51.970 49.525 ;
        RECT 52.150 49.310 52.470 49.640 ;
        RECT 52.670 50.285 52.920 50.875 ;
        RECT 53.100 50.795 53.385 51.595 ;
        RECT 53.565 50.615 53.820 51.285 ;
        RECT 52.670 49.955 53.470 50.285 ;
        RECT 52.670 49.305 52.920 49.955 ;
        RECT 53.640 49.755 53.820 50.615 ;
        RECT 54.365 50.505 56.955 51.595 ;
        RECT 53.565 49.555 53.820 49.755 ;
        RECT 54.365 49.815 55.575 50.335 ;
        RECT 55.745 49.985 56.955 50.505 ;
        RECT 57.585 51.005 58.285 51.425 ;
        RECT 58.485 51.235 58.815 51.595 ;
        RECT 58.985 51.005 59.315 51.405 ;
        RECT 57.585 50.775 59.315 51.005 ;
        RECT 53.100 49.045 53.385 49.505 ;
        RECT 53.565 49.385 53.905 49.555 ;
        RECT 53.565 49.225 53.820 49.385 ;
        RECT 54.365 49.045 56.955 49.815 ;
        RECT 57.585 49.805 57.790 50.775 ;
        RECT 57.960 50.035 58.290 50.575 ;
        RECT 58.465 50.285 58.790 50.575 ;
        RECT 58.985 50.555 59.315 50.775 ;
        RECT 59.485 50.285 59.655 51.210 ;
        RECT 59.835 50.535 60.165 51.595 ;
        RECT 60.345 50.505 61.555 51.595 ;
        RECT 61.780 50.725 62.065 51.595 ;
        RECT 62.235 50.965 62.495 51.425 ;
        RECT 62.670 51.135 62.925 51.595 ;
        RECT 63.095 50.965 63.355 51.425 ;
        RECT 62.235 50.795 63.355 50.965 ;
        RECT 63.525 50.795 63.835 51.595 ;
        RECT 62.235 50.545 62.495 50.795 ;
        RECT 62.705 50.745 62.875 50.795 ;
        RECT 64.005 50.625 64.315 51.425 ;
        RECT 64.485 51.160 69.830 51.595 ;
        RECT 58.465 49.955 58.960 50.285 ;
        RECT 59.280 49.955 59.655 50.285 ;
        RECT 59.865 49.955 60.175 50.285 ;
        RECT 57.585 49.215 58.295 49.805 ;
        RECT 60.345 49.795 60.865 50.335 ;
        RECT 61.035 49.965 61.555 50.505 ;
        RECT 61.740 50.375 62.495 50.545 ;
        RECT 63.285 50.455 64.315 50.625 ;
        RECT 61.740 49.865 62.145 50.375 ;
        RECT 63.285 50.205 63.455 50.455 ;
        RECT 62.315 50.035 63.455 50.205 ;
        RECT 58.805 49.575 60.165 49.785 ;
        RECT 58.805 49.215 59.135 49.575 ;
        RECT 59.335 49.045 59.665 49.405 ;
        RECT 59.835 49.215 60.165 49.575 ;
        RECT 60.345 49.045 61.555 49.795 ;
        RECT 61.740 49.695 63.390 49.865 ;
        RECT 63.625 49.715 63.975 50.285 ;
        RECT 61.785 49.045 62.065 49.525 ;
        RECT 62.235 49.305 62.495 49.695 ;
        RECT 62.670 49.045 62.925 49.525 ;
        RECT 63.095 49.305 63.390 49.695 ;
        RECT 64.145 49.545 64.315 50.455 ;
        RECT 66.070 49.590 66.410 50.420 ;
        RECT 67.890 49.910 68.240 51.160 ;
        RECT 70.005 50.430 70.295 51.595 ;
        RECT 70.465 51.160 75.810 51.595 ;
        RECT 63.570 49.045 63.845 49.525 ;
        RECT 64.015 49.215 64.315 49.545 ;
        RECT 64.485 49.045 69.830 49.590 ;
        RECT 70.005 49.045 70.295 49.770 ;
        RECT 72.050 49.590 72.390 50.420 ;
        RECT 73.870 49.910 74.220 51.160 ;
        RECT 76.965 50.455 77.175 51.595 ;
        RECT 77.345 50.445 77.675 51.425 ;
        RECT 77.845 50.455 78.075 51.595 ;
        RECT 78.285 50.505 81.795 51.595 ;
        RECT 81.965 50.505 83.175 51.595 ;
        RECT 70.465 49.045 75.810 49.590 ;
        RECT 76.965 49.045 77.175 49.865 ;
        RECT 77.345 49.845 77.595 50.445 ;
        RECT 77.765 50.035 78.095 50.285 ;
        RECT 77.345 49.215 77.675 49.845 ;
        RECT 77.845 49.045 78.075 49.865 ;
        RECT 78.285 49.815 79.935 50.335 ;
        RECT 80.105 49.985 81.795 50.505 ;
        RECT 78.285 49.045 81.795 49.815 ;
        RECT 81.965 49.795 82.485 50.335 ;
        RECT 82.655 49.965 83.175 50.505 ;
        RECT 83.550 50.625 83.880 51.425 ;
        RECT 84.050 50.795 84.380 51.595 ;
        RECT 84.680 50.625 85.010 51.425 ;
        RECT 85.655 50.795 85.905 51.595 ;
        RECT 83.550 50.455 85.985 50.625 ;
        RECT 86.175 50.455 86.345 51.595 ;
        RECT 86.515 50.455 86.855 51.425 ;
        RECT 87.025 51.160 92.370 51.595 ;
        RECT 83.345 50.035 83.695 50.285 ;
        RECT 83.880 49.825 84.050 50.455 ;
        RECT 84.220 50.035 84.550 50.235 ;
        RECT 84.720 50.035 85.050 50.235 ;
        RECT 85.220 50.035 85.640 50.235 ;
        RECT 85.815 50.205 85.985 50.455 ;
        RECT 85.815 50.035 86.510 50.205 ;
        RECT 81.965 49.045 83.175 49.795 ;
        RECT 83.550 49.215 84.050 49.825 ;
        RECT 84.680 49.695 85.905 49.865 ;
        RECT 86.680 49.845 86.855 50.455 ;
        RECT 84.680 49.215 85.010 49.695 ;
        RECT 85.180 49.045 85.405 49.505 ;
        RECT 85.575 49.215 85.905 49.695 ;
        RECT 86.095 49.045 86.345 49.845 ;
        RECT 86.515 49.215 86.855 49.845 ;
        RECT 88.610 49.590 88.950 50.420 ;
        RECT 90.430 49.910 90.780 51.160 ;
        RECT 92.545 50.505 95.135 51.595 ;
        RECT 92.545 49.815 93.755 50.335 ;
        RECT 93.925 49.985 95.135 50.505 ;
        RECT 95.765 50.430 96.055 51.595 ;
        RECT 96.225 50.505 99.735 51.595 ;
        RECT 99.905 50.505 101.115 51.595 ;
        RECT 96.225 49.815 97.875 50.335 ;
        RECT 98.045 49.985 99.735 50.505 ;
        RECT 87.025 49.045 92.370 49.590 ;
        RECT 92.545 49.045 95.135 49.815 ;
        RECT 95.765 49.045 96.055 49.770 ;
        RECT 96.225 49.045 99.735 49.815 ;
        RECT 99.905 49.795 100.425 50.335 ;
        RECT 100.595 49.965 101.115 50.505 ;
        RECT 101.290 50.455 101.625 51.425 ;
        RECT 101.795 50.455 101.965 51.595 ;
        RECT 102.135 51.255 104.165 51.425 ;
        RECT 99.905 49.045 101.115 49.795 ;
        RECT 101.290 49.785 101.460 50.455 ;
        RECT 102.135 50.285 102.305 51.255 ;
        RECT 101.630 49.955 101.885 50.285 ;
        RECT 102.110 49.955 102.305 50.285 ;
        RECT 102.475 50.915 103.600 51.085 ;
        RECT 101.715 49.785 101.885 49.955 ;
        RECT 102.475 49.785 102.645 50.915 ;
        RECT 101.290 49.215 101.545 49.785 ;
        RECT 101.715 49.615 102.645 49.785 ;
        RECT 102.815 50.575 103.825 50.745 ;
        RECT 102.815 49.775 102.985 50.575 ;
        RECT 103.190 50.235 103.465 50.375 ;
        RECT 103.185 50.065 103.465 50.235 ;
        RECT 102.470 49.580 102.645 49.615 ;
        RECT 101.715 49.045 102.045 49.445 ;
        RECT 102.470 49.215 103.000 49.580 ;
        RECT 103.190 49.215 103.465 50.065 ;
        RECT 103.635 49.215 103.825 50.575 ;
        RECT 103.995 50.590 104.165 51.255 ;
        RECT 104.335 50.835 104.505 51.595 ;
        RECT 104.740 50.835 105.255 51.245 ;
        RECT 105.425 51.160 110.770 51.595 ;
        RECT 103.995 50.400 104.745 50.590 ;
        RECT 104.915 50.025 105.255 50.835 ;
        RECT 104.025 49.855 105.255 50.025 ;
        RECT 104.005 49.045 104.515 49.580 ;
        RECT 104.735 49.250 104.980 49.855 ;
        RECT 107.010 49.590 107.350 50.420 ;
        RECT 108.830 49.910 109.180 51.160 ;
        RECT 110.945 50.505 112.155 51.595 ;
        RECT 110.945 49.795 111.465 50.335 ;
        RECT 111.635 49.965 112.155 50.505 ;
        RECT 112.325 50.505 113.535 51.595 ;
        RECT 112.325 49.965 112.845 50.505 ;
        RECT 113.015 49.795 113.535 50.335 ;
        RECT 105.425 49.045 110.770 49.590 ;
        RECT 110.945 49.045 112.155 49.795 ;
        RECT 112.325 49.045 113.535 49.795 ;
        RECT 5.520 48.875 113.620 49.045 ;
        RECT 5.605 48.125 6.815 48.875 ;
        RECT 6.985 48.125 8.195 48.875 ;
        RECT 8.370 48.165 8.625 48.695 ;
        RECT 8.795 48.415 9.100 48.875 ;
        RECT 9.345 48.495 10.415 48.665 ;
        RECT 5.605 47.585 6.125 48.125 ;
        RECT 6.295 47.415 6.815 47.955 ;
        RECT 6.985 47.585 7.505 48.125 ;
        RECT 7.675 47.415 8.195 47.955 ;
        RECT 5.605 46.325 6.815 47.415 ;
        RECT 6.985 46.325 8.195 47.415 ;
        RECT 8.370 47.515 8.580 48.165 ;
        RECT 9.345 48.140 9.665 48.495 ;
        RECT 9.340 47.965 9.665 48.140 ;
        RECT 8.750 47.665 9.665 47.965 ;
        RECT 9.835 47.925 10.075 48.325 ;
        RECT 10.245 48.265 10.415 48.495 ;
        RECT 10.585 48.435 10.775 48.875 ;
        RECT 10.945 48.425 11.895 48.705 ;
        RECT 12.115 48.515 12.465 48.685 ;
        RECT 10.245 48.095 10.775 48.265 ;
        RECT 8.750 47.635 9.490 47.665 ;
        RECT 8.370 46.635 8.625 47.515 ;
        RECT 8.795 46.325 9.100 47.465 ;
        RECT 9.320 47.045 9.490 47.635 ;
        RECT 9.835 47.555 10.375 47.925 ;
        RECT 10.555 47.815 10.775 48.095 ;
        RECT 10.945 47.645 11.115 48.425 ;
        RECT 10.710 47.475 11.115 47.645 ;
        RECT 11.285 47.635 11.635 48.255 ;
        RECT 10.710 47.385 10.880 47.475 ;
        RECT 11.805 47.465 12.015 48.255 ;
        RECT 9.660 47.215 10.880 47.385 ;
        RECT 11.340 47.305 12.015 47.465 ;
        RECT 9.320 46.875 10.120 47.045 ;
        RECT 9.440 46.325 9.770 46.705 ;
        RECT 9.950 46.585 10.120 46.875 ;
        RECT 10.710 46.835 10.880 47.215 ;
        RECT 11.050 47.295 12.015 47.305 ;
        RECT 12.205 48.125 12.465 48.515 ;
        RECT 12.675 48.415 13.005 48.875 ;
        RECT 13.880 48.485 14.735 48.655 ;
        RECT 14.940 48.485 15.435 48.655 ;
        RECT 15.605 48.515 15.935 48.875 ;
        RECT 12.205 47.435 12.375 48.125 ;
        RECT 12.545 47.775 12.715 47.955 ;
        RECT 12.885 47.945 13.675 48.195 ;
        RECT 13.880 47.775 14.050 48.485 ;
        RECT 14.220 47.975 14.575 48.195 ;
        RECT 12.545 47.605 14.235 47.775 ;
        RECT 11.050 47.005 11.510 47.295 ;
        RECT 12.205 47.265 13.705 47.435 ;
        RECT 12.205 47.125 12.375 47.265 ;
        RECT 11.815 46.955 12.375 47.125 ;
        RECT 10.290 46.325 10.540 46.785 ;
        RECT 10.710 46.495 11.580 46.835 ;
        RECT 11.815 46.495 11.985 46.955 ;
        RECT 12.820 46.925 13.895 47.095 ;
        RECT 12.155 46.325 12.525 46.785 ;
        RECT 12.820 46.585 12.990 46.925 ;
        RECT 13.160 46.325 13.490 46.755 ;
        RECT 13.725 46.585 13.895 46.925 ;
        RECT 14.065 46.825 14.235 47.605 ;
        RECT 14.405 47.385 14.575 47.975 ;
        RECT 14.745 47.575 15.095 48.195 ;
        RECT 14.405 46.995 14.870 47.385 ;
        RECT 15.265 47.125 15.435 48.485 ;
        RECT 15.605 47.295 16.065 48.345 ;
        RECT 15.040 46.955 15.435 47.125 ;
        RECT 15.040 46.825 15.210 46.955 ;
        RECT 14.065 46.495 14.745 46.825 ;
        RECT 14.960 46.495 15.210 46.825 ;
        RECT 15.380 46.325 15.630 46.785 ;
        RECT 15.800 46.510 16.125 47.295 ;
        RECT 16.295 46.495 16.465 48.615 ;
        RECT 16.635 48.495 16.965 48.875 ;
        RECT 17.135 48.325 17.390 48.615 ;
        RECT 16.640 48.155 17.390 48.325 ;
        RECT 18.115 48.325 18.285 48.705 ;
        RECT 18.465 48.495 18.795 48.875 ;
        RECT 18.115 48.155 18.780 48.325 ;
        RECT 18.975 48.200 19.235 48.705 ;
        RECT 16.640 47.165 16.870 48.155 ;
        RECT 17.040 47.335 17.390 47.985 ;
        RECT 18.045 47.605 18.375 47.975 ;
        RECT 18.610 47.900 18.780 48.155 ;
        RECT 18.610 47.570 18.895 47.900 ;
        RECT 18.610 47.425 18.780 47.570 ;
        RECT 18.115 47.255 18.780 47.425 ;
        RECT 19.065 47.400 19.235 48.200 ;
        RECT 19.415 48.225 19.745 48.700 ;
        RECT 19.915 48.395 20.085 48.875 ;
        RECT 20.255 48.225 20.585 48.700 ;
        RECT 20.755 48.395 20.925 48.875 ;
        RECT 21.095 48.225 21.425 48.700 ;
        RECT 21.595 48.395 21.765 48.875 ;
        RECT 21.935 48.225 22.265 48.700 ;
        RECT 22.435 48.395 22.605 48.875 ;
        RECT 22.775 48.225 23.105 48.700 ;
        RECT 23.275 48.395 23.445 48.875 ;
        RECT 23.615 48.700 23.865 48.705 ;
        RECT 23.615 48.225 23.945 48.700 ;
        RECT 24.115 48.395 24.285 48.875 ;
        RECT 24.535 48.700 24.705 48.705 ;
        RECT 24.455 48.225 24.785 48.700 ;
        RECT 24.955 48.395 25.125 48.875 ;
        RECT 25.375 48.700 25.545 48.705 ;
        RECT 25.295 48.225 25.625 48.700 ;
        RECT 25.795 48.395 25.965 48.875 ;
        RECT 26.135 48.225 26.465 48.700 ;
        RECT 26.635 48.395 26.805 48.875 ;
        RECT 26.975 48.225 27.305 48.700 ;
        RECT 27.475 48.395 27.645 48.875 ;
        RECT 27.815 48.225 28.145 48.700 ;
        RECT 28.315 48.395 28.485 48.875 ;
        RECT 28.655 48.225 28.985 48.700 ;
        RECT 29.155 48.395 29.325 48.875 ;
        RECT 29.495 48.225 29.825 48.700 ;
        RECT 29.995 48.395 30.165 48.875 ;
        RECT 19.415 48.055 20.925 48.225 ;
        RECT 21.095 48.055 23.445 48.225 ;
        RECT 23.615 48.055 30.275 48.225 ;
        RECT 31.365 48.150 31.655 48.875 ;
        RECT 20.755 47.885 20.925 48.055 ;
        RECT 23.270 47.885 23.445 48.055 ;
        RECT 19.410 47.685 20.585 47.885 ;
        RECT 20.755 47.685 23.065 47.885 ;
        RECT 23.270 47.685 29.830 47.885 ;
        RECT 20.755 47.515 20.925 47.685 ;
        RECT 23.270 47.515 23.445 47.685 ;
        RECT 30.000 47.515 30.275 48.055 ;
        RECT 31.825 48.125 33.035 48.875 ;
        RECT 33.210 48.325 33.465 48.615 ;
        RECT 33.635 48.495 33.965 48.875 ;
        RECT 33.210 48.155 33.960 48.325 ;
        RECT 31.825 47.585 32.345 48.125 ;
        RECT 16.640 46.995 17.390 47.165 ;
        RECT 16.635 46.325 16.965 46.825 ;
        RECT 17.135 46.495 17.390 46.995 ;
        RECT 18.115 46.495 18.285 47.255 ;
        RECT 18.465 46.325 18.795 47.085 ;
        RECT 18.965 46.495 19.235 47.400 ;
        RECT 19.415 47.345 20.925 47.515 ;
        RECT 21.095 47.345 23.445 47.515 ;
        RECT 23.615 47.345 30.275 47.515 ;
        RECT 19.415 46.495 19.745 47.345 ;
        RECT 19.915 46.325 20.085 47.175 ;
        RECT 20.255 46.495 20.585 47.345 ;
        RECT 20.755 46.325 20.925 47.175 ;
        RECT 21.095 46.495 21.425 47.345 ;
        RECT 21.595 46.325 21.765 47.125 ;
        RECT 21.935 46.495 22.265 47.345 ;
        RECT 22.435 46.325 22.605 47.125 ;
        RECT 22.775 46.495 23.105 47.345 ;
        RECT 23.275 46.325 23.445 47.125 ;
        RECT 23.615 46.495 23.945 47.345 ;
        RECT 24.115 46.325 24.285 47.125 ;
        RECT 24.455 46.495 24.785 47.345 ;
        RECT 24.955 46.325 25.125 47.125 ;
        RECT 25.295 46.495 25.625 47.345 ;
        RECT 25.795 46.325 25.965 47.125 ;
        RECT 26.135 46.495 26.465 47.345 ;
        RECT 26.635 46.325 26.805 47.125 ;
        RECT 26.975 46.495 27.305 47.345 ;
        RECT 27.475 46.325 27.645 47.125 ;
        RECT 27.815 46.495 28.145 47.345 ;
        RECT 28.315 46.325 28.485 47.125 ;
        RECT 28.655 46.495 28.985 47.345 ;
        RECT 29.155 46.325 29.325 47.125 ;
        RECT 29.495 46.495 29.825 47.345 ;
        RECT 29.995 46.325 30.165 47.125 ;
        RECT 31.365 46.325 31.655 47.490 ;
        RECT 32.515 47.415 33.035 47.955 ;
        RECT 31.825 46.325 33.035 47.415 ;
        RECT 33.210 47.335 33.560 47.985 ;
        RECT 33.730 47.165 33.960 48.155 ;
        RECT 33.210 46.995 33.960 47.165 ;
        RECT 33.210 46.495 33.465 46.995 ;
        RECT 33.635 46.325 33.965 46.825 ;
        RECT 34.135 46.495 34.305 48.615 ;
        RECT 34.665 48.515 34.995 48.875 ;
        RECT 35.165 48.485 35.660 48.655 ;
        RECT 35.865 48.485 36.720 48.655 ;
        RECT 34.535 47.295 34.995 48.345 ;
        RECT 34.475 46.510 34.800 47.295 ;
        RECT 35.165 47.125 35.335 48.485 ;
        RECT 35.505 47.575 35.855 48.195 ;
        RECT 36.025 47.975 36.380 48.195 ;
        RECT 36.025 47.385 36.195 47.975 ;
        RECT 36.550 47.775 36.720 48.485 ;
        RECT 37.595 48.415 37.925 48.875 ;
        RECT 38.135 48.515 38.485 48.685 ;
        RECT 36.925 47.945 37.715 48.195 ;
        RECT 38.135 48.125 38.395 48.515 ;
        RECT 38.705 48.425 39.655 48.705 ;
        RECT 39.825 48.435 40.015 48.875 ;
        RECT 40.185 48.495 41.255 48.665 ;
        RECT 37.885 47.775 38.055 47.955 ;
        RECT 35.165 46.955 35.560 47.125 ;
        RECT 35.730 46.995 36.195 47.385 ;
        RECT 36.365 47.605 38.055 47.775 ;
        RECT 35.390 46.825 35.560 46.955 ;
        RECT 36.365 46.825 36.535 47.605 ;
        RECT 38.225 47.435 38.395 48.125 ;
        RECT 36.895 47.265 38.395 47.435 ;
        RECT 38.585 47.465 38.795 48.255 ;
        RECT 38.965 47.635 39.315 48.255 ;
        RECT 39.485 47.645 39.655 48.425 ;
        RECT 40.185 48.265 40.355 48.495 ;
        RECT 39.825 48.095 40.355 48.265 ;
        RECT 39.825 47.815 40.045 48.095 ;
        RECT 40.525 47.925 40.765 48.325 ;
        RECT 39.485 47.475 39.890 47.645 ;
        RECT 40.225 47.555 40.765 47.925 ;
        RECT 40.935 48.140 41.255 48.495 ;
        RECT 41.500 48.415 41.805 48.875 ;
        RECT 41.975 48.165 42.230 48.695 ;
        RECT 40.935 47.965 41.260 48.140 ;
        RECT 40.935 47.665 41.850 47.965 ;
        RECT 41.110 47.635 41.850 47.665 ;
        RECT 38.585 47.305 39.260 47.465 ;
        RECT 39.720 47.385 39.890 47.475 ;
        RECT 38.585 47.295 39.550 47.305 ;
        RECT 38.225 47.125 38.395 47.265 ;
        RECT 34.970 46.325 35.220 46.785 ;
        RECT 35.390 46.495 35.640 46.825 ;
        RECT 35.855 46.495 36.535 46.825 ;
        RECT 36.705 46.925 37.780 47.095 ;
        RECT 38.225 46.955 38.785 47.125 ;
        RECT 39.090 47.005 39.550 47.295 ;
        RECT 39.720 47.215 40.940 47.385 ;
        RECT 36.705 46.585 36.875 46.925 ;
        RECT 37.110 46.325 37.440 46.755 ;
        RECT 37.610 46.585 37.780 46.925 ;
        RECT 38.075 46.325 38.445 46.785 ;
        RECT 38.615 46.495 38.785 46.955 ;
        RECT 39.720 46.835 39.890 47.215 ;
        RECT 41.110 47.045 41.280 47.635 ;
        RECT 42.020 47.515 42.230 48.165 ;
        RECT 42.465 48.055 42.675 48.875 ;
        RECT 42.845 48.075 43.175 48.705 ;
        RECT 39.020 46.495 39.890 46.835 ;
        RECT 40.480 46.875 41.280 47.045 ;
        RECT 40.060 46.325 40.310 46.785 ;
        RECT 40.480 46.585 40.650 46.875 ;
        RECT 40.830 46.325 41.160 46.705 ;
        RECT 41.500 46.325 41.805 47.465 ;
        RECT 41.975 46.635 42.230 47.515 ;
        RECT 42.845 47.475 43.095 48.075 ;
        RECT 43.345 48.055 43.575 48.875 ;
        RECT 43.785 48.105 47.295 48.875 ;
        RECT 43.265 47.635 43.595 47.885 ;
        RECT 43.785 47.585 45.435 48.105 ;
        RECT 48.425 48.055 48.655 48.875 ;
        RECT 48.825 48.075 49.155 48.705 ;
        RECT 42.465 46.325 42.675 47.465 ;
        RECT 42.845 46.495 43.175 47.475 ;
        RECT 43.345 46.325 43.575 47.465 ;
        RECT 45.605 47.415 47.295 47.935 ;
        RECT 48.405 47.635 48.735 47.885 ;
        RECT 48.905 47.475 49.155 48.075 ;
        RECT 49.325 48.055 49.535 48.875 ;
        RECT 49.765 48.330 55.110 48.875 ;
        RECT 51.350 47.500 51.690 48.330 ;
        RECT 55.285 48.105 56.955 48.875 ;
        RECT 57.125 48.150 57.415 48.875 ;
        RECT 57.585 48.105 59.255 48.875 ;
        RECT 43.785 46.325 47.295 47.415 ;
        RECT 48.425 46.325 48.655 47.465 ;
        RECT 48.825 46.495 49.155 47.475 ;
        RECT 49.325 46.325 49.535 47.465 ;
        RECT 53.170 46.760 53.520 48.010 ;
        RECT 55.285 47.585 56.035 48.105 ;
        RECT 56.205 47.415 56.955 47.935 ;
        RECT 57.585 47.585 58.335 48.105 ;
        RECT 59.430 48.035 59.690 48.875 ;
        RECT 59.865 48.130 60.120 48.705 ;
        RECT 60.290 48.495 60.620 48.875 ;
        RECT 60.835 48.325 61.005 48.705 ;
        RECT 60.290 48.155 61.005 48.325 ;
        RECT 61.355 48.325 61.525 48.705 ;
        RECT 61.740 48.495 62.070 48.875 ;
        RECT 61.355 48.155 62.070 48.325 ;
        RECT 49.765 46.325 55.110 46.760 ;
        RECT 55.285 46.325 56.955 47.415 ;
        RECT 57.125 46.325 57.415 47.490 ;
        RECT 58.505 47.415 59.255 47.935 ;
        RECT 57.585 46.325 59.255 47.415 ;
        RECT 59.430 46.325 59.690 47.475 ;
        RECT 59.865 47.400 60.035 48.130 ;
        RECT 60.290 47.965 60.460 48.155 ;
        RECT 60.205 47.635 60.460 47.965 ;
        RECT 60.290 47.425 60.460 47.635 ;
        RECT 60.740 47.605 61.095 47.975 ;
        RECT 61.265 47.605 61.620 47.975 ;
        RECT 61.900 47.965 62.070 48.155 ;
        RECT 62.240 48.130 62.495 48.705 ;
        RECT 61.900 47.635 62.155 47.965 ;
        RECT 61.900 47.425 62.070 47.635 ;
        RECT 59.865 46.495 60.120 47.400 ;
        RECT 60.290 47.255 61.005 47.425 ;
        RECT 60.290 46.325 60.620 47.085 ;
        RECT 60.835 46.495 61.005 47.255 ;
        RECT 61.355 47.255 62.070 47.425 ;
        RECT 62.325 47.400 62.495 48.130 ;
        RECT 62.670 48.035 62.930 48.875 ;
        RECT 63.105 48.330 68.450 48.875 ;
        RECT 64.690 47.500 65.030 48.330 ;
        RECT 68.625 48.105 72.135 48.875 ;
        RECT 72.775 48.385 73.105 48.875 ;
        RECT 73.275 48.280 73.895 48.705 ;
        RECT 61.355 46.495 61.525 47.255 ;
        RECT 61.740 46.325 62.070 47.085 ;
        RECT 62.240 46.495 62.495 47.400 ;
        RECT 62.670 46.325 62.930 47.475 ;
        RECT 66.510 46.760 66.860 48.010 ;
        RECT 68.625 47.585 70.275 48.105 ;
        RECT 70.445 47.415 72.135 47.935 ;
        RECT 72.765 47.635 73.105 48.215 ;
        RECT 73.275 47.945 73.635 48.280 ;
        RECT 74.355 48.185 74.685 48.875 ;
        RECT 75.730 48.095 76.230 48.705 ;
        RECT 73.275 47.665 74.695 47.945 ;
        RECT 63.105 46.325 68.450 46.760 ;
        RECT 68.625 46.325 72.135 47.415 ;
        RECT 72.775 46.325 73.105 47.465 ;
        RECT 73.275 46.495 73.635 47.665 ;
        RECT 73.835 46.325 74.165 47.495 ;
        RECT 74.365 46.495 74.695 47.665 ;
        RECT 75.525 47.635 75.875 47.885 ;
        RECT 74.895 46.325 75.225 47.495 ;
        RECT 76.060 47.465 76.230 48.095 ;
        RECT 76.860 48.225 77.190 48.705 ;
        RECT 77.360 48.415 77.585 48.875 ;
        RECT 77.755 48.225 78.085 48.705 ;
        RECT 76.860 48.055 78.085 48.225 ;
        RECT 78.275 48.075 78.525 48.875 ;
        RECT 78.695 48.075 79.035 48.705 ;
        RECT 78.805 48.025 79.035 48.075 ;
        RECT 76.400 47.685 76.730 47.885 ;
        RECT 76.900 47.685 77.230 47.885 ;
        RECT 77.400 47.685 77.820 47.885 ;
        RECT 77.995 47.715 78.690 47.885 ;
        RECT 77.995 47.465 78.165 47.715 ;
        RECT 78.860 47.465 79.035 48.025 ;
        RECT 79.205 48.105 82.715 48.875 ;
        RECT 82.885 48.150 83.175 48.875 ;
        RECT 83.345 48.105 85.935 48.875 ;
        RECT 86.110 48.325 86.365 48.615 ;
        RECT 86.535 48.495 86.865 48.875 ;
        RECT 86.110 48.155 86.860 48.325 ;
        RECT 79.205 47.585 80.855 48.105 ;
        RECT 75.730 47.295 78.165 47.465 ;
        RECT 75.730 46.495 76.060 47.295 ;
        RECT 76.230 46.325 76.560 47.125 ;
        RECT 76.860 46.495 77.190 47.295 ;
        RECT 77.835 46.325 78.085 47.125 ;
        RECT 78.355 46.325 78.525 47.465 ;
        RECT 78.695 46.495 79.035 47.465 ;
        RECT 81.025 47.415 82.715 47.935 ;
        RECT 83.345 47.585 84.555 48.105 ;
        RECT 79.205 46.325 82.715 47.415 ;
        RECT 82.885 46.325 83.175 47.490 ;
        RECT 84.725 47.415 85.935 47.935 ;
        RECT 83.345 46.325 85.935 47.415 ;
        RECT 86.110 47.335 86.460 47.985 ;
        RECT 86.630 47.165 86.860 48.155 ;
        RECT 86.110 46.995 86.860 47.165 ;
        RECT 86.110 46.495 86.365 46.995 ;
        RECT 86.535 46.325 86.865 46.825 ;
        RECT 87.035 46.495 87.205 48.615 ;
        RECT 87.565 48.515 87.895 48.875 ;
        RECT 88.065 48.485 88.560 48.655 ;
        RECT 88.765 48.485 89.620 48.655 ;
        RECT 87.435 47.295 87.895 48.345 ;
        RECT 87.375 46.510 87.700 47.295 ;
        RECT 88.065 47.125 88.235 48.485 ;
        RECT 88.405 47.575 88.755 48.195 ;
        RECT 88.925 47.975 89.280 48.195 ;
        RECT 88.925 47.385 89.095 47.975 ;
        RECT 89.450 47.775 89.620 48.485 ;
        RECT 90.495 48.415 90.825 48.875 ;
        RECT 91.035 48.515 91.385 48.685 ;
        RECT 89.825 47.945 90.615 48.195 ;
        RECT 91.035 48.125 91.295 48.515 ;
        RECT 91.605 48.425 92.555 48.705 ;
        RECT 92.725 48.435 92.915 48.875 ;
        RECT 93.085 48.495 94.155 48.665 ;
        RECT 90.785 47.775 90.955 47.955 ;
        RECT 88.065 46.955 88.460 47.125 ;
        RECT 88.630 46.995 89.095 47.385 ;
        RECT 89.265 47.605 90.955 47.775 ;
        RECT 88.290 46.825 88.460 46.955 ;
        RECT 89.265 46.825 89.435 47.605 ;
        RECT 91.125 47.435 91.295 48.125 ;
        RECT 89.795 47.265 91.295 47.435 ;
        RECT 91.485 47.465 91.695 48.255 ;
        RECT 91.865 47.635 92.215 48.255 ;
        RECT 92.385 47.645 92.555 48.425 ;
        RECT 93.085 48.265 93.255 48.495 ;
        RECT 92.725 48.095 93.255 48.265 ;
        RECT 92.725 47.815 92.945 48.095 ;
        RECT 93.425 47.925 93.665 48.325 ;
        RECT 92.385 47.475 92.790 47.645 ;
        RECT 93.125 47.555 93.665 47.925 ;
        RECT 93.835 48.140 94.155 48.495 ;
        RECT 94.400 48.415 94.705 48.875 ;
        RECT 94.875 48.165 95.130 48.695 ;
        RECT 93.835 47.965 94.160 48.140 ;
        RECT 93.835 47.665 94.750 47.965 ;
        RECT 94.010 47.635 94.750 47.665 ;
        RECT 91.485 47.305 92.160 47.465 ;
        RECT 92.620 47.385 92.790 47.475 ;
        RECT 91.485 47.295 92.450 47.305 ;
        RECT 91.125 47.125 91.295 47.265 ;
        RECT 87.870 46.325 88.120 46.785 ;
        RECT 88.290 46.495 88.540 46.825 ;
        RECT 88.755 46.495 89.435 46.825 ;
        RECT 89.605 46.925 90.680 47.095 ;
        RECT 91.125 46.955 91.685 47.125 ;
        RECT 91.990 47.005 92.450 47.295 ;
        RECT 92.620 47.215 93.840 47.385 ;
        RECT 89.605 46.585 89.775 46.925 ;
        RECT 90.010 46.325 90.340 46.755 ;
        RECT 90.510 46.585 90.680 46.925 ;
        RECT 90.975 46.325 91.345 46.785 ;
        RECT 91.515 46.495 91.685 46.955 ;
        RECT 92.620 46.835 92.790 47.215 ;
        RECT 94.010 47.045 94.180 47.635 ;
        RECT 94.920 47.515 95.130 48.165 ;
        RECT 95.315 48.225 95.645 48.700 ;
        RECT 95.815 48.395 95.985 48.875 ;
        RECT 96.155 48.225 96.485 48.700 ;
        RECT 96.655 48.395 96.825 48.875 ;
        RECT 96.995 48.225 97.325 48.700 ;
        RECT 97.495 48.395 97.665 48.875 ;
        RECT 97.835 48.225 98.165 48.700 ;
        RECT 98.335 48.395 98.505 48.875 ;
        RECT 98.675 48.225 99.005 48.700 ;
        RECT 99.175 48.395 99.345 48.875 ;
        RECT 99.515 48.700 99.765 48.705 ;
        RECT 99.515 48.225 99.845 48.700 ;
        RECT 100.015 48.395 100.185 48.875 ;
        RECT 100.435 48.700 100.605 48.705 ;
        RECT 100.355 48.225 100.685 48.700 ;
        RECT 100.855 48.395 101.025 48.875 ;
        RECT 101.275 48.700 101.445 48.705 ;
        RECT 101.195 48.225 101.525 48.700 ;
        RECT 101.695 48.395 101.865 48.875 ;
        RECT 102.035 48.225 102.365 48.700 ;
        RECT 102.535 48.395 102.705 48.875 ;
        RECT 102.875 48.225 103.205 48.700 ;
        RECT 103.375 48.395 103.545 48.875 ;
        RECT 103.715 48.225 104.045 48.700 ;
        RECT 104.215 48.395 104.385 48.875 ;
        RECT 104.555 48.225 104.885 48.700 ;
        RECT 105.055 48.395 105.225 48.875 ;
        RECT 105.395 48.225 105.725 48.700 ;
        RECT 105.895 48.395 106.065 48.875 ;
        RECT 95.315 48.055 96.825 48.225 ;
        RECT 96.995 48.055 99.345 48.225 ;
        RECT 99.515 48.055 106.175 48.225 ;
        RECT 96.655 47.885 96.825 48.055 ;
        RECT 99.170 47.885 99.345 48.055 ;
        RECT 95.310 47.685 96.485 47.885 ;
        RECT 96.655 47.685 98.965 47.885 ;
        RECT 99.170 47.685 105.730 47.885 ;
        RECT 96.655 47.515 96.825 47.685 ;
        RECT 99.170 47.515 99.345 47.685 ;
        RECT 105.900 47.515 106.175 48.055 ;
        RECT 106.345 48.105 108.015 48.875 ;
        RECT 108.645 48.150 108.935 48.875 ;
        RECT 109.105 48.105 111.695 48.875 ;
        RECT 112.325 48.125 113.535 48.875 ;
        RECT 106.345 47.585 107.095 48.105 ;
        RECT 91.920 46.495 92.790 46.835 ;
        RECT 93.380 46.875 94.180 47.045 ;
        RECT 92.960 46.325 93.210 46.785 ;
        RECT 93.380 46.585 93.550 46.875 ;
        RECT 93.730 46.325 94.060 46.705 ;
        RECT 94.400 46.325 94.705 47.465 ;
        RECT 94.875 46.635 95.130 47.515 ;
        RECT 95.315 47.345 96.825 47.515 ;
        RECT 96.995 47.345 99.345 47.515 ;
        RECT 99.515 47.345 106.175 47.515 ;
        RECT 107.265 47.415 108.015 47.935 ;
        RECT 109.105 47.585 110.315 48.105 ;
        RECT 95.315 46.495 95.645 47.345 ;
        RECT 95.815 46.325 95.985 47.175 ;
        RECT 96.155 46.495 96.485 47.345 ;
        RECT 96.655 46.325 96.825 47.175 ;
        RECT 96.995 46.495 97.325 47.345 ;
        RECT 97.495 46.325 97.665 47.125 ;
        RECT 97.835 46.495 98.165 47.345 ;
        RECT 98.335 46.325 98.505 47.125 ;
        RECT 98.675 46.495 99.005 47.345 ;
        RECT 99.175 46.325 99.345 47.125 ;
        RECT 99.515 46.495 99.845 47.345 ;
        RECT 100.015 46.325 100.185 47.125 ;
        RECT 100.355 46.495 100.685 47.345 ;
        RECT 100.855 46.325 101.025 47.125 ;
        RECT 101.195 46.495 101.525 47.345 ;
        RECT 101.695 46.325 101.865 47.125 ;
        RECT 102.035 46.495 102.365 47.345 ;
        RECT 102.535 46.325 102.705 47.125 ;
        RECT 102.875 46.495 103.205 47.345 ;
        RECT 103.375 46.325 103.545 47.125 ;
        RECT 103.715 46.495 104.045 47.345 ;
        RECT 104.215 46.325 104.385 47.125 ;
        RECT 104.555 46.495 104.885 47.345 ;
        RECT 105.055 46.325 105.225 47.125 ;
        RECT 105.395 46.495 105.725 47.345 ;
        RECT 105.895 46.325 106.065 47.125 ;
        RECT 106.345 46.325 108.015 47.415 ;
        RECT 108.645 46.325 108.935 47.490 ;
        RECT 110.485 47.415 111.695 47.935 ;
        RECT 109.105 46.325 111.695 47.415 ;
        RECT 112.325 47.415 112.845 47.955 ;
        RECT 113.015 47.585 113.535 48.125 ;
        RECT 112.325 46.325 113.535 47.415 ;
        RECT 5.520 46.155 113.620 46.325 ;
        RECT 5.605 45.065 6.815 46.155 ;
        RECT 6.985 45.720 12.330 46.155 ;
        RECT 5.605 44.355 6.125 44.895 ;
        RECT 6.295 44.525 6.815 45.065 ;
        RECT 5.605 43.605 6.815 44.355 ;
        RECT 8.570 44.150 8.910 44.980 ;
        RECT 10.390 44.470 10.740 45.720 ;
        RECT 12.505 45.065 16.015 46.155 ;
        RECT 12.505 44.375 14.155 44.895 ;
        RECT 14.325 44.545 16.015 45.065 ;
        RECT 17.165 45.015 17.375 46.155 ;
        RECT 17.545 45.005 17.875 45.985 ;
        RECT 18.045 45.015 18.275 46.155 ;
        RECT 6.985 43.605 12.330 44.150 ;
        RECT 12.505 43.605 16.015 44.375 ;
        RECT 17.165 43.605 17.375 44.425 ;
        RECT 17.545 44.405 17.795 45.005 ;
        RECT 18.485 44.990 18.775 46.155 ;
        RECT 19.005 45.015 19.215 46.155 ;
        RECT 19.385 45.005 19.715 45.985 ;
        RECT 19.885 45.015 20.115 46.155 ;
        RECT 20.325 45.080 20.595 45.985 ;
        RECT 20.765 45.395 21.095 46.155 ;
        RECT 21.275 45.225 21.445 45.985 ;
        RECT 21.710 45.485 21.965 45.985 ;
        RECT 22.135 45.655 22.465 46.155 ;
        RECT 21.710 45.315 22.460 45.485 ;
        RECT 17.965 44.595 18.295 44.845 ;
        RECT 17.545 43.775 17.875 44.405 ;
        RECT 18.045 43.605 18.275 44.425 ;
        RECT 18.485 43.605 18.775 44.330 ;
        RECT 19.005 43.605 19.215 44.425 ;
        RECT 19.385 44.405 19.635 45.005 ;
        RECT 19.805 44.595 20.135 44.845 ;
        RECT 19.385 43.775 19.715 44.405 ;
        RECT 19.885 43.605 20.115 44.425 ;
        RECT 20.325 44.280 20.495 45.080 ;
        RECT 20.780 45.055 21.445 45.225 ;
        RECT 20.780 44.910 20.950 45.055 ;
        RECT 20.665 44.580 20.950 44.910 ;
        RECT 20.780 44.325 20.950 44.580 ;
        RECT 21.185 44.505 21.515 44.875 ;
        RECT 21.710 44.495 22.060 45.145 ;
        RECT 22.230 44.325 22.460 45.315 ;
        RECT 20.325 43.775 20.585 44.280 ;
        RECT 20.780 44.155 21.445 44.325 ;
        RECT 20.765 43.605 21.095 43.985 ;
        RECT 21.275 43.775 21.445 44.155 ;
        RECT 21.710 44.155 22.460 44.325 ;
        RECT 21.710 43.865 21.965 44.155 ;
        RECT 22.135 43.605 22.465 43.985 ;
        RECT 22.635 43.865 22.805 45.985 ;
        RECT 22.975 45.185 23.300 45.970 ;
        RECT 23.470 45.695 23.720 46.155 ;
        RECT 23.890 45.655 24.140 45.985 ;
        RECT 24.355 45.655 25.035 45.985 ;
        RECT 23.890 45.525 24.060 45.655 ;
        RECT 23.665 45.355 24.060 45.525 ;
        RECT 23.035 44.135 23.495 45.185 ;
        RECT 23.665 43.995 23.835 45.355 ;
        RECT 24.230 45.095 24.695 45.485 ;
        RECT 24.005 44.285 24.355 44.905 ;
        RECT 24.525 44.505 24.695 45.095 ;
        RECT 24.865 44.875 25.035 45.655 ;
        RECT 25.205 45.555 25.375 45.895 ;
        RECT 25.610 45.725 25.940 46.155 ;
        RECT 26.110 45.555 26.280 45.895 ;
        RECT 26.575 45.695 26.945 46.155 ;
        RECT 25.205 45.385 26.280 45.555 ;
        RECT 27.115 45.525 27.285 45.985 ;
        RECT 27.520 45.645 28.390 45.985 ;
        RECT 28.560 45.695 28.810 46.155 ;
        RECT 26.725 45.355 27.285 45.525 ;
        RECT 26.725 45.215 26.895 45.355 ;
        RECT 25.395 45.045 26.895 45.215 ;
        RECT 27.590 45.185 28.050 45.475 ;
        RECT 24.865 44.705 26.555 44.875 ;
        RECT 24.525 44.285 24.880 44.505 ;
        RECT 25.050 43.995 25.220 44.705 ;
        RECT 25.425 44.285 26.215 44.535 ;
        RECT 26.385 44.525 26.555 44.705 ;
        RECT 26.725 44.355 26.895 45.045 ;
        RECT 23.165 43.605 23.495 43.965 ;
        RECT 23.665 43.825 24.160 43.995 ;
        RECT 24.365 43.825 25.220 43.995 ;
        RECT 26.095 43.605 26.425 44.065 ;
        RECT 26.635 43.965 26.895 44.355 ;
        RECT 27.085 45.175 28.050 45.185 ;
        RECT 28.220 45.265 28.390 45.645 ;
        RECT 28.980 45.605 29.150 45.895 ;
        RECT 29.330 45.775 29.660 46.155 ;
        RECT 28.980 45.435 29.780 45.605 ;
        RECT 27.085 45.015 27.760 45.175 ;
        RECT 28.220 45.095 29.440 45.265 ;
        RECT 27.085 44.225 27.295 45.015 ;
        RECT 28.220 45.005 28.390 45.095 ;
        RECT 27.465 44.225 27.815 44.845 ;
        RECT 27.985 44.835 28.390 45.005 ;
        RECT 27.985 44.055 28.155 44.835 ;
        RECT 28.325 44.385 28.545 44.665 ;
        RECT 28.725 44.555 29.265 44.925 ;
        RECT 29.610 44.845 29.780 45.435 ;
        RECT 30.000 45.015 30.305 46.155 ;
        RECT 30.475 44.965 30.730 45.845 ;
        RECT 30.965 45.015 31.175 46.155 ;
        RECT 29.610 44.815 30.350 44.845 ;
        RECT 28.325 44.215 28.855 44.385 ;
        RECT 26.635 43.795 26.985 43.965 ;
        RECT 27.205 43.775 28.155 44.055 ;
        RECT 28.325 43.605 28.515 44.045 ;
        RECT 28.685 43.985 28.855 44.215 ;
        RECT 29.025 44.155 29.265 44.555 ;
        RECT 29.435 44.515 30.350 44.815 ;
        RECT 29.435 44.340 29.760 44.515 ;
        RECT 29.435 43.985 29.755 44.340 ;
        RECT 30.520 44.315 30.730 44.965 ;
        RECT 31.345 45.005 31.675 45.985 ;
        RECT 31.845 45.015 32.075 46.155 ;
        RECT 32.285 45.720 37.630 46.155 ;
        RECT 28.685 43.815 29.755 43.985 ;
        RECT 30.000 43.605 30.305 44.065 ;
        RECT 30.475 43.785 30.730 44.315 ;
        RECT 30.965 43.605 31.175 44.425 ;
        RECT 31.345 44.405 31.595 45.005 ;
        RECT 31.765 44.595 32.095 44.845 ;
        RECT 31.345 43.775 31.675 44.405 ;
        RECT 31.845 43.605 32.075 44.425 ;
        RECT 33.870 44.150 34.210 44.980 ;
        RECT 35.690 44.470 36.040 45.720 ;
        RECT 38.265 45.185 38.525 46.155 ;
        RECT 32.285 43.605 37.630 44.150 ;
        RECT 38.265 43.895 38.505 44.845 ;
        RECT 38.695 44.810 39.025 45.985 ;
        RECT 39.195 45.185 39.475 46.155 ;
        RECT 39.645 45.065 43.155 46.155 ;
        RECT 38.695 44.280 39.475 44.810 ;
        RECT 39.645 44.375 41.295 44.895 ;
        RECT 41.465 44.545 43.155 45.065 ;
        RECT 44.245 44.990 44.535 46.155 ;
        RECT 44.855 45.005 45.185 46.155 ;
        RECT 45.355 45.135 45.525 45.985 ;
        RECT 45.695 45.355 46.025 46.155 ;
        RECT 46.195 45.135 46.365 45.985 ;
        RECT 46.545 45.355 46.785 46.155 ;
        RECT 46.955 45.175 47.285 45.985 ;
        RECT 45.355 44.965 46.365 45.135 ;
        RECT 46.570 45.005 47.285 45.175 ;
        RECT 48.130 45.185 48.460 45.985 ;
        RECT 48.630 45.355 48.960 46.155 ;
        RECT 49.260 45.185 49.590 45.985 ;
        RECT 50.235 45.355 50.485 46.155 ;
        RECT 48.130 45.015 50.565 45.185 ;
        RECT 50.755 45.015 50.925 46.155 ;
        RECT 51.095 45.015 51.435 45.985 ;
        RECT 51.605 45.065 55.115 46.155 ;
        RECT 55.285 45.065 56.495 46.155 ;
        RECT 45.355 44.455 45.850 44.965 ;
        RECT 46.570 44.765 46.740 45.005 ;
        RECT 46.240 44.595 46.740 44.765 ;
        RECT 46.910 44.595 47.290 44.835 ;
        RECT 47.925 44.595 48.275 44.845 ;
        RECT 45.355 44.425 45.855 44.455 ;
        RECT 46.570 44.425 46.740 44.595 ;
        RECT 38.695 43.775 39.020 44.280 ;
        RECT 39.190 43.605 39.475 44.110 ;
        RECT 39.645 43.605 43.155 44.375 ;
        RECT 44.245 43.605 44.535 44.330 ;
        RECT 44.855 43.605 45.185 44.405 ;
        RECT 45.355 44.255 46.365 44.425 ;
        RECT 46.570 44.255 47.205 44.425 ;
        RECT 48.460 44.385 48.630 45.015 ;
        RECT 48.800 44.595 49.130 44.795 ;
        RECT 49.300 44.595 49.630 44.795 ;
        RECT 49.800 44.595 50.220 44.795 ;
        RECT 50.395 44.765 50.565 45.015 ;
        RECT 50.395 44.595 51.090 44.765 ;
        RECT 45.355 43.775 45.525 44.255 ;
        RECT 45.695 43.605 46.025 44.085 ;
        RECT 46.195 43.775 46.365 44.255 ;
        RECT 46.615 43.605 46.855 44.085 ;
        RECT 47.035 43.775 47.205 44.255 ;
        RECT 48.130 43.775 48.630 44.385 ;
        RECT 49.260 44.255 50.485 44.425 ;
        RECT 51.260 44.405 51.435 45.015 ;
        RECT 49.260 43.775 49.590 44.255 ;
        RECT 49.760 43.605 49.985 44.065 ;
        RECT 50.155 43.775 50.485 44.255 ;
        RECT 50.675 43.605 50.925 44.405 ;
        RECT 51.095 43.775 51.435 44.405 ;
        RECT 51.605 44.375 53.255 44.895 ;
        RECT 53.425 44.545 55.115 45.065 ;
        RECT 51.605 43.605 55.115 44.375 ;
        RECT 55.285 44.355 55.805 44.895 ;
        RECT 55.975 44.525 56.495 45.065 ;
        RECT 56.670 45.005 56.930 46.155 ;
        RECT 57.105 45.080 57.360 45.985 ;
        RECT 57.530 45.395 57.860 46.155 ;
        RECT 58.075 45.225 58.245 45.985 ;
        RECT 55.285 43.605 56.495 44.355 ;
        RECT 56.670 43.605 56.930 44.445 ;
        RECT 57.105 44.350 57.275 45.080 ;
        RECT 57.530 45.055 58.245 45.225 ;
        RECT 58.595 45.225 58.765 45.985 ;
        RECT 58.980 45.395 59.310 46.155 ;
        RECT 58.595 45.055 59.310 45.225 ;
        RECT 59.480 45.080 59.735 45.985 ;
        RECT 57.530 44.845 57.700 45.055 ;
        RECT 57.445 44.515 57.700 44.845 ;
        RECT 57.105 43.775 57.360 44.350 ;
        RECT 57.530 44.325 57.700 44.515 ;
        RECT 57.980 44.505 58.335 44.875 ;
        RECT 58.505 44.505 58.860 44.875 ;
        RECT 59.140 44.845 59.310 45.055 ;
        RECT 59.140 44.515 59.395 44.845 ;
        RECT 59.140 44.325 59.310 44.515 ;
        RECT 59.565 44.350 59.735 45.080 ;
        RECT 59.910 45.005 60.170 46.155 ;
        RECT 60.350 45.005 60.610 46.155 ;
        RECT 60.785 45.080 61.040 45.985 ;
        RECT 61.210 45.395 61.540 46.155 ;
        RECT 61.755 45.225 61.925 45.985 ;
        RECT 57.530 44.155 58.245 44.325 ;
        RECT 57.530 43.605 57.860 43.985 ;
        RECT 58.075 43.775 58.245 44.155 ;
        RECT 58.595 44.155 59.310 44.325 ;
        RECT 58.595 43.775 58.765 44.155 ;
        RECT 58.980 43.605 59.310 43.985 ;
        RECT 59.480 43.775 59.735 44.350 ;
        RECT 59.910 43.605 60.170 44.445 ;
        RECT 60.350 43.605 60.610 44.445 ;
        RECT 60.785 44.350 60.955 45.080 ;
        RECT 61.210 45.055 61.925 45.225 ;
        RECT 62.275 45.225 62.445 45.985 ;
        RECT 62.660 45.395 62.990 46.155 ;
        RECT 62.275 45.055 62.990 45.225 ;
        RECT 63.160 45.080 63.415 45.985 ;
        RECT 61.210 44.845 61.380 45.055 ;
        RECT 61.125 44.515 61.380 44.845 ;
        RECT 60.785 43.775 61.040 44.350 ;
        RECT 61.210 44.325 61.380 44.515 ;
        RECT 61.660 44.505 62.015 44.875 ;
        RECT 62.185 44.505 62.540 44.875 ;
        RECT 62.820 44.845 62.990 45.055 ;
        RECT 62.820 44.515 63.075 44.845 ;
        RECT 62.820 44.325 62.990 44.515 ;
        RECT 63.245 44.350 63.415 45.080 ;
        RECT 63.590 45.005 63.850 46.155 ;
        RECT 64.115 45.225 64.285 45.985 ;
        RECT 64.500 45.395 64.830 46.155 ;
        RECT 64.115 45.055 64.830 45.225 ;
        RECT 65.000 45.080 65.255 45.985 ;
        RECT 64.025 44.505 64.380 44.875 ;
        RECT 64.660 44.845 64.830 45.055 ;
        RECT 64.660 44.515 64.915 44.845 ;
        RECT 61.210 44.155 61.925 44.325 ;
        RECT 61.210 43.605 61.540 43.985 ;
        RECT 61.755 43.775 61.925 44.155 ;
        RECT 62.275 44.155 62.990 44.325 ;
        RECT 62.275 43.775 62.445 44.155 ;
        RECT 62.660 43.605 62.990 43.985 ;
        RECT 63.160 43.775 63.415 44.350 ;
        RECT 63.590 43.605 63.850 44.445 ;
        RECT 64.660 44.325 64.830 44.515 ;
        RECT 65.085 44.350 65.255 45.080 ;
        RECT 65.430 45.005 65.690 46.155 ;
        RECT 65.865 45.065 69.375 46.155 ;
        RECT 64.115 44.155 64.830 44.325 ;
        RECT 64.115 43.775 64.285 44.155 ;
        RECT 64.500 43.605 64.830 43.985 ;
        RECT 65.000 43.775 65.255 44.350 ;
        RECT 65.430 43.605 65.690 44.445 ;
        RECT 65.865 44.375 67.515 44.895 ;
        RECT 67.685 44.545 69.375 45.065 ;
        RECT 70.005 44.990 70.295 46.155 ;
        RECT 70.465 45.065 72.135 46.155 ;
        RECT 72.775 45.345 73.070 46.155 ;
        RECT 70.465 44.375 71.215 44.895 ;
        RECT 71.385 44.545 72.135 45.065 ;
        RECT 73.250 44.845 73.495 45.985 ;
        RECT 73.670 45.345 73.930 46.155 ;
        RECT 74.530 46.150 80.805 46.155 ;
        RECT 74.110 44.845 74.360 45.980 ;
        RECT 74.530 45.355 74.790 46.150 ;
        RECT 74.960 45.255 75.220 45.980 ;
        RECT 75.390 45.425 75.650 46.150 ;
        RECT 75.820 45.255 76.080 45.980 ;
        RECT 76.250 45.425 76.510 46.150 ;
        RECT 76.680 45.255 76.940 45.980 ;
        RECT 77.110 45.425 77.370 46.150 ;
        RECT 77.540 45.255 77.800 45.980 ;
        RECT 77.970 45.425 78.215 46.150 ;
        RECT 78.385 45.255 78.645 45.980 ;
        RECT 78.830 45.425 79.075 46.150 ;
        RECT 79.245 45.255 79.505 45.980 ;
        RECT 79.690 45.425 79.935 46.150 ;
        RECT 80.105 45.255 80.365 45.980 ;
        RECT 80.550 45.425 80.805 46.150 ;
        RECT 74.960 45.240 80.365 45.255 ;
        RECT 80.975 45.240 81.265 45.980 ;
        RECT 81.435 45.410 81.705 46.155 ;
        RECT 74.960 45.015 81.705 45.240 ;
        RECT 65.865 43.605 69.375 44.375 ;
        RECT 70.005 43.605 70.295 44.330 ;
        RECT 70.465 43.605 72.135 44.375 ;
        RECT 72.765 44.285 73.080 44.845 ;
        RECT 73.250 44.595 80.370 44.845 ;
        RECT 72.765 43.605 73.070 44.115 ;
        RECT 73.250 43.785 73.500 44.595 ;
        RECT 73.670 43.605 73.930 44.130 ;
        RECT 74.110 43.785 74.360 44.595 ;
        RECT 80.540 44.425 81.705 45.015 ;
        RECT 74.960 44.255 81.705 44.425 ;
        RECT 81.965 45.015 82.305 45.985 ;
        RECT 82.475 45.015 82.645 46.155 ;
        RECT 82.915 45.355 83.165 46.155 ;
        RECT 83.810 45.185 84.140 45.985 ;
        RECT 84.440 45.355 84.770 46.155 ;
        RECT 84.940 45.185 85.270 45.985 ;
        RECT 82.835 45.015 85.270 45.185 ;
        RECT 85.645 45.015 85.985 45.985 ;
        RECT 86.155 45.015 86.325 46.155 ;
        RECT 86.595 45.355 86.845 46.155 ;
        RECT 87.490 45.185 87.820 45.985 ;
        RECT 88.120 45.355 88.450 46.155 ;
        RECT 88.620 45.185 88.950 45.985 ;
        RECT 86.515 45.015 88.950 45.185 ;
        RECT 89.325 45.015 89.665 45.985 ;
        RECT 89.835 45.015 90.005 46.155 ;
        RECT 90.275 45.355 90.525 46.155 ;
        RECT 91.170 45.185 91.500 45.985 ;
        RECT 91.800 45.355 92.130 46.155 ;
        RECT 92.300 45.185 92.630 45.985 ;
        RECT 90.195 45.015 92.630 45.185 ;
        RECT 93.005 45.065 95.595 46.155 ;
        RECT 81.965 44.405 82.140 45.015 ;
        RECT 82.835 44.765 83.005 45.015 ;
        RECT 82.310 44.595 83.005 44.765 ;
        RECT 83.180 44.595 83.600 44.795 ;
        RECT 83.770 44.595 84.100 44.795 ;
        RECT 84.270 44.595 84.600 44.795 ;
        RECT 74.530 43.605 74.790 44.165 ;
        RECT 74.960 43.800 75.220 44.255 ;
        RECT 75.390 43.605 75.650 44.085 ;
        RECT 75.820 43.800 76.080 44.255 ;
        RECT 76.250 43.605 76.510 44.085 ;
        RECT 76.680 43.800 76.940 44.255 ;
        RECT 77.110 43.605 77.355 44.085 ;
        RECT 77.525 43.800 77.800 44.255 ;
        RECT 77.970 43.605 78.215 44.085 ;
        RECT 78.385 43.800 78.645 44.255 ;
        RECT 78.825 43.605 79.075 44.085 ;
        RECT 79.245 43.800 79.505 44.255 ;
        RECT 79.685 43.605 79.935 44.085 ;
        RECT 80.105 43.800 80.365 44.255 ;
        RECT 80.545 43.605 80.805 44.085 ;
        RECT 80.975 43.800 81.235 44.255 ;
        RECT 81.405 43.605 81.705 44.085 ;
        RECT 81.965 43.775 82.305 44.405 ;
        RECT 82.475 43.605 82.725 44.405 ;
        RECT 82.915 44.255 84.140 44.425 ;
        RECT 82.915 43.775 83.245 44.255 ;
        RECT 83.415 43.605 83.640 44.065 ;
        RECT 83.810 43.775 84.140 44.255 ;
        RECT 84.770 44.385 84.940 45.015 ;
        RECT 85.125 44.595 85.475 44.845 ;
        RECT 85.645 44.405 85.820 45.015 ;
        RECT 86.515 44.765 86.685 45.015 ;
        RECT 85.990 44.595 86.685 44.765 ;
        RECT 86.860 44.595 87.280 44.795 ;
        RECT 87.450 44.595 87.780 44.795 ;
        RECT 87.950 44.595 88.280 44.795 ;
        RECT 84.770 43.775 85.270 44.385 ;
        RECT 85.645 43.775 85.985 44.405 ;
        RECT 86.155 43.605 86.405 44.405 ;
        RECT 86.595 44.255 87.820 44.425 ;
        RECT 86.595 43.775 86.925 44.255 ;
        RECT 87.095 43.605 87.320 44.065 ;
        RECT 87.490 43.775 87.820 44.255 ;
        RECT 88.450 44.385 88.620 45.015 ;
        RECT 88.805 44.595 89.155 44.845 ;
        RECT 89.325 44.405 89.500 45.015 ;
        RECT 90.195 44.765 90.365 45.015 ;
        RECT 89.670 44.595 90.365 44.765 ;
        RECT 90.540 44.595 90.960 44.795 ;
        RECT 91.130 44.595 91.460 44.795 ;
        RECT 91.630 44.595 91.960 44.795 ;
        RECT 88.450 43.775 88.950 44.385 ;
        RECT 89.325 43.775 89.665 44.405 ;
        RECT 89.835 43.605 90.085 44.405 ;
        RECT 90.275 44.255 91.500 44.425 ;
        RECT 90.275 43.775 90.605 44.255 ;
        RECT 90.775 43.605 91.000 44.065 ;
        RECT 91.170 43.775 91.500 44.255 ;
        RECT 92.130 44.385 92.300 45.015 ;
        RECT 92.485 44.595 92.835 44.845 ;
        RECT 92.130 43.775 92.630 44.385 ;
        RECT 93.005 44.375 94.215 44.895 ;
        RECT 94.385 44.545 95.595 45.065 ;
        RECT 95.765 44.990 96.055 46.155 ;
        RECT 96.235 45.345 96.530 46.155 ;
        RECT 96.710 44.845 96.955 45.985 ;
        RECT 97.130 45.345 97.390 46.155 ;
        RECT 97.990 46.150 104.265 46.155 ;
        RECT 97.570 44.845 97.820 45.980 ;
        RECT 97.990 45.355 98.250 46.150 ;
        RECT 98.420 45.255 98.680 45.980 ;
        RECT 98.850 45.425 99.110 46.150 ;
        RECT 99.280 45.255 99.540 45.980 ;
        RECT 99.710 45.425 99.970 46.150 ;
        RECT 100.140 45.255 100.400 45.980 ;
        RECT 100.570 45.425 100.830 46.150 ;
        RECT 101.000 45.255 101.260 45.980 ;
        RECT 101.430 45.425 101.675 46.150 ;
        RECT 101.845 45.255 102.105 45.980 ;
        RECT 102.290 45.425 102.535 46.150 ;
        RECT 102.705 45.255 102.965 45.980 ;
        RECT 103.150 45.425 103.395 46.150 ;
        RECT 103.565 45.255 103.825 45.980 ;
        RECT 104.010 45.425 104.265 46.150 ;
        RECT 98.420 45.240 103.825 45.255 ;
        RECT 104.435 45.240 104.725 45.980 ;
        RECT 104.895 45.410 105.165 46.155 ;
        RECT 105.425 45.720 110.770 46.155 ;
        RECT 98.420 45.015 105.165 45.240 ;
        RECT 93.005 43.605 95.595 44.375 ;
        RECT 95.765 43.605 96.055 44.330 ;
        RECT 96.225 44.285 96.540 44.845 ;
        RECT 96.710 44.595 103.830 44.845 ;
        RECT 96.225 43.605 96.530 44.115 ;
        RECT 96.710 43.785 96.960 44.595 ;
        RECT 97.130 43.605 97.390 44.130 ;
        RECT 97.570 43.785 97.820 44.595 ;
        RECT 104.000 44.425 105.165 45.015 ;
        RECT 98.420 44.255 105.165 44.425 ;
        RECT 97.990 43.605 98.250 44.165 ;
        RECT 98.420 43.800 98.680 44.255 ;
        RECT 98.850 43.605 99.110 44.085 ;
        RECT 99.280 43.800 99.540 44.255 ;
        RECT 99.710 43.605 99.970 44.085 ;
        RECT 100.140 43.800 100.400 44.255 ;
        RECT 100.570 43.605 100.815 44.085 ;
        RECT 100.985 43.800 101.260 44.255 ;
        RECT 101.430 43.605 101.675 44.085 ;
        RECT 101.845 43.800 102.105 44.255 ;
        RECT 102.285 43.605 102.535 44.085 ;
        RECT 102.705 43.800 102.965 44.255 ;
        RECT 103.145 43.605 103.395 44.085 ;
        RECT 103.565 43.800 103.825 44.255 ;
        RECT 104.005 43.605 104.265 44.085 ;
        RECT 104.435 43.800 104.695 44.255 ;
        RECT 107.010 44.150 107.350 44.980 ;
        RECT 108.830 44.470 109.180 45.720 ;
        RECT 110.945 45.065 112.155 46.155 ;
        RECT 110.945 44.355 111.465 44.895 ;
        RECT 111.635 44.525 112.155 45.065 ;
        RECT 112.325 45.065 113.535 46.155 ;
        RECT 112.325 44.525 112.845 45.065 ;
        RECT 113.015 44.355 113.535 44.895 ;
        RECT 104.865 43.605 105.165 44.085 ;
        RECT 105.425 43.605 110.770 44.150 ;
        RECT 110.945 43.605 112.155 44.355 ;
        RECT 112.325 43.605 113.535 44.355 ;
        RECT 5.520 43.435 113.620 43.605 ;
        RECT 5.605 42.685 6.815 43.435 ;
        RECT 6.985 42.890 12.330 43.435 ;
        RECT 5.605 42.145 6.125 42.685 ;
        RECT 6.295 41.975 6.815 42.515 ;
        RECT 8.570 42.060 8.910 42.890 ;
        RECT 12.505 42.665 16.015 43.435 ;
        RECT 5.605 40.885 6.815 41.975 ;
        RECT 10.390 41.320 10.740 42.570 ;
        RECT 12.505 42.145 14.155 42.665 ;
        RECT 17.310 42.655 17.810 43.265 ;
        RECT 14.325 41.975 16.015 42.495 ;
        RECT 17.105 42.195 17.455 42.445 ;
        RECT 17.640 42.025 17.810 42.655 ;
        RECT 18.440 42.785 18.770 43.265 ;
        RECT 18.940 42.975 19.165 43.435 ;
        RECT 19.335 42.785 19.665 43.265 ;
        RECT 18.440 42.615 19.665 42.785 ;
        RECT 19.855 42.635 20.105 43.435 ;
        RECT 20.275 42.635 20.615 43.265 ;
        RECT 20.990 42.655 21.490 43.265 ;
        RECT 17.980 42.245 18.310 42.445 ;
        RECT 18.480 42.245 18.810 42.445 ;
        RECT 18.980 42.245 19.400 42.445 ;
        RECT 19.575 42.275 20.270 42.445 ;
        RECT 19.575 42.025 19.745 42.275 ;
        RECT 20.440 42.025 20.615 42.635 ;
        RECT 20.785 42.195 21.135 42.445 ;
        RECT 21.320 42.025 21.490 42.655 ;
        RECT 22.120 42.785 22.450 43.265 ;
        RECT 22.620 42.975 22.845 43.435 ;
        RECT 23.015 42.785 23.345 43.265 ;
        RECT 22.120 42.615 23.345 42.785 ;
        RECT 23.535 42.635 23.785 43.435 ;
        RECT 23.955 42.635 24.295 43.265 ;
        RECT 21.660 42.245 21.990 42.445 ;
        RECT 22.160 42.245 22.490 42.445 ;
        RECT 22.660 42.245 23.080 42.445 ;
        RECT 23.255 42.275 23.950 42.445 ;
        RECT 23.255 42.025 23.425 42.275 ;
        RECT 24.120 42.025 24.295 42.635 ;
        RECT 24.465 42.665 26.135 43.435 ;
        RECT 24.465 42.145 25.215 42.665 ;
        RECT 26.510 42.655 27.010 43.265 ;
        RECT 6.985 40.885 12.330 41.320 ;
        RECT 12.505 40.885 16.015 41.975 ;
        RECT 17.310 41.855 19.745 42.025 ;
        RECT 17.310 41.055 17.640 41.855 ;
        RECT 17.810 40.885 18.140 41.685 ;
        RECT 18.440 41.055 18.770 41.855 ;
        RECT 19.415 40.885 19.665 41.685 ;
        RECT 19.935 40.885 20.105 42.025 ;
        RECT 20.275 41.055 20.615 42.025 ;
        RECT 20.990 41.855 23.425 42.025 ;
        RECT 20.990 41.055 21.320 41.855 ;
        RECT 21.490 40.885 21.820 41.685 ;
        RECT 22.120 41.055 22.450 41.855 ;
        RECT 23.095 40.885 23.345 41.685 ;
        RECT 23.615 40.885 23.785 42.025 ;
        RECT 23.955 41.055 24.295 42.025 ;
        RECT 25.385 41.975 26.135 42.495 ;
        RECT 26.305 42.195 26.655 42.445 ;
        RECT 26.840 42.025 27.010 42.655 ;
        RECT 27.640 42.785 27.970 43.265 ;
        RECT 28.140 42.975 28.365 43.435 ;
        RECT 28.535 42.785 28.865 43.265 ;
        RECT 27.640 42.615 28.865 42.785 ;
        RECT 29.055 42.635 29.305 43.435 ;
        RECT 29.475 42.635 29.815 43.265 ;
        RECT 27.180 42.245 27.510 42.445 ;
        RECT 27.680 42.245 28.010 42.445 ;
        RECT 28.180 42.245 28.600 42.445 ;
        RECT 28.775 42.275 29.470 42.445 ;
        RECT 28.775 42.025 28.945 42.275 ;
        RECT 29.640 42.025 29.815 42.635 ;
        RECT 29.985 42.685 31.195 43.435 ;
        RECT 31.365 42.710 31.655 43.435 ;
        RECT 29.985 42.145 30.505 42.685 ;
        RECT 31.825 42.635 32.165 43.265 ;
        RECT 32.335 42.635 32.585 43.435 ;
        RECT 32.775 42.785 33.105 43.265 ;
        RECT 33.275 42.975 33.500 43.435 ;
        RECT 33.670 42.785 34.000 43.265 ;
        RECT 24.465 40.885 26.135 41.975 ;
        RECT 26.510 41.855 28.945 42.025 ;
        RECT 26.510 41.055 26.840 41.855 ;
        RECT 27.010 40.885 27.340 41.685 ;
        RECT 27.640 41.055 27.970 41.855 ;
        RECT 28.615 40.885 28.865 41.685 ;
        RECT 29.135 40.885 29.305 42.025 ;
        RECT 29.475 41.055 29.815 42.025 ;
        RECT 30.675 41.975 31.195 42.515 ;
        RECT 29.985 40.885 31.195 41.975 ;
        RECT 31.365 40.885 31.655 42.050 ;
        RECT 31.825 42.025 32.000 42.635 ;
        RECT 32.775 42.615 34.000 42.785 ;
        RECT 34.630 42.655 35.130 43.265 ;
        RECT 32.170 42.275 32.865 42.445 ;
        RECT 32.695 42.025 32.865 42.275 ;
        RECT 33.040 42.245 33.460 42.445 ;
        RECT 33.630 42.245 33.960 42.445 ;
        RECT 34.130 42.245 34.460 42.445 ;
        RECT 34.630 42.025 34.800 42.655 ;
        RECT 35.545 42.615 35.775 43.435 ;
        RECT 35.945 42.635 36.275 43.265 ;
        RECT 34.985 42.195 35.335 42.445 ;
        RECT 35.525 42.195 35.855 42.445 ;
        RECT 36.025 42.035 36.275 42.635 ;
        RECT 36.445 42.615 36.655 43.435 ;
        RECT 36.885 42.685 38.095 43.435 ;
        RECT 38.355 42.955 38.655 43.435 ;
        RECT 38.825 42.785 39.085 43.240 ;
        RECT 39.255 42.955 39.515 43.435 ;
        RECT 39.695 42.785 39.955 43.240 ;
        RECT 40.125 42.955 40.375 43.435 ;
        RECT 40.555 42.785 40.815 43.240 ;
        RECT 40.985 42.955 41.235 43.435 ;
        RECT 41.415 42.785 41.675 43.240 ;
        RECT 41.845 42.955 42.090 43.435 ;
        RECT 42.260 42.785 42.535 43.240 ;
        RECT 42.705 42.955 42.950 43.435 ;
        RECT 43.120 42.785 43.380 43.240 ;
        RECT 43.550 42.955 43.810 43.435 ;
        RECT 43.980 42.785 44.240 43.240 ;
        RECT 44.410 42.955 44.670 43.435 ;
        RECT 44.840 42.785 45.100 43.240 ;
        RECT 45.270 42.875 45.530 43.435 ;
        RECT 38.355 42.755 45.100 42.785 ;
        RECT 36.885 42.145 37.405 42.685 ;
        RECT 38.325 42.615 45.100 42.755 ;
        RECT 38.325 42.585 39.520 42.615 ;
        RECT 31.825 41.055 32.165 42.025 ;
        RECT 32.335 40.885 32.505 42.025 ;
        RECT 32.695 41.855 35.130 42.025 ;
        RECT 32.775 40.885 33.025 41.685 ;
        RECT 33.670 41.055 34.000 41.855 ;
        RECT 34.300 40.885 34.630 41.685 ;
        RECT 34.800 41.055 35.130 41.855 ;
        RECT 35.545 40.885 35.775 42.025 ;
        RECT 35.945 41.055 36.275 42.035 ;
        RECT 36.445 40.885 36.655 42.025 ;
        RECT 37.575 41.975 38.095 42.515 ;
        RECT 36.885 40.885 38.095 41.975 ;
        RECT 38.355 42.025 39.520 42.585 ;
        RECT 45.700 42.445 45.950 43.255 ;
        RECT 46.130 42.910 46.390 43.435 ;
        RECT 46.560 42.445 46.810 43.255 ;
        RECT 46.990 42.925 47.295 43.435 ;
        RECT 39.690 42.195 46.810 42.445 ;
        RECT 46.980 42.195 47.295 42.755 ;
        RECT 48.590 42.655 49.090 43.265 ;
        RECT 48.385 42.195 48.735 42.445 ;
        RECT 38.355 41.800 45.100 42.025 ;
        RECT 38.355 40.885 38.625 41.630 ;
        RECT 38.795 41.060 39.085 41.800 ;
        RECT 39.695 41.785 45.100 41.800 ;
        RECT 39.255 40.890 39.510 41.615 ;
        RECT 39.695 41.060 39.955 41.785 ;
        RECT 40.125 40.890 40.370 41.615 ;
        RECT 40.555 41.060 40.815 41.785 ;
        RECT 40.985 40.890 41.230 41.615 ;
        RECT 41.415 41.060 41.675 41.785 ;
        RECT 41.845 40.890 42.090 41.615 ;
        RECT 42.260 41.060 42.520 41.785 ;
        RECT 42.690 40.890 42.950 41.615 ;
        RECT 43.120 41.060 43.380 41.785 ;
        RECT 43.550 40.890 43.810 41.615 ;
        RECT 43.980 41.060 44.240 41.785 ;
        RECT 44.410 40.890 44.670 41.615 ;
        RECT 44.840 41.060 45.100 41.785 ;
        RECT 45.270 40.890 45.530 41.685 ;
        RECT 45.700 41.060 45.950 42.195 ;
        RECT 39.255 40.885 45.530 40.890 ;
        RECT 46.130 40.885 46.390 41.695 ;
        RECT 46.565 41.055 46.810 42.195 ;
        RECT 48.920 42.025 49.090 42.655 ;
        RECT 49.720 42.785 50.050 43.265 ;
        RECT 50.220 42.975 50.445 43.435 ;
        RECT 50.615 42.785 50.945 43.265 ;
        RECT 49.720 42.615 50.945 42.785 ;
        RECT 51.135 42.635 51.385 43.435 ;
        RECT 51.555 42.635 51.895 43.265 ;
        RECT 52.270 42.655 52.770 43.265 ;
        RECT 49.260 42.245 49.590 42.445 ;
        RECT 49.760 42.245 50.090 42.445 ;
        RECT 50.260 42.245 50.680 42.445 ;
        RECT 50.855 42.275 51.550 42.445 ;
        RECT 50.855 42.025 51.025 42.275 ;
        RECT 51.720 42.025 51.895 42.635 ;
        RECT 52.065 42.195 52.415 42.445 ;
        RECT 52.600 42.025 52.770 42.655 ;
        RECT 53.400 42.785 53.730 43.265 ;
        RECT 53.900 42.975 54.125 43.435 ;
        RECT 54.295 42.785 54.625 43.265 ;
        RECT 53.400 42.615 54.625 42.785 ;
        RECT 54.815 42.635 55.065 43.435 ;
        RECT 55.235 42.635 55.575 43.265 ;
        RECT 52.940 42.245 53.270 42.445 ;
        RECT 53.440 42.245 53.770 42.445 ;
        RECT 53.940 42.245 54.360 42.445 ;
        RECT 54.535 42.275 55.230 42.445 ;
        RECT 54.535 42.025 54.705 42.275 ;
        RECT 55.400 42.025 55.575 42.635 ;
        RECT 55.745 42.685 56.955 43.435 ;
        RECT 57.125 42.710 57.415 43.435 ;
        RECT 55.745 42.145 56.265 42.685 ;
        RECT 57.585 42.675 58.295 43.265 ;
        RECT 58.805 42.905 59.135 43.265 ;
        RECT 59.335 43.075 59.665 43.435 ;
        RECT 59.835 42.905 60.165 43.265 ;
        RECT 58.805 42.695 60.165 42.905 ;
        RECT 60.345 42.685 61.555 43.435 ;
        RECT 61.725 42.935 62.025 43.265 ;
        RECT 62.195 42.955 62.470 43.435 ;
        RECT 48.590 41.855 51.025 42.025 ;
        RECT 46.990 40.885 47.285 41.695 ;
        RECT 48.590 41.055 48.920 41.855 ;
        RECT 49.090 40.885 49.420 41.685 ;
        RECT 49.720 41.055 50.050 41.855 ;
        RECT 50.695 40.885 50.945 41.685 ;
        RECT 51.215 40.885 51.385 42.025 ;
        RECT 51.555 41.055 51.895 42.025 ;
        RECT 52.270 41.855 54.705 42.025 ;
        RECT 52.270 41.055 52.600 41.855 ;
        RECT 52.770 40.885 53.100 41.685 ;
        RECT 53.400 41.055 53.730 41.855 ;
        RECT 54.375 40.885 54.625 41.685 ;
        RECT 54.895 40.885 55.065 42.025 ;
        RECT 55.235 41.055 55.575 42.025 ;
        RECT 56.435 41.975 56.955 42.515 ;
        RECT 55.745 40.885 56.955 41.975 ;
        RECT 57.125 40.885 57.415 42.050 ;
        RECT 57.585 41.705 57.790 42.675 ;
        RECT 57.960 41.905 58.290 42.445 ;
        RECT 58.465 42.195 58.960 42.525 ;
        RECT 59.280 42.195 59.655 42.525 ;
        RECT 59.865 42.195 60.175 42.525 ;
        RECT 58.465 41.905 58.790 42.195 ;
        RECT 58.985 41.705 59.315 41.925 ;
        RECT 57.585 41.475 59.315 41.705 ;
        RECT 57.585 41.055 58.285 41.475 ;
        RECT 58.485 40.885 58.815 41.245 ;
        RECT 58.985 41.075 59.315 41.475 ;
        RECT 59.485 41.270 59.655 42.195 ;
        RECT 60.345 42.145 60.865 42.685 ;
        RECT 61.035 41.975 61.555 42.515 ;
        RECT 59.835 40.885 60.165 41.945 ;
        RECT 60.345 40.885 61.555 41.975 ;
        RECT 61.725 42.025 61.895 42.935 ;
        RECT 62.650 42.785 62.945 43.175 ;
        RECT 63.115 42.955 63.370 43.435 ;
        RECT 63.545 42.785 63.805 43.175 ;
        RECT 63.975 42.955 64.255 43.435 ;
        RECT 64.950 42.885 65.205 43.175 ;
        RECT 65.375 43.055 65.705 43.435 ;
        RECT 62.065 42.195 62.415 42.765 ;
        RECT 62.650 42.615 64.300 42.785 ;
        RECT 64.950 42.715 65.700 42.885 ;
        RECT 62.585 42.275 63.725 42.445 ;
        RECT 62.585 42.025 62.755 42.275 ;
        RECT 63.895 42.105 64.300 42.615 ;
        RECT 61.725 41.855 62.755 42.025 ;
        RECT 63.545 41.935 64.300 42.105 ;
        RECT 61.725 41.055 62.035 41.855 ;
        RECT 63.545 41.685 63.805 41.935 ;
        RECT 64.950 41.895 65.300 42.545 ;
        RECT 62.205 40.885 62.515 41.685 ;
        RECT 62.685 41.515 63.805 41.685 ;
        RECT 62.685 41.055 62.945 41.515 ;
        RECT 63.115 40.885 63.370 41.345 ;
        RECT 63.545 41.055 63.805 41.515 ;
        RECT 63.975 40.885 64.260 41.755 ;
        RECT 65.470 41.725 65.700 42.715 ;
        RECT 64.950 41.555 65.700 41.725 ;
        RECT 64.950 41.055 65.205 41.555 ;
        RECT 65.375 40.885 65.705 41.385 ;
        RECT 65.875 41.055 66.045 43.175 ;
        RECT 66.405 43.075 66.735 43.435 ;
        RECT 66.905 43.045 67.400 43.215 ;
        RECT 67.605 43.045 68.460 43.215 ;
        RECT 66.275 41.855 66.735 42.905 ;
        RECT 66.215 41.070 66.540 41.855 ;
        RECT 66.905 41.685 67.075 43.045 ;
        RECT 67.245 42.135 67.595 42.755 ;
        RECT 67.765 42.535 68.120 42.755 ;
        RECT 67.765 41.945 67.935 42.535 ;
        RECT 68.290 42.335 68.460 43.045 ;
        RECT 69.335 42.975 69.665 43.435 ;
        RECT 69.875 43.075 70.225 43.245 ;
        RECT 68.665 42.505 69.455 42.755 ;
        RECT 69.875 42.685 70.135 43.075 ;
        RECT 70.445 42.985 71.395 43.265 ;
        RECT 71.565 42.995 71.755 43.435 ;
        RECT 71.925 43.055 72.995 43.225 ;
        RECT 69.625 42.335 69.795 42.515 ;
        RECT 66.905 41.515 67.300 41.685 ;
        RECT 67.470 41.555 67.935 41.945 ;
        RECT 68.105 42.165 69.795 42.335 ;
        RECT 67.130 41.385 67.300 41.515 ;
        RECT 68.105 41.385 68.275 42.165 ;
        RECT 69.965 41.995 70.135 42.685 ;
        RECT 68.635 41.825 70.135 41.995 ;
        RECT 70.325 42.025 70.535 42.815 ;
        RECT 70.705 42.195 71.055 42.815 ;
        RECT 71.225 42.205 71.395 42.985 ;
        RECT 71.925 42.825 72.095 43.055 ;
        RECT 71.565 42.655 72.095 42.825 ;
        RECT 71.565 42.375 71.785 42.655 ;
        RECT 72.265 42.485 72.505 42.885 ;
        RECT 71.225 42.035 71.630 42.205 ;
        RECT 71.965 42.115 72.505 42.485 ;
        RECT 72.675 42.700 72.995 43.055 ;
        RECT 73.240 42.975 73.545 43.435 ;
        RECT 73.715 42.725 73.970 43.255 ;
        RECT 72.675 42.525 73.000 42.700 ;
        RECT 72.675 42.225 73.590 42.525 ;
        RECT 72.850 42.195 73.590 42.225 ;
        RECT 70.325 41.865 71.000 42.025 ;
        RECT 71.460 41.945 71.630 42.035 ;
        RECT 70.325 41.855 71.290 41.865 ;
        RECT 69.965 41.685 70.135 41.825 ;
        RECT 66.710 40.885 66.960 41.345 ;
        RECT 67.130 41.055 67.380 41.385 ;
        RECT 67.595 41.055 68.275 41.385 ;
        RECT 68.445 41.485 69.520 41.655 ;
        RECT 69.965 41.515 70.525 41.685 ;
        RECT 70.830 41.565 71.290 41.855 ;
        RECT 71.460 41.775 72.680 41.945 ;
        RECT 68.445 41.145 68.615 41.485 ;
        RECT 68.850 40.885 69.180 41.315 ;
        RECT 69.350 41.145 69.520 41.485 ;
        RECT 69.815 40.885 70.185 41.345 ;
        RECT 70.355 41.055 70.525 41.515 ;
        RECT 71.460 41.395 71.630 41.775 ;
        RECT 72.850 41.605 73.020 42.195 ;
        RECT 73.760 42.075 73.970 42.725 ;
        RECT 70.760 41.055 71.630 41.395 ;
        RECT 72.220 41.435 73.020 41.605 ;
        RECT 71.800 40.885 72.050 41.345 ;
        RECT 72.220 41.145 72.390 41.435 ;
        RECT 72.570 40.885 72.900 41.265 ;
        RECT 73.240 40.885 73.545 42.025 ;
        RECT 73.715 41.195 73.970 42.075 ;
        RECT 74.150 42.695 74.405 43.265 ;
        RECT 74.575 43.035 74.905 43.435 ;
        RECT 75.330 42.900 75.860 43.265 ;
        RECT 75.330 42.865 75.505 42.900 ;
        RECT 74.575 42.695 75.505 42.865 ;
        RECT 74.150 42.025 74.320 42.695 ;
        RECT 74.575 42.525 74.745 42.695 ;
        RECT 74.490 42.195 74.745 42.525 ;
        RECT 74.970 42.195 75.165 42.525 ;
        RECT 74.150 41.055 74.485 42.025 ;
        RECT 74.655 40.885 74.825 42.025 ;
        RECT 74.995 41.225 75.165 42.195 ;
        RECT 75.335 41.565 75.505 42.695 ;
        RECT 75.675 41.905 75.845 42.705 ;
        RECT 76.050 42.415 76.325 43.265 ;
        RECT 76.045 42.245 76.325 42.415 ;
        RECT 76.050 42.105 76.325 42.245 ;
        RECT 76.495 41.905 76.685 43.265 ;
        RECT 76.865 42.900 77.375 43.435 ;
        RECT 77.595 42.625 77.840 43.230 ;
        RECT 78.285 42.635 78.625 43.265 ;
        RECT 78.795 42.635 79.045 43.435 ;
        RECT 79.235 42.785 79.565 43.265 ;
        RECT 79.735 42.975 79.960 43.435 ;
        RECT 80.130 42.785 80.460 43.265 ;
        RECT 76.885 42.455 78.115 42.625 ;
        RECT 75.675 41.735 76.685 41.905 ;
        RECT 76.855 41.890 77.605 42.080 ;
        RECT 75.335 41.395 76.460 41.565 ;
        RECT 76.855 41.225 77.025 41.890 ;
        RECT 77.775 41.645 78.115 42.455 ;
        RECT 74.995 41.055 77.025 41.225 ;
        RECT 77.195 40.885 77.365 41.645 ;
        RECT 77.600 41.235 78.115 41.645 ;
        RECT 78.285 42.025 78.460 42.635 ;
        RECT 79.235 42.615 80.460 42.785 ;
        RECT 81.090 42.655 81.590 43.265 ;
        RECT 82.885 42.710 83.175 43.435 ;
        RECT 83.350 42.885 83.605 43.175 ;
        RECT 83.775 43.055 84.105 43.435 ;
        RECT 83.350 42.715 84.100 42.885 ;
        RECT 78.630 42.275 79.325 42.445 ;
        RECT 79.155 42.025 79.325 42.275 ;
        RECT 79.500 42.245 79.920 42.445 ;
        RECT 80.090 42.245 80.420 42.445 ;
        RECT 80.590 42.245 80.920 42.445 ;
        RECT 81.090 42.025 81.260 42.655 ;
        RECT 81.445 42.195 81.795 42.445 ;
        RECT 78.285 41.055 78.625 42.025 ;
        RECT 78.795 40.885 78.965 42.025 ;
        RECT 79.155 41.855 81.590 42.025 ;
        RECT 79.235 40.885 79.485 41.685 ;
        RECT 80.130 41.055 80.460 41.855 ;
        RECT 80.760 40.885 81.090 41.685 ;
        RECT 81.260 41.055 81.590 41.855 ;
        RECT 82.885 40.885 83.175 42.050 ;
        RECT 83.350 41.895 83.700 42.545 ;
        RECT 83.870 41.725 84.100 42.715 ;
        RECT 83.350 41.555 84.100 41.725 ;
        RECT 83.350 41.055 83.605 41.555 ;
        RECT 83.775 40.885 84.105 41.385 ;
        RECT 84.275 41.055 84.445 43.175 ;
        RECT 84.805 43.075 85.135 43.435 ;
        RECT 85.305 43.045 85.800 43.215 ;
        RECT 86.005 43.045 86.860 43.215 ;
        RECT 84.675 41.855 85.135 42.905 ;
        RECT 84.615 41.070 84.940 41.855 ;
        RECT 85.305 41.685 85.475 43.045 ;
        RECT 85.645 42.135 85.995 42.755 ;
        RECT 86.165 42.535 86.520 42.755 ;
        RECT 86.165 41.945 86.335 42.535 ;
        RECT 86.690 42.335 86.860 43.045 ;
        RECT 87.735 42.975 88.065 43.435 ;
        RECT 88.275 43.075 88.625 43.245 ;
        RECT 87.065 42.505 87.855 42.755 ;
        RECT 88.275 42.685 88.535 43.075 ;
        RECT 88.845 42.985 89.795 43.265 ;
        RECT 89.965 42.995 90.155 43.435 ;
        RECT 90.325 43.055 91.395 43.225 ;
        RECT 88.025 42.335 88.195 42.515 ;
        RECT 85.305 41.515 85.700 41.685 ;
        RECT 85.870 41.555 86.335 41.945 ;
        RECT 86.505 42.165 88.195 42.335 ;
        RECT 85.530 41.385 85.700 41.515 ;
        RECT 86.505 41.385 86.675 42.165 ;
        RECT 88.365 41.995 88.535 42.685 ;
        RECT 87.035 41.825 88.535 41.995 ;
        RECT 88.725 42.025 88.935 42.815 ;
        RECT 89.105 42.195 89.455 42.815 ;
        RECT 89.625 42.205 89.795 42.985 ;
        RECT 90.325 42.825 90.495 43.055 ;
        RECT 89.965 42.655 90.495 42.825 ;
        RECT 89.965 42.375 90.185 42.655 ;
        RECT 90.665 42.485 90.905 42.885 ;
        RECT 89.625 42.035 90.030 42.205 ;
        RECT 90.365 42.115 90.905 42.485 ;
        RECT 91.075 42.700 91.395 43.055 ;
        RECT 91.640 42.975 91.945 43.435 ;
        RECT 92.115 42.725 92.370 43.255 ;
        RECT 91.075 42.525 91.400 42.700 ;
        RECT 91.075 42.225 91.990 42.525 ;
        RECT 91.250 42.195 91.990 42.225 ;
        RECT 88.725 41.865 89.400 42.025 ;
        RECT 89.860 41.945 90.030 42.035 ;
        RECT 88.725 41.855 89.690 41.865 ;
        RECT 88.365 41.685 88.535 41.825 ;
        RECT 85.110 40.885 85.360 41.345 ;
        RECT 85.530 41.055 85.780 41.385 ;
        RECT 85.995 41.055 86.675 41.385 ;
        RECT 86.845 41.485 87.920 41.655 ;
        RECT 88.365 41.515 88.925 41.685 ;
        RECT 89.230 41.565 89.690 41.855 ;
        RECT 89.860 41.775 91.080 41.945 ;
        RECT 86.845 41.145 87.015 41.485 ;
        RECT 87.250 40.885 87.580 41.315 ;
        RECT 87.750 41.145 87.920 41.485 ;
        RECT 88.215 40.885 88.585 41.345 ;
        RECT 88.755 41.055 88.925 41.515 ;
        RECT 89.860 41.395 90.030 41.775 ;
        RECT 91.250 41.605 91.420 42.195 ;
        RECT 92.160 42.075 92.370 42.725 ;
        RECT 89.160 41.055 90.030 41.395 ;
        RECT 90.620 41.435 91.420 41.605 ;
        RECT 90.200 40.885 90.450 41.345 ;
        RECT 90.620 41.145 90.790 41.435 ;
        RECT 90.970 40.885 91.300 41.265 ;
        RECT 91.640 40.885 91.945 42.025 ;
        RECT 92.115 41.195 92.370 42.075 ;
        RECT 92.545 42.635 92.885 43.265 ;
        RECT 93.055 42.635 93.305 43.435 ;
        RECT 93.495 42.785 93.825 43.265 ;
        RECT 93.995 42.975 94.220 43.435 ;
        RECT 94.390 42.785 94.720 43.265 ;
        RECT 92.545 42.025 92.720 42.635 ;
        RECT 93.495 42.615 94.720 42.785 ;
        RECT 95.350 42.655 95.850 43.265 ;
        RECT 96.230 42.885 96.485 43.175 ;
        RECT 96.655 43.055 96.985 43.435 ;
        RECT 96.230 42.715 96.980 42.885 ;
        RECT 92.890 42.275 93.585 42.445 ;
        RECT 93.415 42.025 93.585 42.275 ;
        RECT 93.760 42.245 94.180 42.445 ;
        RECT 94.350 42.245 94.680 42.445 ;
        RECT 94.850 42.245 95.180 42.445 ;
        RECT 95.350 42.025 95.520 42.655 ;
        RECT 95.705 42.195 96.055 42.445 ;
        RECT 92.545 41.055 92.885 42.025 ;
        RECT 93.055 40.885 93.225 42.025 ;
        RECT 93.415 41.855 95.850 42.025 ;
        RECT 96.230 41.895 96.580 42.545 ;
        RECT 93.495 40.885 93.745 41.685 ;
        RECT 94.390 41.055 94.720 41.855 ;
        RECT 95.020 40.885 95.350 41.685 ;
        RECT 95.520 41.055 95.850 41.855 ;
        RECT 96.750 41.725 96.980 42.715 ;
        RECT 96.230 41.555 96.980 41.725 ;
        RECT 96.230 41.055 96.485 41.555 ;
        RECT 96.655 40.885 96.985 41.385 ;
        RECT 97.155 41.055 97.325 43.175 ;
        RECT 97.685 43.075 98.015 43.435 ;
        RECT 98.185 43.045 98.680 43.215 ;
        RECT 98.885 43.045 99.740 43.215 ;
        RECT 97.555 41.855 98.015 42.905 ;
        RECT 97.495 41.070 97.820 41.855 ;
        RECT 98.185 41.685 98.355 43.045 ;
        RECT 98.525 42.135 98.875 42.755 ;
        RECT 99.045 42.535 99.400 42.755 ;
        RECT 99.045 41.945 99.215 42.535 ;
        RECT 99.570 42.335 99.740 43.045 ;
        RECT 100.615 42.975 100.945 43.435 ;
        RECT 101.155 43.075 101.505 43.245 ;
        RECT 99.945 42.505 100.735 42.755 ;
        RECT 101.155 42.685 101.415 43.075 ;
        RECT 101.725 42.985 102.675 43.265 ;
        RECT 102.845 42.995 103.035 43.435 ;
        RECT 103.205 43.055 104.275 43.225 ;
        RECT 100.905 42.335 101.075 42.515 ;
        RECT 98.185 41.515 98.580 41.685 ;
        RECT 98.750 41.555 99.215 41.945 ;
        RECT 99.385 42.165 101.075 42.335 ;
        RECT 98.410 41.385 98.580 41.515 ;
        RECT 99.385 41.385 99.555 42.165 ;
        RECT 101.245 41.995 101.415 42.685 ;
        RECT 99.915 41.825 101.415 41.995 ;
        RECT 101.605 42.025 101.815 42.815 ;
        RECT 101.985 42.195 102.335 42.815 ;
        RECT 102.505 42.205 102.675 42.985 ;
        RECT 103.205 42.825 103.375 43.055 ;
        RECT 102.845 42.655 103.375 42.825 ;
        RECT 102.845 42.375 103.065 42.655 ;
        RECT 103.545 42.485 103.785 42.885 ;
        RECT 102.505 42.035 102.910 42.205 ;
        RECT 103.245 42.115 103.785 42.485 ;
        RECT 103.955 42.700 104.275 43.055 ;
        RECT 104.520 42.975 104.825 43.435 ;
        RECT 104.995 42.725 105.250 43.255 ;
        RECT 103.955 42.525 104.280 42.700 ;
        RECT 103.955 42.225 104.870 42.525 ;
        RECT 104.130 42.195 104.870 42.225 ;
        RECT 101.605 41.865 102.280 42.025 ;
        RECT 102.740 41.945 102.910 42.035 ;
        RECT 101.605 41.855 102.570 41.865 ;
        RECT 101.245 41.685 101.415 41.825 ;
        RECT 97.990 40.885 98.240 41.345 ;
        RECT 98.410 41.055 98.660 41.385 ;
        RECT 98.875 41.055 99.555 41.385 ;
        RECT 99.725 41.485 100.800 41.655 ;
        RECT 101.245 41.515 101.805 41.685 ;
        RECT 102.110 41.565 102.570 41.855 ;
        RECT 102.740 41.775 103.960 41.945 ;
        RECT 99.725 41.145 99.895 41.485 ;
        RECT 100.130 40.885 100.460 41.315 ;
        RECT 100.630 41.145 100.800 41.485 ;
        RECT 101.095 40.885 101.465 41.345 ;
        RECT 101.635 41.055 101.805 41.515 ;
        RECT 102.740 41.395 102.910 41.775 ;
        RECT 104.130 41.605 104.300 42.195 ;
        RECT 105.040 42.075 105.250 42.725 ;
        RECT 105.465 42.615 105.695 43.435 ;
        RECT 105.865 42.635 106.195 43.265 ;
        RECT 105.445 42.195 105.775 42.445 ;
        RECT 102.040 41.055 102.910 41.395 ;
        RECT 103.500 41.435 104.300 41.605 ;
        RECT 103.080 40.885 103.330 41.345 ;
        RECT 103.500 41.145 103.670 41.435 ;
        RECT 103.850 40.885 104.180 41.265 ;
        RECT 104.520 40.885 104.825 42.025 ;
        RECT 104.995 41.195 105.250 42.075 ;
        RECT 105.945 42.035 106.195 42.635 ;
        RECT 106.365 42.615 106.575 43.435 ;
        RECT 106.805 42.665 108.475 43.435 ;
        RECT 108.645 42.710 108.935 43.435 ;
        RECT 109.105 42.665 111.695 43.435 ;
        RECT 112.325 42.685 113.535 43.435 ;
        RECT 106.805 42.145 107.555 42.665 ;
        RECT 105.465 40.885 105.695 42.025 ;
        RECT 105.865 41.055 106.195 42.035 ;
        RECT 106.365 40.885 106.575 42.025 ;
        RECT 107.725 41.975 108.475 42.495 ;
        RECT 109.105 42.145 110.315 42.665 ;
        RECT 106.805 40.885 108.475 41.975 ;
        RECT 108.645 40.885 108.935 42.050 ;
        RECT 110.485 41.975 111.695 42.495 ;
        RECT 109.105 40.885 111.695 41.975 ;
        RECT 112.325 41.975 112.845 42.515 ;
        RECT 113.015 42.145 113.535 42.685 ;
        RECT 112.325 40.885 113.535 41.975 ;
        RECT 5.520 40.715 113.620 40.885 ;
        RECT 5.605 39.625 6.815 40.715 ;
        RECT 6.985 39.625 10.495 40.715 ;
        RECT 5.605 38.915 6.125 39.455 ;
        RECT 6.295 39.085 6.815 39.625 ;
        RECT 6.985 38.935 8.635 39.455 ;
        RECT 8.805 39.105 10.495 39.625 ;
        RECT 11.585 39.640 11.855 40.545 ;
        RECT 12.025 39.955 12.355 40.715 ;
        RECT 12.535 39.785 12.705 40.545 ;
        RECT 5.605 38.165 6.815 38.915 ;
        RECT 6.985 38.165 10.495 38.935 ;
        RECT 11.585 38.840 11.755 39.640 ;
        RECT 12.040 39.615 12.705 39.785 ;
        RECT 12.965 39.640 13.235 40.545 ;
        RECT 13.405 39.955 13.735 40.715 ;
        RECT 13.915 39.785 14.085 40.545 ;
        RECT 12.040 39.470 12.210 39.615 ;
        RECT 11.925 39.140 12.210 39.470 ;
        RECT 12.040 38.885 12.210 39.140 ;
        RECT 12.445 39.065 12.775 39.435 ;
        RECT 11.585 38.335 11.845 38.840 ;
        RECT 12.040 38.715 12.705 38.885 ;
        RECT 12.025 38.165 12.355 38.545 ;
        RECT 12.535 38.335 12.705 38.715 ;
        RECT 12.965 38.840 13.135 39.640 ;
        RECT 13.420 39.615 14.085 39.785 ;
        RECT 13.420 39.470 13.590 39.615 ;
        RECT 14.405 39.575 14.615 40.715 ;
        RECT 13.305 39.140 13.590 39.470 ;
        RECT 14.785 39.565 15.115 40.545 ;
        RECT 15.285 39.575 15.515 40.715 ;
        RECT 15.785 39.575 15.995 40.715 ;
        RECT 16.165 39.565 16.495 40.545 ;
        RECT 16.665 39.575 16.895 40.715 ;
        RECT 17.105 39.625 18.315 40.715 ;
        RECT 13.420 38.885 13.590 39.140 ;
        RECT 13.825 39.065 14.155 39.435 ;
        RECT 12.965 38.335 13.225 38.840 ;
        RECT 13.420 38.715 14.085 38.885 ;
        RECT 13.405 38.165 13.735 38.545 ;
        RECT 13.915 38.335 14.085 38.715 ;
        RECT 14.405 38.165 14.615 38.985 ;
        RECT 14.785 38.965 15.035 39.565 ;
        RECT 15.205 39.155 15.535 39.405 ;
        RECT 14.785 38.335 15.115 38.965 ;
        RECT 15.285 38.165 15.515 38.985 ;
        RECT 15.785 38.165 15.995 38.985 ;
        RECT 16.165 38.965 16.415 39.565 ;
        RECT 16.585 39.155 16.915 39.405 ;
        RECT 16.165 38.335 16.495 38.965 ;
        RECT 16.665 38.165 16.895 38.985 ;
        RECT 17.105 38.915 17.625 39.455 ;
        RECT 17.795 39.085 18.315 39.625 ;
        RECT 18.485 39.550 18.775 40.715 ;
        RECT 18.945 39.625 22.455 40.715 ;
        RECT 18.945 38.935 20.595 39.455 ;
        RECT 20.765 39.105 22.455 39.625 ;
        RECT 22.830 39.745 23.160 40.545 ;
        RECT 23.330 39.915 23.660 40.715 ;
        RECT 23.960 39.745 24.290 40.545 ;
        RECT 24.935 39.915 25.185 40.715 ;
        RECT 22.830 39.575 25.265 39.745 ;
        RECT 25.455 39.575 25.625 40.715 ;
        RECT 25.795 39.575 26.135 40.545 ;
        RECT 22.625 39.155 22.975 39.405 ;
        RECT 23.160 38.945 23.330 39.575 ;
        RECT 23.500 39.155 23.830 39.355 ;
        RECT 24.000 39.155 24.330 39.355 ;
        RECT 24.500 39.155 24.920 39.355 ;
        RECT 25.095 39.325 25.265 39.575 ;
        RECT 25.095 39.155 25.790 39.325 ;
        RECT 17.105 38.165 18.315 38.915 ;
        RECT 18.485 38.165 18.775 38.890 ;
        RECT 18.945 38.165 22.455 38.935 ;
        RECT 22.830 38.335 23.330 38.945 ;
        RECT 23.960 38.815 25.185 38.985 ;
        RECT 25.960 38.965 26.135 39.575 ;
        RECT 23.960 38.335 24.290 38.815 ;
        RECT 24.460 38.165 24.685 38.625 ;
        RECT 24.855 38.335 25.185 38.815 ;
        RECT 25.375 38.165 25.625 38.965 ;
        RECT 25.795 38.335 26.135 38.965 ;
        RECT 26.305 39.575 26.645 40.545 ;
        RECT 26.815 39.575 26.985 40.715 ;
        RECT 27.255 39.915 27.505 40.715 ;
        RECT 28.150 39.745 28.480 40.545 ;
        RECT 28.780 39.915 29.110 40.715 ;
        RECT 29.280 39.745 29.610 40.545 ;
        RECT 30.450 40.045 30.705 40.545 ;
        RECT 30.875 40.215 31.205 40.715 ;
        RECT 30.450 39.875 31.200 40.045 ;
        RECT 27.175 39.575 29.610 39.745 ;
        RECT 26.305 38.965 26.480 39.575 ;
        RECT 27.175 39.325 27.345 39.575 ;
        RECT 26.650 39.155 27.345 39.325 ;
        RECT 27.520 39.155 27.940 39.355 ;
        RECT 28.110 39.155 28.440 39.355 ;
        RECT 28.610 39.155 28.940 39.355 ;
        RECT 26.305 38.335 26.645 38.965 ;
        RECT 26.815 38.165 27.065 38.965 ;
        RECT 27.255 38.815 28.480 38.985 ;
        RECT 27.255 38.335 27.585 38.815 ;
        RECT 27.755 38.165 27.980 38.625 ;
        RECT 28.150 38.335 28.480 38.815 ;
        RECT 29.110 38.945 29.280 39.575 ;
        RECT 29.465 39.155 29.815 39.405 ;
        RECT 30.450 39.055 30.800 39.705 ;
        RECT 29.110 38.335 29.610 38.945 ;
        RECT 30.970 38.885 31.200 39.875 ;
        RECT 30.450 38.715 31.200 38.885 ;
        RECT 30.450 38.425 30.705 38.715 ;
        RECT 30.875 38.165 31.205 38.545 ;
        RECT 31.375 38.425 31.545 40.545 ;
        RECT 31.715 39.745 32.040 40.530 ;
        RECT 32.210 40.255 32.460 40.715 ;
        RECT 32.630 40.215 32.880 40.545 ;
        RECT 33.095 40.215 33.775 40.545 ;
        RECT 32.630 40.085 32.800 40.215 ;
        RECT 32.405 39.915 32.800 40.085 ;
        RECT 31.775 38.695 32.235 39.745 ;
        RECT 32.405 38.555 32.575 39.915 ;
        RECT 32.970 39.655 33.435 40.045 ;
        RECT 32.745 38.845 33.095 39.465 ;
        RECT 33.265 39.065 33.435 39.655 ;
        RECT 33.605 39.435 33.775 40.215 ;
        RECT 33.945 40.115 34.115 40.455 ;
        RECT 34.350 40.285 34.680 40.715 ;
        RECT 34.850 40.115 35.020 40.455 ;
        RECT 35.315 40.255 35.685 40.715 ;
        RECT 33.945 39.945 35.020 40.115 ;
        RECT 35.855 40.085 36.025 40.545 ;
        RECT 36.260 40.205 37.130 40.545 ;
        RECT 37.300 40.255 37.550 40.715 ;
        RECT 35.465 39.915 36.025 40.085 ;
        RECT 35.465 39.775 35.635 39.915 ;
        RECT 34.135 39.605 35.635 39.775 ;
        RECT 36.330 39.745 36.790 40.035 ;
        RECT 33.605 39.265 35.295 39.435 ;
        RECT 33.265 38.845 33.620 39.065 ;
        RECT 33.790 38.555 33.960 39.265 ;
        RECT 34.165 38.845 34.955 39.095 ;
        RECT 35.125 39.085 35.295 39.265 ;
        RECT 35.465 38.915 35.635 39.605 ;
        RECT 31.905 38.165 32.235 38.525 ;
        RECT 32.405 38.385 32.900 38.555 ;
        RECT 33.105 38.385 33.960 38.555 ;
        RECT 34.835 38.165 35.165 38.625 ;
        RECT 35.375 38.525 35.635 38.915 ;
        RECT 35.825 39.735 36.790 39.745 ;
        RECT 36.960 39.825 37.130 40.205 ;
        RECT 37.720 40.165 37.890 40.455 ;
        RECT 38.070 40.335 38.400 40.715 ;
        RECT 37.720 39.995 38.520 40.165 ;
        RECT 35.825 39.575 36.500 39.735 ;
        RECT 36.960 39.655 38.180 39.825 ;
        RECT 35.825 38.785 36.035 39.575 ;
        RECT 36.960 39.565 37.130 39.655 ;
        RECT 36.205 38.785 36.555 39.405 ;
        RECT 36.725 39.395 37.130 39.565 ;
        RECT 36.725 38.615 36.895 39.395 ;
        RECT 37.065 38.945 37.285 39.225 ;
        RECT 37.465 39.115 38.005 39.485 ;
        RECT 38.350 39.405 38.520 39.995 ;
        RECT 38.740 39.575 39.045 40.715 ;
        RECT 39.215 39.525 39.470 40.405 ;
        RECT 38.350 39.375 39.090 39.405 ;
        RECT 37.065 38.775 37.595 38.945 ;
        RECT 35.375 38.355 35.725 38.525 ;
        RECT 35.945 38.335 36.895 38.615 ;
        RECT 37.065 38.165 37.255 38.605 ;
        RECT 37.425 38.545 37.595 38.775 ;
        RECT 37.765 38.715 38.005 39.115 ;
        RECT 38.175 39.075 39.090 39.375 ;
        RECT 38.175 38.900 38.500 39.075 ;
        RECT 38.175 38.545 38.495 38.900 ;
        RECT 39.260 38.875 39.470 39.525 ;
        RECT 37.425 38.375 38.495 38.545 ;
        RECT 38.740 38.165 39.045 38.625 ;
        RECT 39.215 38.345 39.470 38.875 ;
        RECT 40.565 39.640 40.835 40.545 ;
        RECT 41.005 39.955 41.335 40.715 ;
        RECT 41.515 39.785 41.685 40.545 ;
        RECT 40.565 38.840 40.735 39.640 ;
        RECT 41.020 39.615 41.685 39.785 ;
        RECT 41.945 39.625 43.615 40.715 ;
        RECT 41.020 39.470 41.190 39.615 ;
        RECT 40.905 39.140 41.190 39.470 ;
        RECT 41.020 38.885 41.190 39.140 ;
        RECT 41.425 39.065 41.755 39.435 ;
        RECT 41.945 38.935 42.695 39.455 ;
        RECT 42.865 39.105 43.615 39.625 ;
        RECT 44.245 39.550 44.535 40.715 ;
        RECT 44.710 39.575 45.045 40.545 ;
        RECT 45.215 39.575 45.385 40.715 ;
        RECT 45.555 40.375 47.585 40.545 ;
        RECT 40.565 38.335 40.825 38.840 ;
        RECT 41.020 38.715 41.685 38.885 ;
        RECT 41.005 38.165 41.335 38.545 ;
        RECT 41.515 38.335 41.685 38.715 ;
        RECT 41.945 38.165 43.615 38.935 ;
        RECT 44.710 38.905 44.880 39.575 ;
        RECT 45.555 39.405 45.725 40.375 ;
        RECT 45.050 39.075 45.305 39.405 ;
        RECT 45.530 39.075 45.725 39.405 ;
        RECT 45.895 40.035 47.020 40.205 ;
        RECT 45.135 38.905 45.305 39.075 ;
        RECT 45.895 38.905 46.065 40.035 ;
        RECT 44.245 38.165 44.535 38.890 ;
        RECT 44.710 38.335 44.965 38.905 ;
        RECT 45.135 38.735 46.065 38.905 ;
        RECT 46.235 39.695 47.245 39.865 ;
        RECT 46.235 38.895 46.405 39.695 ;
        RECT 46.610 39.355 46.885 39.495 ;
        RECT 46.605 39.185 46.885 39.355 ;
        RECT 45.890 38.700 46.065 38.735 ;
        RECT 45.135 38.165 45.465 38.565 ;
        RECT 45.890 38.335 46.420 38.700 ;
        RECT 46.610 38.335 46.885 39.185 ;
        RECT 47.055 38.335 47.245 39.695 ;
        RECT 47.415 39.710 47.585 40.375 ;
        RECT 47.755 39.955 47.925 40.715 ;
        RECT 48.160 39.955 48.675 40.365 ;
        RECT 47.415 39.520 48.165 39.710 ;
        RECT 48.335 39.145 48.675 39.955 ;
        RECT 49.050 39.745 49.380 40.545 ;
        RECT 49.550 39.915 49.880 40.715 ;
        RECT 50.180 39.745 50.510 40.545 ;
        RECT 51.155 39.915 51.405 40.715 ;
        RECT 49.050 39.575 51.485 39.745 ;
        RECT 51.675 39.575 51.845 40.715 ;
        RECT 52.015 39.575 52.355 40.545 ;
        RECT 52.580 39.845 52.865 40.715 ;
        RECT 53.035 40.085 53.295 40.545 ;
        RECT 53.470 40.255 53.725 40.715 ;
        RECT 53.895 40.085 54.155 40.545 ;
        RECT 53.035 39.915 54.155 40.085 ;
        RECT 54.325 39.915 54.635 40.715 ;
        RECT 53.035 39.665 53.295 39.915 ;
        RECT 54.805 39.745 55.115 40.545 ;
        RECT 48.845 39.155 49.195 39.405 ;
        RECT 47.445 38.975 48.675 39.145 ;
        RECT 47.425 38.165 47.935 38.700 ;
        RECT 48.155 38.370 48.400 38.975 ;
        RECT 49.380 38.945 49.550 39.575 ;
        RECT 49.720 39.155 50.050 39.355 ;
        RECT 50.220 39.155 50.550 39.355 ;
        RECT 50.720 39.155 51.140 39.355 ;
        RECT 51.315 39.325 51.485 39.575 ;
        RECT 51.315 39.155 52.010 39.325 ;
        RECT 49.050 38.335 49.550 38.945 ;
        RECT 50.180 38.815 51.405 38.985 ;
        RECT 52.180 38.965 52.355 39.575 ;
        RECT 50.180 38.335 50.510 38.815 ;
        RECT 50.680 38.165 50.905 38.625 ;
        RECT 51.075 38.335 51.405 38.815 ;
        RECT 51.595 38.165 51.845 38.965 ;
        RECT 52.015 38.335 52.355 38.965 ;
        RECT 52.540 39.495 53.295 39.665 ;
        RECT 54.085 39.575 55.115 39.745 ;
        RECT 55.285 39.625 57.875 40.715 ;
        RECT 58.755 40.265 59.085 40.715 ;
        RECT 52.540 38.985 52.945 39.495 ;
        RECT 54.085 39.325 54.255 39.575 ;
        RECT 53.115 39.155 54.255 39.325 ;
        RECT 52.540 38.815 54.190 38.985 ;
        RECT 54.425 38.835 54.775 39.405 ;
        RECT 52.585 38.165 52.865 38.645 ;
        RECT 53.035 38.425 53.295 38.815 ;
        RECT 53.470 38.165 53.725 38.645 ;
        RECT 53.895 38.425 54.190 38.815 ;
        RECT 54.945 38.665 55.115 39.575 ;
        RECT 54.370 38.165 54.645 38.645 ;
        RECT 54.815 38.335 55.115 38.665 ;
        RECT 55.285 38.935 56.495 39.455 ;
        RECT 56.665 39.105 57.875 39.625 ;
        RECT 58.045 39.875 60.655 40.085 ;
        RECT 55.285 38.165 57.875 38.935 ;
        RECT 58.045 38.905 58.215 39.875 ;
        RECT 58.385 39.075 58.735 39.695 ;
        RECT 58.905 39.075 59.225 39.695 ;
        RECT 59.395 39.075 59.725 39.695 ;
        RECT 59.895 39.075 60.195 39.695 ;
        RECT 60.435 39.075 60.655 39.875 ;
        RECT 60.835 38.905 61.095 40.530 ;
        RECT 62.335 39.565 62.665 40.715 ;
        RECT 62.835 39.695 63.005 40.545 ;
        RECT 63.175 39.915 63.505 40.715 ;
        RECT 63.675 39.695 63.845 40.545 ;
        RECT 64.025 39.915 64.265 40.715 ;
        RECT 64.435 39.735 64.765 40.545 ;
        RECT 62.835 39.525 63.845 39.695 ;
        RECT 64.050 39.565 64.765 39.735 ;
        RECT 65.005 39.575 65.215 40.715 ;
        RECT 65.385 39.565 65.715 40.545 ;
        RECT 65.885 39.575 66.115 40.715 ;
        RECT 66.415 39.785 66.585 40.545 ;
        RECT 66.765 39.955 67.095 40.715 ;
        RECT 66.415 39.615 67.080 39.785 ;
        RECT 67.265 39.640 67.535 40.545 ;
        RECT 62.835 39.015 63.330 39.525 ;
        RECT 64.050 39.325 64.220 39.565 ;
        RECT 63.720 39.155 64.220 39.325 ;
        RECT 64.390 39.155 64.770 39.395 ;
        RECT 62.835 38.985 63.335 39.015 ;
        RECT 64.050 38.985 64.220 39.155 ;
        RECT 58.045 38.735 58.520 38.905 ;
        RECT 58.350 38.485 58.520 38.735 ;
        RECT 58.755 38.165 59.085 38.905 ;
        RECT 59.255 38.735 61.095 38.905 ;
        RECT 59.255 38.390 59.455 38.735 ;
        RECT 59.625 38.165 59.955 38.565 ;
        RECT 60.125 38.380 60.325 38.735 ;
        RECT 60.495 38.165 60.825 38.560 ;
        RECT 62.335 38.165 62.665 38.965 ;
        RECT 62.835 38.815 63.845 38.985 ;
        RECT 64.050 38.815 64.685 38.985 ;
        RECT 62.835 38.335 63.005 38.815 ;
        RECT 63.175 38.165 63.505 38.645 ;
        RECT 63.675 38.335 63.845 38.815 ;
        RECT 64.095 38.165 64.335 38.645 ;
        RECT 64.515 38.335 64.685 38.815 ;
        RECT 65.005 38.165 65.215 38.985 ;
        RECT 65.385 38.965 65.635 39.565 ;
        RECT 66.910 39.470 67.080 39.615 ;
        RECT 65.805 39.155 66.135 39.405 ;
        RECT 66.345 39.065 66.675 39.435 ;
        RECT 66.910 39.140 67.195 39.470 ;
        RECT 65.385 38.335 65.715 38.965 ;
        RECT 65.885 38.165 66.115 38.985 ;
        RECT 66.910 38.885 67.080 39.140 ;
        RECT 66.415 38.715 67.080 38.885 ;
        RECT 67.365 38.840 67.535 39.640 ;
        RECT 66.415 38.335 66.585 38.715 ;
        RECT 66.765 38.165 67.095 38.545 ;
        RECT 67.275 38.335 67.535 38.840 ;
        RECT 67.705 39.640 67.975 40.545 ;
        RECT 68.145 39.955 68.475 40.715 ;
        RECT 68.655 39.785 68.825 40.545 ;
        RECT 67.705 38.840 67.875 39.640 ;
        RECT 68.160 39.615 68.825 39.785 ;
        RECT 68.160 39.470 68.330 39.615 ;
        RECT 70.005 39.550 70.295 40.715 ;
        RECT 70.525 39.575 70.735 40.715 ;
        RECT 70.905 39.565 71.235 40.545 ;
        RECT 71.405 39.575 71.635 40.715 ;
        RECT 72.310 39.575 72.645 40.545 ;
        RECT 72.815 39.575 72.985 40.715 ;
        RECT 73.155 40.375 75.185 40.545 ;
        RECT 68.045 39.140 68.330 39.470 ;
        RECT 68.160 38.885 68.330 39.140 ;
        RECT 68.565 39.065 68.895 39.435 ;
        RECT 67.705 38.335 67.965 38.840 ;
        RECT 68.160 38.715 68.825 38.885 ;
        RECT 68.145 38.165 68.475 38.545 ;
        RECT 68.655 38.335 68.825 38.715 ;
        RECT 70.005 38.165 70.295 38.890 ;
        RECT 70.525 38.165 70.735 38.985 ;
        RECT 70.905 38.965 71.155 39.565 ;
        RECT 71.325 39.155 71.655 39.405 ;
        RECT 70.905 38.335 71.235 38.965 ;
        RECT 71.405 38.165 71.635 38.985 ;
        RECT 72.310 38.905 72.480 39.575 ;
        RECT 73.155 39.405 73.325 40.375 ;
        RECT 72.650 39.075 72.905 39.405 ;
        RECT 73.130 39.075 73.325 39.405 ;
        RECT 73.495 40.035 74.620 40.205 ;
        RECT 72.735 38.905 72.905 39.075 ;
        RECT 73.495 38.905 73.665 40.035 ;
        RECT 72.310 38.335 72.565 38.905 ;
        RECT 72.735 38.735 73.665 38.905 ;
        RECT 73.835 39.695 74.845 39.865 ;
        RECT 73.835 38.895 74.005 39.695 ;
        RECT 74.210 39.015 74.485 39.495 ;
        RECT 74.205 38.845 74.485 39.015 ;
        RECT 73.490 38.700 73.665 38.735 ;
        RECT 72.735 38.165 73.065 38.565 ;
        RECT 73.490 38.335 74.020 38.700 ;
        RECT 74.210 38.335 74.485 38.845 ;
        RECT 74.655 38.335 74.845 39.695 ;
        RECT 75.015 39.710 75.185 40.375 ;
        RECT 75.355 39.955 75.525 40.715 ;
        RECT 75.760 39.955 76.275 40.365 ;
        RECT 75.015 39.520 75.765 39.710 ;
        RECT 75.935 39.145 76.275 39.955 ;
        RECT 76.445 39.625 78.115 40.715 ;
        RECT 75.045 38.975 76.275 39.145 ;
        RECT 75.025 38.165 75.535 38.700 ;
        RECT 75.755 38.370 76.000 38.975 ;
        RECT 76.445 38.935 77.195 39.455 ;
        RECT 77.365 39.105 78.115 39.625 ;
        RECT 78.490 39.745 78.820 40.545 ;
        RECT 78.990 39.915 79.320 40.715 ;
        RECT 79.620 39.745 79.950 40.545 ;
        RECT 80.595 39.915 80.845 40.715 ;
        RECT 78.490 39.575 80.925 39.745 ;
        RECT 81.115 39.575 81.285 40.715 ;
        RECT 81.455 39.575 81.795 40.545 ;
        RECT 78.285 39.155 78.635 39.405 ;
        RECT 78.820 38.945 78.990 39.575 ;
        RECT 79.160 39.155 79.490 39.355 ;
        RECT 79.660 39.155 79.990 39.355 ;
        RECT 80.160 39.155 80.580 39.355 ;
        RECT 80.755 39.325 80.925 39.575 ;
        RECT 80.755 39.155 81.450 39.325 ;
        RECT 76.445 38.165 78.115 38.935 ;
        RECT 78.490 38.335 78.990 38.945 ;
        RECT 79.620 38.815 80.845 38.985 ;
        RECT 81.620 38.965 81.795 39.575 ;
        RECT 82.425 39.955 82.940 40.365 ;
        RECT 83.175 39.955 83.345 40.715 ;
        RECT 83.515 40.375 85.545 40.545 ;
        RECT 82.425 39.145 82.765 39.955 ;
        RECT 83.515 39.710 83.685 40.375 ;
        RECT 84.080 40.035 85.205 40.205 ;
        RECT 82.935 39.520 83.685 39.710 ;
        RECT 83.855 39.695 84.865 39.865 ;
        RECT 82.425 38.975 83.655 39.145 ;
        RECT 79.620 38.335 79.950 38.815 ;
        RECT 80.120 38.165 80.345 38.625 ;
        RECT 80.515 38.335 80.845 38.815 ;
        RECT 81.035 38.165 81.285 38.965 ;
        RECT 81.455 38.335 81.795 38.965 ;
        RECT 82.700 38.370 82.945 38.975 ;
        RECT 83.165 38.165 83.675 38.700 ;
        RECT 83.855 38.335 84.045 39.695 ;
        RECT 84.215 38.675 84.490 39.495 ;
        RECT 84.695 38.895 84.865 39.695 ;
        RECT 85.035 38.905 85.205 40.035 ;
        RECT 85.375 39.405 85.545 40.375 ;
        RECT 85.715 39.575 85.885 40.715 ;
        RECT 86.055 39.575 86.390 40.545 ;
        RECT 85.375 39.075 85.570 39.405 ;
        RECT 85.795 39.075 86.050 39.405 ;
        RECT 85.795 38.905 85.965 39.075 ;
        RECT 86.220 38.905 86.390 39.575 ;
        RECT 85.035 38.735 85.965 38.905 ;
        RECT 85.035 38.700 85.210 38.735 ;
        RECT 84.215 38.505 84.495 38.675 ;
        RECT 84.215 38.335 84.490 38.505 ;
        RECT 84.680 38.335 85.210 38.700 ;
        RECT 85.635 38.165 85.965 38.565 ;
        RECT 86.135 38.335 86.390 38.905 ;
        RECT 86.565 39.640 86.835 40.545 ;
        RECT 87.005 39.955 87.335 40.715 ;
        RECT 87.515 39.785 87.685 40.545 ;
        RECT 86.565 38.840 86.735 39.640 ;
        RECT 87.020 39.615 87.685 39.785 ;
        RECT 88.150 39.745 88.480 40.545 ;
        RECT 88.650 39.915 88.980 40.715 ;
        RECT 89.280 39.745 89.610 40.545 ;
        RECT 90.255 39.915 90.505 40.715 ;
        RECT 87.020 39.470 87.190 39.615 ;
        RECT 88.150 39.575 90.585 39.745 ;
        RECT 90.775 39.575 90.945 40.715 ;
        RECT 91.115 39.575 91.455 40.545 ;
        RECT 86.905 39.140 87.190 39.470 ;
        RECT 87.020 38.885 87.190 39.140 ;
        RECT 87.425 39.065 87.755 39.435 ;
        RECT 87.945 39.155 88.295 39.405 ;
        RECT 88.480 38.945 88.650 39.575 ;
        RECT 88.820 39.155 89.150 39.355 ;
        RECT 89.320 39.155 89.650 39.355 ;
        RECT 89.820 39.155 90.240 39.355 ;
        RECT 90.415 39.325 90.585 39.575 ;
        RECT 90.415 39.155 91.110 39.325 ;
        RECT 86.565 38.335 86.825 38.840 ;
        RECT 87.020 38.715 87.685 38.885 ;
        RECT 87.005 38.165 87.335 38.545 ;
        RECT 87.515 38.335 87.685 38.715 ;
        RECT 88.150 38.335 88.650 38.945 ;
        RECT 89.280 38.815 90.505 38.985 ;
        RECT 91.280 38.965 91.455 39.575 ;
        RECT 91.625 39.955 92.140 40.365 ;
        RECT 92.375 39.955 92.545 40.715 ;
        RECT 92.715 40.375 94.745 40.545 ;
        RECT 91.625 39.145 91.965 39.955 ;
        RECT 92.715 39.710 92.885 40.375 ;
        RECT 93.280 40.035 94.405 40.205 ;
        RECT 92.135 39.520 92.885 39.710 ;
        RECT 93.055 39.695 94.065 39.865 ;
        RECT 91.625 38.975 92.855 39.145 ;
        RECT 89.280 38.335 89.610 38.815 ;
        RECT 89.780 38.165 90.005 38.625 ;
        RECT 90.175 38.335 90.505 38.815 ;
        RECT 90.695 38.165 90.945 38.965 ;
        RECT 91.115 38.335 91.455 38.965 ;
        RECT 91.900 38.370 92.145 38.975 ;
        RECT 92.365 38.165 92.875 38.700 ;
        RECT 93.055 38.335 93.245 39.695 ;
        RECT 93.415 39.355 93.690 39.495 ;
        RECT 93.415 39.185 93.695 39.355 ;
        RECT 93.415 38.335 93.690 39.185 ;
        RECT 93.895 38.895 94.065 39.695 ;
        RECT 94.235 38.905 94.405 40.035 ;
        RECT 94.575 39.405 94.745 40.375 ;
        RECT 94.915 39.575 95.085 40.715 ;
        RECT 95.255 39.575 95.590 40.545 ;
        RECT 94.575 39.075 94.770 39.405 ;
        RECT 94.995 39.075 95.250 39.405 ;
        RECT 94.995 38.905 95.165 39.075 ;
        RECT 95.420 38.905 95.590 39.575 ;
        RECT 95.765 39.550 96.055 40.715 ;
        RECT 94.235 38.735 95.165 38.905 ;
        RECT 94.235 38.700 94.410 38.735 ;
        RECT 93.880 38.335 94.410 38.700 ;
        RECT 94.835 38.165 95.165 38.565 ;
        RECT 95.335 38.335 95.590 38.905 ;
        RECT 96.690 39.525 96.945 40.405 ;
        RECT 97.115 39.575 97.420 40.715 ;
        RECT 97.760 40.335 98.090 40.715 ;
        RECT 98.270 40.165 98.440 40.455 ;
        RECT 98.610 40.255 98.860 40.715 ;
        RECT 97.640 39.995 98.440 40.165 ;
        RECT 99.030 40.205 99.900 40.545 ;
        RECT 95.765 38.165 96.055 38.890 ;
        RECT 96.690 38.875 96.900 39.525 ;
        RECT 97.640 39.405 97.810 39.995 ;
        RECT 99.030 39.825 99.200 40.205 ;
        RECT 100.135 40.085 100.305 40.545 ;
        RECT 100.475 40.255 100.845 40.715 ;
        RECT 101.140 40.115 101.310 40.455 ;
        RECT 101.480 40.285 101.810 40.715 ;
        RECT 102.045 40.115 102.215 40.455 ;
        RECT 97.980 39.655 99.200 39.825 ;
        RECT 99.370 39.745 99.830 40.035 ;
        RECT 100.135 39.915 100.695 40.085 ;
        RECT 101.140 39.945 102.215 40.115 ;
        RECT 102.385 40.215 103.065 40.545 ;
        RECT 103.280 40.215 103.530 40.545 ;
        RECT 103.700 40.255 103.950 40.715 ;
        RECT 100.525 39.775 100.695 39.915 ;
        RECT 99.370 39.735 100.335 39.745 ;
        RECT 99.030 39.565 99.200 39.655 ;
        RECT 99.660 39.575 100.335 39.735 ;
        RECT 97.070 39.375 97.810 39.405 ;
        RECT 97.070 39.075 97.985 39.375 ;
        RECT 97.660 38.900 97.985 39.075 ;
        RECT 96.690 38.345 96.945 38.875 ;
        RECT 97.115 38.165 97.420 38.625 ;
        RECT 97.665 38.545 97.985 38.900 ;
        RECT 98.155 39.115 98.695 39.485 ;
        RECT 99.030 39.395 99.435 39.565 ;
        RECT 98.155 38.715 98.395 39.115 ;
        RECT 98.875 38.945 99.095 39.225 ;
        RECT 98.565 38.775 99.095 38.945 ;
        RECT 98.565 38.545 98.735 38.775 ;
        RECT 99.265 38.615 99.435 39.395 ;
        RECT 99.605 38.785 99.955 39.405 ;
        RECT 100.125 38.785 100.335 39.575 ;
        RECT 100.525 39.605 102.025 39.775 ;
        RECT 100.525 38.915 100.695 39.605 ;
        RECT 102.385 39.435 102.555 40.215 ;
        RECT 103.360 40.085 103.530 40.215 ;
        RECT 100.865 39.265 102.555 39.435 ;
        RECT 102.725 39.655 103.190 40.045 ;
        RECT 103.360 39.915 103.755 40.085 ;
        RECT 100.865 39.085 101.035 39.265 ;
        RECT 97.665 38.375 98.735 38.545 ;
        RECT 98.905 38.165 99.095 38.605 ;
        RECT 99.265 38.335 100.215 38.615 ;
        RECT 100.525 38.525 100.785 38.915 ;
        RECT 101.205 38.845 101.995 39.095 ;
        RECT 100.435 38.355 100.785 38.525 ;
        RECT 100.995 38.165 101.325 38.625 ;
        RECT 102.200 38.555 102.370 39.265 ;
        RECT 102.725 39.065 102.895 39.655 ;
        RECT 102.540 38.845 102.895 39.065 ;
        RECT 103.065 38.845 103.415 39.465 ;
        RECT 103.585 38.555 103.755 39.915 ;
        RECT 104.120 39.745 104.445 40.530 ;
        RECT 103.925 38.695 104.385 39.745 ;
        RECT 102.200 38.385 103.055 38.555 ;
        RECT 103.260 38.385 103.755 38.555 ;
        RECT 103.925 38.165 104.255 38.525 ;
        RECT 104.615 38.425 104.785 40.545 ;
        RECT 104.955 40.215 105.285 40.715 ;
        RECT 105.455 40.045 105.710 40.545 ;
        RECT 105.885 40.280 111.230 40.715 ;
        RECT 104.960 39.875 105.710 40.045 ;
        RECT 104.960 38.885 105.190 39.875 ;
        RECT 105.360 39.055 105.710 39.705 ;
        RECT 104.960 38.715 105.710 38.885 ;
        RECT 104.955 38.165 105.285 38.545 ;
        RECT 105.455 38.425 105.710 38.715 ;
        RECT 107.470 38.710 107.810 39.540 ;
        RECT 109.290 39.030 109.640 40.280 ;
        RECT 112.325 39.625 113.535 40.715 ;
        RECT 112.325 39.085 112.845 39.625 ;
        RECT 113.015 38.915 113.535 39.455 ;
        RECT 105.885 38.165 111.230 38.710 ;
        RECT 112.325 38.165 113.535 38.915 ;
        RECT 5.520 37.995 113.620 38.165 ;
        RECT 5.605 37.245 6.815 37.995 ;
        RECT 6.985 37.245 8.195 37.995 ;
        RECT 8.370 37.445 8.625 37.735 ;
        RECT 8.795 37.615 9.125 37.995 ;
        RECT 8.370 37.275 9.120 37.445 ;
        RECT 5.605 36.705 6.125 37.245 ;
        RECT 6.295 36.535 6.815 37.075 ;
        RECT 6.985 36.705 7.505 37.245 ;
        RECT 7.675 36.535 8.195 37.075 ;
        RECT 5.605 35.445 6.815 36.535 ;
        RECT 6.985 35.445 8.195 36.535 ;
        RECT 8.370 36.455 8.720 37.105 ;
        RECT 8.890 36.285 9.120 37.275 ;
        RECT 8.370 36.115 9.120 36.285 ;
        RECT 8.370 35.615 8.625 36.115 ;
        RECT 8.795 35.445 9.125 35.945 ;
        RECT 9.295 35.615 9.465 37.735 ;
        RECT 9.825 37.635 10.155 37.995 ;
        RECT 10.325 37.605 10.820 37.775 ;
        RECT 11.025 37.605 11.880 37.775 ;
        RECT 9.695 36.415 10.155 37.465 ;
        RECT 9.635 35.630 9.960 36.415 ;
        RECT 10.325 36.245 10.495 37.605 ;
        RECT 10.665 36.695 11.015 37.315 ;
        RECT 11.185 37.095 11.540 37.315 ;
        RECT 11.185 36.505 11.355 37.095 ;
        RECT 11.710 36.895 11.880 37.605 ;
        RECT 12.755 37.535 13.085 37.995 ;
        RECT 13.295 37.635 13.645 37.805 ;
        RECT 12.085 37.065 12.875 37.315 ;
        RECT 13.295 37.245 13.555 37.635 ;
        RECT 13.865 37.545 14.815 37.825 ;
        RECT 14.985 37.555 15.175 37.995 ;
        RECT 15.345 37.615 16.415 37.785 ;
        RECT 13.045 36.895 13.215 37.075 ;
        RECT 10.325 36.075 10.720 36.245 ;
        RECT 10.890 36.115 11.355 36.505 ;
        RECT 11.525 36.725 13.215 36.895 ;
        RECT 10.550 35.945 10.720 36.075 ;
        RECT 11.525 35.945 11.695 36.725 ;
        RECT 13.385 36.555 13.555 37.245 ;
        RECT 12.055 36.385 13.555 36.555 ;
        RECT 13.745 36.585 13.955 37.375 ;
        RECT 14.125 36.755 14.475 37.375 ;
        RECT 14.645 36.765 14.815 37.545 ;
        RECT 15.345 37.385 15.515 37.615 ;
        RECT 14.985 37.215 15.515 37.385 ;
        RECT 14.985 36.935 15.205 37.215 ;
        RECT 15.685 37.045 15.925 37.445 ;
        RECT 14.645 36.595 15.050 36.765 ;
        RECT 15.385 36.675 15.925 37.045 ;
        RECT 16.095 37.260 16.415 37.615 ;
        RECT 16.660 37.535 16.965 37.995 ;
        RECT 17.135 37.285 17.390 37.815 ;
        RECT 16.095 37.085 16.420 37.260 ;
        RECT 16.095 36.785 17.010 37.085 ;
        RECT 16.270 36.755 17.010 36.785 ;
        RECT 13.745 36.425 14.420 36.585 ;
        RECT 14.880 36.505 15.050 36.595 ;
        RECT 13.745 36.415 14.710 36.425 ;
        RECT 13.385 36.245 13.555 36.385 ;
        RECT 10.130 35.445 10.380 35.905 ;
        RECT 10.550 35.615 10.800 35.945 ;
        RECT 11.015 35.615 11.695 35.945 ;
        RECT 11.865 36.045 12.940 36.215 ;
        RECT 13.385 36.075 13.945 36.245 ;
        RECT 14.250 36.125 14.710 36.415 ;
        RECT 14.880 36.335 16.100 36.505 ;
        RECT 11.865 35.705 12.035 36.045 ;
        RECT 12.270 35.445 12.600 35.875 ;
        RECT 12.770 35.705 12.940 36.045 ;
        RECT 13.235 35.445 13.605 35.905 ;
        RECT 13.775 35.615 13.945 36.075 ;
        RECT 14.880 35.955 15.050 36.335 ;
        RECT 16.270 36.165 16.440 36.755 ;
        RECT 17.180 36.635 17.390 37.285 ;
        RECT 14.180 35.615 15.050 35.955 ;
        RECT 15.640 35.995 16.440 36.165 ;
        RECT 15.220 35.445 15.470 35.905 ;
        RECT 15.640 35.705 15.810 35.995 ;
        RECT 15.990 35.445 16.320 35.825 ;
        RECT 16.660 35.445 16.965 36.585 ;
        RECT 17.135 35.755 17.390 36.635 ;
        RECT 17.570 37.255 17.825 37.825 ;
        RECT 17.995 37.595 18.325 37.995 ;
        RECT 18.750 37.460 19.280 37.825 ;
        RECT 19.470 37.655 19.745 37.825 ;
        RECT 19.465 37.485 19.745 37.655 ;
        RECT 18.750 37.425 18.925 37.460 ;
        RECT 17.995 37.255 18.925 37.425 ;
        RECT 17.570 36.585 17.740 37.255 ;
        RECT 17.995 37.085 18.165 37.255 ;
        RECT 17.910 36.755 18.165 37.085 ;
        RECT 18.390 36.755 18.585 37.085 ;
        RECT 17.570 35.615 17.905 36.585 ;
        RECT 18.075 35.445 18.245 36.585 ;
        RECT 18.415 35.785 18.585 36.755 ;
        RECT 18.755 36.125 18.925 37.255 ;
        RECT 19.095 36.465 19.265 37.265 ;
        RECT 19.470 36.665 19.745 37.485 ;
        RECT 19.915 36.465 20.105 37.825 ;
        RECT 20.285 37.460 20.795 37.995 ;
        RECT 21.015 37.185 21.260 37.790 ;
        RECT 21.705 37.225 24.295 37.995 ;
        RECT 24.470 37.255 24.725 37.825 ;
        RECT 24.895 37.595 25.225 37.995 ;
        RECT 25.650 37.460 26.180 37.825 ;
        RECT 25.650 37.425 25.825 37.460 ;
        RECT 24.895 37.255 25.825 37.425 ;
        RECT 20.305 37.015 21.535 37.185 ;
        RECT 19.095 36.295 20.105 36.465 ;
        RECT 20.275 36.450 21.025 36.640 ;
        RECT 18.755 35.955 19.880 36.125 ;
        RECT 20.275 35.785 20.445 36.450 ;
        RECT 21.195 36.205 21.535 37.015 ;
        RECT 21.705 36.705 22.915 37.225 ;
        RECT 23.085 36.535 24.295 37.055 ;
        RECT 18.415 35.615 20.445 35.785 ;
        RECT 20.615 35.445 20.785 36.205 ;
        RECT 21.020 35.795 21.535 36.205 ;
        RECT 21.705 35.445 24.295 36.535 ;
        RECT 24.470 36.585 24.640 37.255 ;
        RECT 24.895 37.085 25.065 37.255 ;
        RECT 24.810 36.755 25.065 37.085 ;
        RECT 25.290 36.755 25.485 37.085 ;
        RECT 24.470 35.615 24.805 36.585 ;
        RECT 24.975 35.445 25.145 36.585 ;
        RECT 25.315 35.785 25.485 36.755 ;
        RECT 25.655 36.125 25.825 37.255 ;
        RECT 25.995 36.465 26.165 37.265 ;
        RECT 26.370 36.975 26.645 37.825 ;
        RECT 26.365 36.805 26.645 36.975 ;
        RECT 26.370 36.665 26.645 36.805 ;
        RECT 26.815 36.465 27.005 37.825 ;
        RECT 27.185 37.460 27.695 37.995 ;
        RECT 27.915 37.185 28.160 37.790 ;
        RECT 29.155 37.445 29.325 37.825 ;
        RECT 29.505 37.615 29.835 37.995 ;
        RECT 29.155 37.275 29.820 37.445 ;
        RECT 30.015 37.320 30.275 37.825 ;
        RECT 27.205 37.015 28.435 37.185 ;
        RECT 25.995 36.295 27.005 36.465 ;
        RECT 27.175 36.450 27.925 36.640 ;
        RECT 25.655 35.955 26.780 36.125 ;
        RECT 27.175 35.785 27.345 36.450 ;
        RECT 28.095 36.205 28.435 37.015 ;
        RECT 29.085 36.725 29.415 37.095 ;
        RECT 29.650 37.020 29.820 37.275 ;
        RECT 29.650 36.690 29.935 37.020 ;
        RECT 29.650 36.545 29.820 36.690 ;
        RECT 25.315 35.615 27.345 35.785 ;
        RECT 27.515 35.445 27.685 36.205 ;
        RECT 27.920 35.795 28.435 36.205 ;
        RECT 29.155 36.375 29.820 36.545 ;
        RECT 30.105 36.520 30.275 37.320 ;
        RECT 31.365 37.270 31.655 37.995 ;
        RECT 31.830 37.255 32.085 37.825 ;
        RECT 32.255 37.595 32.585 37.995 ;
        RECT 33.010 37.460 33.540 37.825 ;
        RECT 33.010 37.425 33.185 37.460 ;
        RECT 32.255 37.255 33.185 37.425 ;
        RECT 29.155 35.615 29.325 36.375 ;
        RECT 29.505 35.445 29.835 36.205 ;
        RECT 30.005 35.615 30.275 36.520 ;
        RECT 31.365 35.445 31.655 36.610 ;
        RECT 31.830 36.585 32.000 37.255 ;
        RECT 32.255 37.085 32.425 37.255 ;
        RECT 32.170 36.755 32.425 37.085 ;
        RECT 32.650 36.755 32.845 37.085 ;
        RECT 31.830 35.615 32.165 36.585 ;
        RECT 32.335 35.445 32.505 36.585 ;
        RECT 32.675 35.785 32.845 36.755 ;
        RECT 33.015 36.125 33.185 37.255 ;
        RECT 33.355 36.465 33.525 37.265 ;
        RECT 33.730 36.975 34.005 37.825 ;
        RECT 33.725 36.805 34.005 36.975 ;
        RECT 33.730 36.665 34.005 36.805 ;
        RECT 34.175 36.465 34.365 37.825 ;
        RECT 34.545 37.460 35.055 37.995 ;
        RECT 35.275 37.185 35.520 37.790 ;
        RECT 35.965 37.225 37.635 37.995 ;
        RECT 38.270 37.445 38.525 37.735 ;
        RECT 38.695 37.615 39.025 37.995 ;
        RECT 38.270 37.275 39.020 37.445 ;
        RECT 34.565 37.015 35.795 37.185 ;
        RECT 33.355 36.295 34.365 36.465 ;
        RECT 34.535 36.450 35.285 36.640 ;
        RECT 33.015 35.955 34.140 36.125 ;
        RECT 34.535 35.785 34.705 36.450 ;
        RECT 35.455 36.205 35.795 37.015 ;
        RECT 35.965 36.705 36.715 37.225 ;
        RECT 36.885 36.535 37.635 37.055 ;
        RECT 32.675 35.615 34.705 35.785 ;
        RECT 34.875 35.445 35.045 36.205 ;
        RECT 35.280 35.795 35.795 36.205 ;
        RECT 35.965 35.445 37.635 36.535 ;
        RECT 38.270 36.455 38.620 37.105 ;
        RECT 38.790 36.285 39.020 37.275 ;
        RECT 38.270 36.115 39.020 36.285 ;
        RECT 38.270 35.615 38.525 36.115 ;
        RECT 38.695 35.445 39.025 35.945 ;
        RECT 39.195 35.615 39.365 37.735 ;
        RECT 39.725 37.635 40.055 37.995 ;
        RECT 40.225 37.605 40.720 37.775 ;
        RECT 40.925 37.605 41.780 37.775 ;
        RECT 39.595 36.415 40.055 37.465 ;
        RECT 39.535 35.630 39.860 36.415 ;
        RECT 40.225 36.245 40.395 37.605 ;
        RECT 40.565 36.695 40.915 37.315 ;
        RECT 41.085 37.095 41.440 37.315 ;
        RECT 41.085 36.505 41.255 37.095 ;
        RECT 41.610 36.895 41.780 37.605 ;
        RECT 42.655 37.535 42.985 37.995 ;
        RECT 43.195 37.635 43.545 37.805 ;
        RECT 41.985 37.065 42.775 37.315 ;
        RECT 43.195 37.245 43.455 37.635 ;
        RECT 43.765 37.545 44.715 37.825 ;
        RECT 44.885 37.555 45.075 37.995 ;
        RECT 45.245 37.615 46.315 37.785 ;
        RECT 42.945 36.895 43.115 37.075 ;
        RECT 40.225 36.075 40.620 36.245 ;
        RECT 40.790 36.115 41.255 36.505 ;
        RECT 41.425 36.725 43.115 36.895 ;
        RECT 40.450 35.945 40.620 36.075 ;
        RECT 41.425 35.945 41.595 36.725 ;
        RECT 43.285 36.555 43.455 37.245 ;
        RECT 41.955 36.385 43.455 36.555 ;
        RECT 43.645 36.585 43.855 37.375 ;
        RECT 44.025 36.755 44.375 37.375 ;
        RECT 44.545 36.765 44.715 37.545 ;
        RECT 45.245 37.385 45.415 37.615 ;
        RECT 44.885 37.215 45.415 37.385 ;
        RECT 44.885 36.935 45.105 37.215 ;
        RECT 45.585 37.045 45.825 37.445 ;
        RECT 44.545 36.595 44.950 36.765 ;
        RECT 45.285 36.675 45.825 37.045 ;
        RECT 45.995 37.260 46.315 37.615 ;
        RECT 46.560 37.535 46.865 37.995 ;
        RECT 47.035 37.285 47.290 37.815 ;
        RECT 45.995 37.085 46.320 37.260 ;
        RECT 45.995 36.785 46.910 37.085 ;
        RECT 46.170 36.755 46.910 36.785 ;
        RECT 43.645 36.425 44.320 36.585 ;
        RECT 44.780 36.505 44.950 36.595 ;
        RECT 43.645 36.415 44.610 36.425 ;
        RECT 43.285 36.245 43.455 36.385 ;
        RECT 40.030 35.445 40.280 35.905 ;
        RECT 40.450 35.615 40.700 35.945 ;
        RECT 40.915 35.615 41.595 35.945 ;
        RECT 41.765 36.045 42.840 36.215 ;
        RECT 43.285 36.075 43.845 36.245 ;
        RECT 44.150 36.125 44.610 36.415 ;
        RECT 44.780 36.335 46.000 36.505 ;
        RECT 41.765 35.705 41.935 36.045 ;
        RECT 42.170 35.445 42.500 35.875 ;
        RECT 42.670 35.705 42.840 36.045 ;
        RECT 43.135 35.445 43.505 35.905 ;
        RECT 43.675 35.615 43.845 36.075 ;
        RECT 44.780 35.955 44.950 36.335 ;
        RECT 46.170 36.165 46.340 36.755 ;
        RECT 47.080 36.635 47.290 37.285 ;
        RECT 47.505 37.175 47.735 37.995 ;
        RECT 47.905 37.195 48.235 37.825 ;
        RECT 47.485 36.755 47.815 37.005 ;
        RECT 44.080 35.615 44.950 35.955 ;
        RECT 45.540 35.995 46.340 36.165 ;
        RECT 45.120 35.445 45.370 35.905 ;
        RECT 45.540 35.705 45.710 35.995 ;
        RECT 45.890 35.445 46.220 35.825 ;
        RECT 46.560 35.445 46.865 36.585 ;
        RECT 47.035 35.755 47.290 36.635 ;
        RECT 47.985 36.595 48.235 37.195 ;
        RECT 48.405 37.175 48.615 37.995 ;
        RECT 48.845 37.450 54.190 37.995 ;
        RECT 50.430 36.620 50.770 37.450 ;
        RECT 54.365 37.225 56.955 37.995 ;
        RECT 57.125 37.270 57.415 37.995 ;
        RECT 47.505 35.445 47.735 36.585 ;
        RECT 47.905 35.615 48.235 36.595 ;
        RECT 48.405 35.445 48.615 36.585 ;
        RECT 52.250 35.880 52.600 37.130 ;
        RECT 54.365 36.705 55.575 37.225 ;
        RECT 58.505 37.175 58.765 37.995 ;
        RECT 58.935 37.355 59.265 37.825 ;
        RECT 59.435 37.525 59.605 37.995 ;
        RECT 59.775 37.355 60.105 37.825 ;
        RECT 60.275 37.525 61.000 37.995 ;
        RECT 61.170 37.355 61.500 37.825 ;
        RECT 61.670 37.525 61.840 37.995 ;
        RECT 62.010 37.355 62.340 37.825 ;
        RECT 58.935 37.175 62.340 37.355 ;
        RECT 62.510 37.185 62.715 37.995 ;
        RECT 55.745 36.535 56.955 37.055 ;
        RECT 62.135 37.005 62.340 37.175 ;
        RECT 62.885 37.175 63.240 37.700 ;
        RECT 63.410 37.255 63.660 37.995 ;
        RECT 64.025 37.225 67.535 37.995 ;
        RECT 67.705 37.245 68.915 37.995 ;
        RECT 69.090 37.445 69.345 37.735 ;
        RECT 69.515 37.615 69.845 37.995 ;
        RECT 69.090 37.275 69.840 37.445 ;
        RECT 62.885 37.005 63.055 37.175 ;
        RECT 58.520 36.795 59.660 37.005 ;
        RECT 59.840 36.795 61.055 37.005 ;
        RECT 61.235 36.795 61.955 37.005 ;
        RECT 62.135 36.625 62.455 37.005 ;
        RECT 62.740 36.835 63.055 37.005 ;
        RECT 48.845 35.445 54.190 35.880 ;
        RECT 54.365 35.445 56.955 36.535 ;
        RECT 57.125 35.445 57.415 36.610 ;
        RECT 58.505 36.455 60.525 36.625 ;
        RECT 58.505 35.615 58.845 36.455 ;
        RECT 59.015 35.445 59.225 36.285 ;
        RECT 59.395 35.615 59.645 36.455 ;
        RECT 59.815 35.785 60.025 36.285 ;
        RECT 60.195 35.955 60.525 36.455 ;
        RECT 60.695 36.455 61.880 36.625 ;
        RECT 60.695 35.955 61.080 36.455 ;
        RECT 61.250 35.785 61.460 36.285 ;
        RECT 59.815 35.615 61.460 35.785 ;
        RECT 61.630 35.785 61.880 36.455 ;
        RECT 62.050 36.455 62.455 36.625 ;
        RECT 62.050 35.955 62.300 36.455 ;
        RECT 62.470 35.785 62.715 36.285 ;
        RECT 61.630 35.615 62.715 35.785 ;
        RECT 62.885 36.045 63.055 36.835 ;
        RECT 63.225 36.795 63.855 37.005 ;
        RECT 63.605 36.125 63.855 36.795 ;
        RECT 64.025 36.705 65.675 37.225 ;
        RECT 65.845 36.535 67.535 37.055 ;
        RECT 67.705 36.705 68.225 37.245 ;
        RECT 68.395 36.535 68.915 37.075 ;
        RECT 62.885 35.630 63.240 36.045 ;
        RECT 63.410 35.445 63.660 35.945 ;
        RECT 64.025 35.445 67.535 36.535 ;
        RECT 67.705 35.445 68.915 36.535 ;
        RECT 69.090 36.455 69.440 37.105 ;
        RECT 69.610 36.285 69.840 37.275 ;
        RECT 69.090 36.115 69.840 36.285 ;
        RECT 69.090 35.615 69.345 36.115 ;
        RECT 69.515 35.445 69.845 35.945 ;
        RECT 70.015 35.615 70.185 37.735 ;
        RECT 70.545 37.635 70.875 37.995 ;
        RECT 71.045 37.605 71.540 37.775 ;
        RECT 71.745 37.605 72.600 37.775 ;
        RECT 70.415 36.415 70.875 37.465 ;
        RECT 70.355 35.630 70.680 36.415 ;
        RECT 71.045 36.245 71.215 37.605 ;
        RECT 71.385 36.695 71.735 37.315 ;
        RECT 71.905 37.095 72.260 37.315 ;
        RECT 71.905 36.505 72.075 37.095 ;
        RECT 72.430 36.895 72.600 37.605 ;
        RECT 73.475 37.535 73.805 37.995 ;
        RECT 74.015 37.635 74.365 37.805 ;
        RECT 72.805 37.065 73.595 37.315 ;
        RECT 74.015 37.245 74.275 37.635 ;
        RECT 74.585 37.545 75.535 37.825 ;
        RECT 75.705 37.555 75.895 37.995 ;
        RECT 76.065 37.615 77.135 37.785 ;
        RECT 73.765 36.895 73.935 37.075 ;
        RECT 71.045 36.075 71.440 36.245 ;
        RECT 71.610 36.115 72.075 36.505 ;
        RECT 72.245 36.725 73.935 36.895 ;
        RECT 71.270 35.945 71.440 36.075 ;
        RECT 72.245 35.945 72.415 36.725 ;
        RECT 74.105 36.555 74.275 37.245 ;
        RECT 72.775 36.385 74.275 36.555 ;
        RECT 74.465 36.585 74.675 37.375 ;
        RECT 74.845 36.755 75.195 37.375 ;
        RECT 75.365 36.765 75.535 37.545 ;
        RECT 76.065 37.385 76.235 37.615 ;
        RECT 75.705 37.215 76.235 37.385 ;
        RECT 75.705 36.935 75.925 37.215 ;
        RECT 76.405 37.045 76.645 37.445 ;
        RECT 75.365 36.595 75.770 36.765 ;
        RECT 76.105 36.675 76.645 37.045 ;
        RECT 76.815 37.260 77.135 37.615 ;
        RECT 77.380 37.535 77.685 37.995 ;
        RECT 77.855 37.285 78.110 37.815 ;
        RECT 76.815 37.085 77.140 37.260 ;
        RECT 76.815 36.785 77.730 37.085 ;
        RECT 76.990 36.755 77.730 36.785 ;
        RECT 74.465 36.425 75.140 36.585 ;
        RECT 75.600 36.505 75.770 36.595 ;
        RECT 74.465 36.415 75.430 36.425 ;
        RECT 74.105 36.245 74.275 36.385 ;
        RECT 70.850 35.445 71.100 35.905 ;
        RECT 71.270 35.615 71.520 35.945 ;
        RECT 71.735 35.615 72.415 35.945 ;
        RECT 72.585 36.045 73.660 36.215 ;
        RECT 74.105 36.075 74.665 36.245 ;
        RECT 74.970 36.125 75.430 36.415 ;
        RECT 75.600 36.335 76.820 36.505 ;
        RECT 72.585 35.705 72.755 36.045 ;
        RECT 72.990 35.445 73.320 35.875 ;
        RECT 73.490 35.705 73.660 36.045 ;
        RECT 73.955 35.445 74.325 35.905 ;
        RECT 74.495 35.615 74.665 36.075 ;
        RECT 75.600 35.955 75.770 36.335 ;
        RECT 76.990 36.165 77.160 36.755 ;
        RECT 77.900 36.635 78.110 37.285 ;
        RECT 78.345 37.175 78.555 37.995 ;
        RECT 78.725 37.195 79.055 37.825 ;
        RECT 74.900 35.615 75.770 35.955 ;
        RECT 76.360 35.995 77.160 36.165 ;
        RECT 75.940 35.445 76.190 35.905 ;
        RECT 76.360 35.705 76.530 35.995 ;
        RECT 76.710 35.445 77.040 35.825 ;
        RECT 77.380 35.445 77.685 36.585 ;
        RECT 77.855 35.755 78.110 36.635 ;
        RECT 78.725 36.595 78.975 37.195 ;
        RECT 79.225 37.175 79.455 37.995 ;
        RECT 79.665 37.225 82.255 37.995 ;
        RECT 82.885 37.270 83.175 37.995 ;
        RECT 83.345 37.225 86.855 37.995 ;
        RECT 79.145 36.755 79.475 37.005 ;
        RECT 79.665 36.705 80.875 37.225 ;
        RECT 78.345 35.445 78.555 36.585 ;
        RECT 78.725 35.615 79.055 36.595 ;
        RECT 79.225 35.445 79.455 36.585 ;
        RECT 81.045 36.535 82.255 37.055 ;
        RECT 83.345 36.705 84.995 37.225 ;
        RECT 87.985 37.175 88.215 37.995 ;
        RECT 88.385 37.195 88.715 37.825 ;
        RECT 79.665 35.445 82.255 36.535 ;
        RECT 82.885 35.445 83.175 36.610 ;
        RECT 85.165 36.535 86.855 37.055 ;
        RECT 87.965 36.755 88.295 37.005 ;
        RECT 88.465 36.595 88.715 37.195 ;
        RECT 88.885 37.175 89.095 37.995 ;
        RECT 90.450 37.215 90.950 37.825 ;
        RECT 90.245 36.755 90.595 37.005 ;
        RECT 83.345 35.445 86.855 36.535 ;
        RECT 87.985 35.445 88.215 36.585 ;
        RECT 88.385 35.615 88.715 36.595 ;
        RECT 90.780 36.585 90.950 37.215 ;
        RECT 91.580 37.345 91.910 37.825 ;
        RECT 92.080 37.535 92.305 37.995 ;
        RECT 92.475 37.345 92.805 37.825 ;
        RECT 91.580 37.175 92.805 37.345 ;
        RECT 92.995 37.195 93.245 37.995 ;
        RECT 93.415 37.195 93.755 37.825 ;
        RECT 94.015 37.445 94.185 37.825 ;
        RECT 94.365 37.615 94.695 37.995 ;
        RECT 94.015 37.275 94.680 37.445 ;
        RECT 94.875 37.320 95.135 37.825 ;
        RECT 91.120 36.805 91.450 37.005 ;
        RECT 91.620 36.805 91.950 37.005 ;
        RECT 92.120 36.805 92.540 37.005 ;
        RECT 92.715 36.835 93.410 37.005 ;
        RECT 92.715 36.585 92.885 36.835 ;
        RECT 93.580 36.585 93.755 37.195 ;
        RECT 93.945 36.725 94.275 37.095 ;
        RECT 94.510 37.020 94.680 37.275 ;
        RECT 88.885 35.445 89.095 36.585 ;
        RECT 90.450 36.415 92.885 36.585 ;
        RECT 90.450 35.615 90.780 36.415 ;
        RECT 90.950 35.445 91.280 36.245 ;
        RECT 91.580 35.615 91.910 36.415 ;
        RECT 92.555 35.445 92.805 36.245 ;
        RECT 93.075 35.445 93.245 36.585 ;
        RECT 93.415 35.615 93.755 36.585 ;
        RECT 94.510 36.690 94.795 37.020 ;
        RECT 94.510 36.545 94.680 36.690 ;
        RECT 94.015 36.375 94.680 36.545 ;
        RECT 94.965 36.520 95.135 37.320 ;
        RECT 95.305 37.245 96.515 37.995 ;
        RECT 95.305 36.705 95.825 37.245 ;
        RECT 96.960 37.185 97.205 37.790 ;
        RECT 97.425 37.460 97.935 37.995 ;
        RECT 95.995 36.535 96.515 37.075 ;
        RECT 94.015 35.615 94.185 36.375 ;
        RECT 94.365 35.445 94.695 36.205 ;
        RECT 94.865 35.615 95.135 36.520 ;
        RECT 95.305 35.445 96.515 36.535 ;
        RECT 96.685 37.015 97.915 37.185 ;
        RECT 96.685 36.205 97.025 37.015 ;
        RECT 97.195 36.450 97.945 36.640 ;
        RECT 96.685 35.795 97.200 36.205 ;
        RECT 97.435 35.445 97.605 36.205 ;
        RECT 97.775 35.785 97.945 36.450 ;
        RECT 98.115 36.465 98.305 37.825 ;
        RECT 98.475 36.975 98.750 37.825 ;
        RECT 98.940 37.460 99.470 37.825 ;
        RECT 99.895 37.595 100.225 37.995 ;
        RECT 99.295 37.425 99.470 37.460 ;
        RECT 98.475 36.805 98.755 36.975 ;
        RECT 98.475 36.665 98.750 36.805 ;
        RECT 98.955 36.465 99.125 37.265 ;
        RECT 98.115 36.295 99.125 36.465 ;
        RECT 99.295 37.255 100.225 37.425 ;
        RECT 100.395 37.255 100.650 37.825 ;
        RECT 100.915 37.445 101.085 37.825 ;
        RECT 101.265 37.615 101.595 37.995 ;
        RECT 100.915 37.275 101.580 37.445 ;
        RECT 101.775 37.320 102.035 37.825 ;
        RECT 99.295 36.125 99.465 37.255 ;
        RECT 100.055 37.085 100.225 37.255 ;
        RECT 98.340 35.955 99.465 36.125 ;
        RECT 99.635 36.755 99.830 37.085 ;
        RECT 100.055 36.755 100.310 37.085 ;
        RECT 99.635 35.785 99.805 36.755 ;
        RECT 100.480 36.585 100.650 37.255 ;
        RECT 100.845 36.725 101.175 37.095 ;
        RECT 101.410 37.020 101.580 37.275 ;
        RECT 97.775 35.615 99.805 35.785 ;
        RECT 99.975 35.445 100.145 36.585 ;
        RECT 100.315 35.615 100.650 36.585 ;
        RECT 101.410 36.690 101.695 37.020 ;
        RECT 101.410 36.545 101.580 36.690 ;
        RECT 100.915 36.375 101.580 36.545 ;
        RECT 101.865 36.520 102.035 37.320 ;
        RECT 102.265 37.175 102.475 37.995 ;
        RECT 102.645 37.195 102.975 37.825 ;
        RECT 102.645 36.595 102.895 37.195 ;
        RECT 103.145 37.175 103.375 37.995 ;
        RECT 103.585 37.225 107.095 37.995 ;
        RECT 107.265 37.245 108.475 37.995 ;
        RECT 108.645 37.270 108.935 37.995 ;
        RECT 103.065 36.755 103.395 37.005 ;
        RECT 103.585 36.705 105.235 37.225 ;
        RECT 100.915 35.615 101.085 36.375 ;
        RECT 101.265 35.445 101.595 36.205 ;
        RECT 101.765 35.615 102.035 36.520 ;
        RECT 102.265 35.445 102.475 36.585 ;
        RECT 102.645 35.615 102.975 36.595 ;
        RECT 103.145 35.445 103.375 36.585 ;
        RECT 105.405 36.535 107.095 37.055 ;
        RECT 107.265 36.705 107.785 37.245 ;
        RECT 109.105 37.225 111.695 37.995 ;
        RECT 112.325 37.245 113.535 37.995 ;
        RECT 107.955 36.535 108.475 37.075 ;
        RECT 109.105 36.705 110.315 37.225 ;
        RECT 103.585 35.445 107.095 36.535 ;
        RECT 107.265 35.445 108.475 36.535 ;
        RECT 108.645 35.445 108.935 36.610 ;
        RECT 110.485 36.535 111.695 37.055 ;
        RECT 109.105 35.445 111.695 36.535 ;
        RECT 112.325 36.535 112.845 37.075 ;
        RECT 113.015 36.705 113.535 37.245 ;
        RECT 112.325 35.445 113.535 36.535 ;
        RECT 5.520 35.275 113.620 35.445 ;
        RECT 5.605 34.185 6.815 35.275 ;
        RECT 6.985 34.185 8.655 35.275 ;
        RECT 8.830 34.605 9.085 35.105 ;
        RECT 9.255 34.775 9.585 35.275 ;
        RECT 8.830 34.435 9.580 34.605 ;
        RECT 5.605 33.475 6.125 34.015 ;
        RECT 6.295 33.645 6.815 34.185 ;
        RECT 6.985 33.495 7.735 34.015 ;
        RECT 7.905 33.665 8.655 34.185 ;
        RECT 8.830 33.615 9.180 34.265 ;
        RECT 5.605 32.725 6.815 33.475 ;
        RECT 6.985 32.725 8.655 33.495 ;
        RECT 9.350 33.445 9.580 34.435 ;
        RECT 8.830 33.275 9.580 33.445 ;
        RECT 8.830 32.985 9.085 33.275 ;
        RECT 9.255 32.725 9.585 33.105 ;
        RECT 9.755 32.985 9.925 35.105 ;
        RECT 10.095 34.305 10.420 35.090 ;
        RECT 10.590 34.815 10.840 35.275 ;
        RECT 11.010 34.775 11.260 35.105 ;
        RECT 11.475 34.775 12.155 35.105 ;
        RECT 11.010 34.645 11.180 34.775 ;
        RECT 10.785 34.475 11.180 34.645 ;
        RECT 10.155 33.255 10.615 34.305 ;
        RECT 10.785 33.115 10.955 34.475 ;
        RECT 11.350 34.215 11.815 34.605 ;
        RECT 11.125 33.405 11.475 34.025 ;
        RECT 11.645 33.625 11.815 34.215 ;
        RECT 11.985 33.995 12.155 34.775 ;
        RECT 12.325 34.675 12.495 35.015 ;
        RECT 12.730 34.845 13.060 35.275 ;
        RECT 13.230 34.675 13.400 35.015 ;
        RECT 13.695 34.815 14.065 35.275 ;
        RECT 12.325 34.505 13.400 34.675 ;
        RECT 14.235 34.645 14.405 35.105 ;
        RECT 14.640 34.765 15.510 35.105 ;
        RECT 15.680 34.815 15.930 35.275 ;
        RECT 13.845 34.475 14.405 34.645 ;
        RECT 13.845 34.335 14.015 34.475 ;
        RECT 12.515 34.165 14.015 34.335 ;
        RECT 14.710 34.305 15.170 34.595 ;
        RECT 11.985 33.825 13.675 33.995 ;
        RECT 11.645 33.405 12.000 33.625 ;
        RECT 12.170 33.115 12.340 33.825 ;
        RECT 12.545 33.405 13.335 33.655 ;
        RECT 13.505 33.645 13.675 33.825 ;
        RECT 13.845 33.475 14.015 34.165 ;
        RECT 10.285 32.725 10.615 33.085 ;
        RECT 10.785 32.945 11.280 33.115 ;
        RECT 11.485 32.945 12.340 33.115 ;
        RECT 13.215 32.725 13.545 33.185 ;
        RECT 13.755 33.085 14.015 33.475 ;
        RECT 14.205 34.295 15.170 34.305 ;
        RECT 15.340 34.385 15.510 34.765 ;
        RECT 16.100 34.725 16.270 35.015 ;
        RECT 16.450 34.895 16.780 35.275 ;
        RECT 16.100 34.555 16.900 34.725 ;
        RECT 14.205 34.135 14.880 34.295 ;
        RECT 15.340 34.215 16.560 34.385 ;
        RECT 14.205 33.345 14.415 34.135 ;
        RECT 15.340 34.125 15.510 34.215 ;
        RECT 14.585 33.345 14.935 33.965 ;
        RECT 15.105 33.955 15.510 34.125 ;
        RECT 15.105 33.175 15.275 33.955 ;
        RECT 15.445 33.505 15.665 33.785 ;
        RECT 15.845 33.675 16.385 34.045 ;
        RECT 16.730 33.965 16.900 34.555 ;
        RECT 17.120 34.135 17.425 35.275 ;
        RECT 17.595 34.085 17.850 34.965 ;
        RECT 18.485 34.110 18.775 35.275 ;
        RECT 18.950 34.135 19.285 35.105 ;
        RECT 19.455 34.135 19.625 35.275 ;
        RECT 19.795 34.935 21.825 35.105 ;
        RECT 16.730 33.935 17.470 33.965 ;
        RECT 15.445 33.335 15.975 33.505 ;
        RECT 13.755 32.915 14.105 33.085 ;
        RECT 14.325 32.895 15.275 33.175 ;
        RECT 15.445 32.725 15.635 33.165 ;
        RECT 15.805 33.105 15.975 33.335 ;
        RECT 16.145 33.275 16.385 33.675 ;
        RECT 16.555 33.635 17.470 33.935 ;
        RECT 16.555 33.460 16.880 33.635 ;
        RECT 16.555 33.105 16.875 33.460 ;
        RECT 17.640 33.435 17.850 34.085 ;
        RECT 18.950 33.465 19.120 34.135 ;
        RECT 19.795 33.965 19.965 34.935 ;
        RECT 19.290 33.635 19.545 33.965 ;
        RECT 19.770 33.635 19.965 33.965 ;
        RECT 20.135 34.595 21.260 34.765 ;
        RECT 19.375 33.465 19.545 33.635 ;
        RECT 20.135 33.465 20.305 34.595 ;
        RECT 15.805 32.935 16.875 33.105 ;
        RECT 17.120 32.725 17.425 33.185 ;
        RECT 17.595 32.905 17.850 33.435 ;
        RECT 18.485 32.725 18.775 33.450 ;
        RECT 18.950 32.895 19.205 33.465 ;
        RECT 19.375 33.295 20.305 33.465 ;
        RECT 20.475 34.255 21.485 34.425 ;
        RECT 20.475 33.455 20.645 34.255 ;
        RECT 20.850 33.915 21.125 34.055 ;
        RECT 20.845 33.745 21.125 33.915 ;
        RECT 20.130 33.260 20.305 33.295 ;
        RECT 19.375 32.725 19.705 33.125 ;
        RECT 20.130 32.895 20.660 33.260 ;
        RECT 20.850 32.895 21.125 33.745 ;
        RECT 21.295 32.895 21.485 34.255 ;
        RECT 21.655 34.270 21.825 34.935 ;
        RECT 21.995 34.515 22.165 35.275 ;
        RECT 22.400 34.515 22.915 34.925 ;
        RECT 21.655 34.080 22.405 34.270 ;
        RECT 22.575 33.705 22.915 34.515 ;
        RECT 24.010 34.605 24.265 35.105 ;
        RECT 24.435 34.775 24.765 35.275 ;
        RECT 24.010 34.435 24.760 34.605 ;
        RECT 21.685 33.535 22.915 33.705 ;
        RECT 24.010 33.615 24.360 34.265 ;
        RECT 21.665 32.725 22.175 33.260 ;
        RECT 22.395 32.930 22.640 33.535 ;
        RECT 24.530 33.445 24.760 34.435 ;
        RECT 24.010 33.275 24.760 33.445 ;
        RECT 24.010 32.985 24.265 33.275 ;
        RECT 24.435 32.725 24.765 33.105 ;
        RECT 24.935 32.985 25.105 35.105 ;
        RECT 25.275 34.305 25.600 35.090 ;
        RECT 25.770 34.815 26.020 35.275 ;
        RECT 26.190 34.775 26.440 35.105 ;
        RECT 26.655 34.775 27.335 35.105 ;
        RECT 26.190 34.645 26.360 34.775 ;
        RECT 25.965 34.475 26.360 34.645 ;
        RECT 25.335 33.255 25.795 34.305 ;
        RECT 25.965 33.115 26.135 34.475 ;
        RECT 26.530 34.215 26.995 34.605 ;
        RECT 26.305 33.405 26.655 34.025 ;
        RECT 26.825 33.625 26.995 34.215 ;
        RECT 27.165 33.995 27.335 34.775 ;
        RECT 27.505 34.675 27.675 35.015 ;
        RECT 27.910 34.845 28.240 35.275 ;
        RECT 28.410 34.675 28.580 35.015 ;
        RECT 28.875 34.815 29.245 35.275 ;
        RECT 27.505 34.505 28.580 34.675 ;
        RECT 29.415 34.645 29.585 35.105 ;
        RECT 29.820 34.765 30.690 35.105 ;
        RECT 30.860 34.815 31.110 35.275 ;
        RECT 29.025 34.475 29.585 34.645 ;
        RECT 29.025 34.335 29.195 34.475 ;
        RECT 27.695 34.165 29.195 34.335 ;
        RECT 29.890 34.305 30.350 34.595 ;
        RECT 27.165 33.825 28.855 33.995 ;
        RECT 26.825 33.405 27.180 33.625 ;
        RECT 27.350 33.115 27.520 33.825 ;
        RECT 27.725 33.405 28.515 33.655 ;
        RECT 28.685 33.645 28.855 33.825 ;
        RECT 29.025 33.475 29.195 34.165 ;
        RECT 25.465 32.725 25.795 33.085 ;
        RECT 25.965 32.945 26.460 33.115 ;
        RECT 26.665 32.945 27.520 33.115 ;
        RECT 28.395 32.725 28.725 33.185 ;
        RECT 28.935 33.085 29.195 33.475 ;
        RECT 29.385 34.295 30.350 34.305 ;
        RECT 30.520 34.385 30.690 34.765 ;
        RECT 31.280 34.725 31.450 35.015 ;
        RECT 31.630 34.895 31.960 35.275 ;
        RECT 31.280 34.555 32.080 34.725 ;
        RECT 29.385 34.135 30.060 34.295 ;
        RECT 30.520 34.215 31.740 34.385 ;
        RECT 29.385 33.345 29.595 34.135 ;
        RECT 30.520 34.125 30.690 34.215 ;
        RECT 29.765 33.345 30.115 33.965 ;
        RECT 30.285 33.955 30.690 34.125 ;
        RECT 30.285 33.175 30.455 33.955 ;
        RECT 30.625 33.505 30.845 33.785 ;
        RECT 31.025 33.675 31.565 34.045 ;
        RECT 31.910 33.965 32.080 34.555 ;
        RECT 32.300 34.135 32.605 35.275 ;
        RECT 32.775 34.085 33.030 34.965 ;
        RECT 33.265 34.135 33.475 35.275 ;
        RECT 31.910 33.935 32.650 33.965 ;
        RECT 30.625 33.335 31.155 33.505 ;
        RECT 28.935 32.915 29.285 33.085 ;
        RECT 29.505 32.895 30.455 33.175 ;
        RECT 30.625 32.725 30.815 33.165 ;
        RECT 30.985 33.105 31.155 33.335 ;
        RECT 31.325 33.275 31.565 33.675 ;
        RECT 31.735 33.635 32.650 33.935 ;
        RECT 31.735 33.460 32.060 33.635 ;
        RECT 31.735 33.105 32.055 33.460 ;
        RECT 32.820 33.435 33.030 34.085 ;
        RECT 33.645 34.125 33.975 35.105 ;
        RECT 34.145 34.135 34.375 35.275 ;
        RECT 34.585 34.840 39.930 35.275 ;
        RECT 30.985 32.935 32.055 33.105 ;
        RECT 32.300 32.725 32.605 33.185 ;
        RECT 32.775 32.905 33.030 33.435 ;
        RECT 33.265 32.725 33.475 33.545 ;
        RECT 33.645 33.525 33.895 34.125 ;
        RECT 34.065 33.715 34.395 33.965 ;
        RECT 33.645 32.895 33.975 33.525 ;
        RECT 34.145 32.725 34.375 33.545 ;
        RECT 36.170 33.270 36.510 34.100 ;
        RECT 37.990 33.590 38.340 34.840 ;
        RECT 40.105 34.185 41.315 35.275 ;
        RECT 40.105 33.475 40.625 34.015 ;
        RECT 40.795 33.645 41.315 34.185 ;
        RECT 41.485 34.200 41.755 35.105 ;
        RECT 41.925 34.515 42.255 35.275 ;
        RECT 42.435 34.345 42.605 35.105 ;
        RECT 34.585 32.725 39.930 33.270 ;
        RECT 40.105 32.725 41.315 33.475 ;
        RECT 41.485 33.400 41.655 34.200 ;
        RECT 41.940 34.175 42.605 34.345 ;
        RECT 42.865 34.185 44.075 35.275 ;
        RECT 41.940 34.030 42.110 34.175 ;
        RECT 41.825 33.700 42.110 34.030 ;
        RECT 41.940 33.445 42.110 33.700 ;
        RECT 42.345 33.625 42.675 33.995 ;
        RECT 42.865 33.475 43.385 34.015 ;
        RECT 43.555 33.645 44.075 34.185 ;
        RECT 44.245 34.110 44.535 35.275 ;
        RECT 44.710 34.135 45.045 35.105 ;
        RECT 45.215 34.135 45.385 35.275 ;
        RECT 45.555 34.935 47.585 35.105 ;
        RECT 41.485 32.895 41.745 33.400 ;
        RECT 41.940 33.275 42.605 33.445 ;
        RECT 41.925 32.725 42.255 33.105 ;
        RECT 42.435 32.895 42.605 33.275 ;
        RECT 42.865 32.725 44.075 33.475 ;
        RECT 44.710 33.465 44.880 34.135 ;
        RECT 45.555 33.965 45.725 34.935 ;
        RECT 45.050 33.635 45.305 33.965 ;
        RECT 45.530 33.635 45.725 33.965 ;
        RECT 45.895 34.595 47.020 34.765 ;
        RECT 45.135 33.465 45.305 33.635 ;
        RECT 45.895 33.465 46.065 34.595 ;
        RECT 44.245 32.725 44.535 33.450 ;
        RECT 44.710 32.895 44.965 33.465 ;
        RECT 45.135 33.295 46.065 33.465 ;
        RECT 46.235 34.255 47.245 34.425 ;
        RECT 46.235 33.455 46.405 34.255 ;
        RECT 45.890 33.260 46.065 33.295 ;
        RECT 45.135 32.725 45.465 33.125 ;
        RECT 45.890 32.895 46.420 33.260 ;
        RECT 46.610 33.235 46.885 34.055 ;
        RECT 46.605 33.065 46.885 33.235 ;
        RECT 46.610 32.895 46.885 33.065 ;
        RECT 47.055 32.895 47.245 34.255 ;
        RECT 47.415 34.270 47.585 34.935 ;
        RECT 47.755 34.515 47.925 35.275 ;
        RECT 48.160 34.515 48.675 34.925 ;
        RECT 48.845 34.840 54.190 35.275 ;
        RECT 47.415 34.080 48.165 34.270 ;
        RECT 48.335 33.705 48.675 34.515 ;
        RECT 47.445 33.535 48.675 33.705 ;
        RECT 47.425 32.725 47.935 33.260 ;
        RECT 48.155 32.930 48.400 33.535 ;
        RECT 50.430 33.270 50.770 34.100 ;
        RECT 52.250 33.590 52.600 34.840 ;
        RECT 54.365 34.185 56.955 35.275 ;
        RECT 54.365 33.495 55.575 34.015 ;
        RECT 55.745 33.665 56.955 34.185 ;
        RECT 48.845 32.725 54.190 33.270 ;
        RECT 54.365 32.725 56.955 33.495 ;
        RECT 57.125 32.895 57.385 35.105 ;
        RECT 57.555 34.895 57.885 35.275 ;
        RECT 58.310 34.725 58.480 35.105 ;
        RECT 58.740 34.895 59.070 35.275 ;
        RECT 59.265 34.725 59.435 35.105 ;
        RECT 59.645 34.895 59.975 35.275 ;
        RECT 60.225 34.725 60.415 35.105 ;
        RECT 60.655 34.895 60.985 35.275 ;
        RECT 61.295 34.775 61.555 35.105 ;
        RECT 57.555 34.555 59.505 34.725 ;
        RECT 57.555 33.635 57.725 34.555 ;
        RECT 58.095 33.965 58.290 34.275 ;
        RECT 58.560 33.965 58.745 34.275 ;
        RECT 58.035 33.635 58.290 33.965 ;
        RECT 58.515 33.635 58.745 33.965 ;
        RECT 57.555 32.725 57.885 33.105 ;
        RECT 58.095 33.060 58.290 33.635 ;
        RECT 58.560 33.055 58.745 33.635 ;
        RECT 58.995 33.065 59.165 33.965 ;
        RECT 59.335 33.565 59.505 34.555 ;
        RECT 59.675 34.555 60.415 34.725 ;
        RECT 59.675 34.045 59.845 34.555 ;
        RECT 60.015 34.215 60.595 34.385 ;
        RECT 60.865 34.265 61.215 34.595 ;
        RECT 60.425 34.095 60.595 34.215 ;
        RECT 61.385 34.095 61.555 34.775 ;
        RECT 59.675 33.875 60.245 34.045 ;
        RECT 60.425 33.925 61.555 34.095 ;
        RECT 59.335 33.235 59.885 33.565 ;
        RECT 60.075 33.395 60.245 33.875 ;
        RECT 60.415 33.585 61.035 33.755 ;
        RECT 60.825 33.405 61.035 33.585 ;
        RECT 60.075 33.065 60.475 33.395 ;
        RECT 61.385 33.225 61.555 33.925 ;
        RECT 61.725 33.465 61.985 35.090 ;
        RECT 63.735 34.825 64.065 35.275 ;
        RECT 62.165 34.435 64.775 34.645 ;
        RECT 62.165 33.635 62.385 34.435 ;
        RECT 62.625 33.635 62.925 34.255 ;
        RECT 63.095 33.635 63.425 34.255 ;
        RECT 63.595 33.635 63.915 34.255 ;
        RECT 64.085 33.635 64.435 34.255 ;
        RECT 64.605 33.465 64.775 34.435 ;
        RECT 64.945 34.185 68.455 35.275 ;
        RECT 68.625 34.185 69.835 35.275 ;
        RECT 61.725 33.295 63.565 33.465 ;
        RECT 58.995 32.895 60.475 33.065 ;
        RECT 60.655 32.725 60.985 33.105 ;
        RECT 61.295 32.895 61.555 33.225 ;
        RECT 61.995 32.725 62.325 33.120 ;
        RECT 62.495 32.940 62.695 33.295 ;
        RECT 62.865 32.725 63.195 33.125 ;
        RECT 63.365 32.950 63.565 33.295 ;
        RECT 63.735 32.725 64.065 33.465 ;
        RECT 64.300 33.295 64.775 33.465 ;
        RECT 64.945 33.495 66.595 34.015 ;
        RECT 66.765 33.665 68.455 34.185 ;
        RECT 64.300 33.045 64.470 33.295 ;
        RECT 64.945 32.725 68.455 33.495 ;
        RECT 68.625 33.475 69.145 34.015 ;
        RECT 69.315 33.645 69.835 34.185 ;
        RECT 70.005 34.110 70.295 35.275 ;
        RECT 70.465 34.840 75.810 35.275 ;
        RECT 68.625 32.725 69.835 33.475 ;
        RECT 70.005 32.725 70.295 33.450 ;
        RECT 72.050 33.270 72.390 34.100 ;
        RECT 73.870 33.590 74.220 34.840 ;
        RECT 76.445 34.515 76.960 34.925 ;
        RECT 77.195 34.515 77.365 35.275 ;
        RECT 77.535 34.935 79.565 35.105 ;
        RECT 76.445 33.705 76.785 34.515 ;
        RECT 77.535 34.270 77.705 34.935 ;
        RECT 78.100 34.595 79.225 34.765 ;
        RECT 76.955 34.080 77.705 34.270 ;
        RECT 77.875 34.255 78.885 34.425 ;
        RECT 76.445 33.535 77.675 33.705 ;
        RECT 70.465 32.725 75.810 33.270 ;
        RECT 76.720 32.930 76.965 33.535 ;
        RECT 77.185 32.725 77.695 33.260 ;
        RECT 77.875 32.895 78.065 34.255 ;
        RECT 78.235 33.915 78.510 34.055 ;
        RECT 78.235 33.745 78.515 33.915 ;
        RECT 78.235 32.895 78.510 33.745 ;
        RECT 78.715 33.455 78.885 34.255 ;
        RECT 79.055 33.465 79.225 34.595 ;
        RECT 79.395 33.965 79.565 34.935 ;
        RECT 79.735 34.135 79.905 35.275 ;
        RECT 80.075 34.135 80.410 35.105 ;
        RECT 80.625 34.135 80.855 35.275 ;
        RECT 79.395 33.635 79.590 33.965 ;
        RECT 79.815 33.635 80.070 33.965 ;
        RECT 79.815 33.465 79.985 33.635 ;
        RECT 80.240 33.465 80.410 34.135 ;
        RECT 81.025 34.125 81.355 35.105 ;
        RECT 81.525 34.135 81.735 35.275 ;
        RECT 81.965 34.840 87.310 35.275 ;
        RECT 80.605 33.715 80.935 33.965 ;
        RECT 79.055 33.295 79.985 33.465 ;
        RECT 79.055 33.260 79.230 33.295 ;
        RECT 78.700 32.895 79.230 33.260 ;
        RECT 79.655 32.725 79.985 33.125 ;
        RECT 80.155 32.895 80.410 33.465 ;
        RECT 80.625 32.725 80.855 33.545 ;
        RECT 81.105 33.525 81.355 34.125 ;
        RECT 81.025 32.895 81.355 33.525 ;
        RECT 81.525 32.725 81.735 33.545 ;
        RECT 83.550 33.270 83.890 34.100 ;
        RECT 85.370 33.590 85.720 34.840 ;
        RECT 87.485 34.185 88.695 35.275 ;
        RECT 87.485 33.475 88.005 34.015 ;
        RECT 88.175 33.645 88.695 34.185 ;
        RECT 88.870 34.135 89.205 35.105 ;
        RECT 89.375 34.135 89.545 35.275 ;
        RECT 89.715 34.935 91.745 35.105 ;
        RECT 81.965 32.725 87.310 33.270 ;
        RECT 87.485 32.725 88.695 33.475 ;
        RECT 88.870 33.465 89.040 34.135 ;
        RECT 89.715 33.965 89.885 34.935 ;
        RECT 89.210 33.635 89.465 33.965 ;
        RECT 89.690 33.635 89.885 33.965 ;
        RECT 90.055 34.595 91.180 34.765 ;
        RECT 89.295 33.465 89.465 33.635 ;
        RECT 90.055 33.465 90.225 34.595 ;
        RECT 88.870 32.895 89.125 33.465 ;
        RECT 89.295 33.295 90.225 33.465 ;
        RECT 90.395 34.255 91.405 34.425 ;
        RECT 90.395 33.455 90.565 34.255 ;
        RECT 90.770 33.575 91.045 34.055 ;
        RECT 90.765 33.405 91.045 33.575 ;
        RECT 90.050 33.260 90.225 33.295 ;
        RECT 89.295 32.725 89.625 33.125 ;
        RECT 90.050 32.895 90.580 33.260 ;
        RECT 90.770 32.895 91.045 33.405 ;
        RECT 91.215 32.895 91.405 34.255 ;
        RECT 91.575 34.270 91.745 34.935 ;
        RECT 91.915 34.515 92.085 35.275 ;
        RECT 92.320 34.515 92.835 34.925 ;
        RECT 91.575 34.080 92.325 34.270 ;
        RECT 92.495 33.705 92.835 34.515 ;
        RECT 91.605 33.535 92.835 33.705 ;
        RECT 93.465 34.200 93.735 35.105 ;
        RECT 93.905 34.515 94.235 35.275 ;
        RECT 94.415 34.345 94.585 35.105 ;
        RECT 91.585 32.725 92.095 33.260 ;
        RECT 92.315 32.930 92.560 33.535 ;
        RECT 93.465 33.400 93.635 34.200 ;
        RECT 93.920 34.175 94.585 34.345 ;
        RECT 93.920 34.030 94.090 34.175 ;
        RECT 95.765 34.110 96.055 35.275 ;
        RECT 96.230 34.135 96.565 35.105 ;
        RECT 96.735 34.135 96.905 35.275 ;
        RECT 97.075 34.935 99.105 35.105 ;
        RECT 93.805 33.700 94.090 34.030 ;
        RECT 93.920 33.445 94.090 33.700 ;
        RECT 94.325 33.625 94.655 33.995 ;
        RECT 96.230 33.465 96.400 34.135 ;
        RECT 97.075 33.965 97.245 34.935 ;
        RECT 96.570 33.635 96.825 33.965 ;
        RECT 97.050 33.635 97.245 33.965 ;
        RECT 97.415 34.595 98.540 34.765 ;
        RECT 96.655 33.465 96.825 33.635 ;
        RECT 97.415 33.465 97.585 34.595 ;
        RECT 93.465 32.895 93.725 33.400 ;
        RECT 93.920 33.275 94.585 33.445 ;
        RECT 93.905 32.725 94.235 33.105 ;
        RECT 94.415 32.895 94.585 33.275 ;
        RECT 95.765 32.725 96.055 33.450 ;
        RECT 96.230 32.895 96.485 33.465 ;
        RECT 96.655 33.295 97.585 33.465 ;
        RECT 97.755 34.255 98.765 34.425 ;
        RECT 97.755 33.455 97.925 34.255 ;
        RECT 98.130 33.915 98.405 34.055 ;
        RECT 98.125 33.745 98.405 33.915 ;
        RECT 97.410 33.260 97.585 33.295 ;
        RECT 96.655 32.725 96.985 33.125 ;
        RECT 97.410 32.895 97.940 33.260 ;
        RECT 98.130 32.895 98.405 33.745 ;
        RECT 98.575 32.895 98.765 34.255 ;
        RECT 98.935 34.270 99.105 34.935 ;
        RECT 99.275 34.515 99.445 35.275 ;
        RECT 99.680 34.515 100.195 34.925 ;
        RECT 100.365 34.840 105.710 35.275 ;
        RECT 105.885 34.840 111.230 35.275 ;
        RECT 98.935 34.080 99.685 34.270 ;
        RECT 99.855 33.705 100.195 34.515 ;
        RECT 98.965 33.535 100.195 33.705 ;
        RECT 98.945 32.725 99.455 33.260 ;
        RECT 99.675 32.930 99.920 33.535 ;
        RECT 101.950 33.270 102.290 34.100 ;
        RECT 103.770 33.590 104.120 34.840 ;
        RECT 107.470 33.270 107.810 34.100 ;
        RECT 109.290 33.590 109.640 34.840 ;
        RECT 112.325 34.185 113.535 35.275 ;
        RECT 112.325 33.645 112.845 34.185 ;
        RECT 113.015 33.475 113.535 34.015 ;
        RECT 100.365 32.725 105.710 33.270 ;
        RECT 105.885 32.725 111.230 33.270 ;
        RECT 112.325 32.725 113.535 33.475 ;
        RECT 5.520 32.555 113.620 32.725 ;
        RECT 5.605 31.805 6.815 32.555 ;
        RECT 6.985 32.010 12.330 32.555 ;
        RECT 5.605 31.265 6.125 31.805 ;
        RECT 6.295 31.095 6.815 31.635 ;
        RECT 8.570 31.180 8.910 32.010 ;
        RECT 12.505 31.785 16.015 32.555 ;
        RECT 16.185 31.805 17.395 32.555 ;
        RECT 5.605 30.005 6.815 31.095 ;
        RECT 10.390 30.440 10.740 31.690 ;
        RECT 12.505 31.265 14.155 31.785 ;
        RECT 14.325 31.095 16.015 31.615 ;
        RECT 16.185 31.265 16.705 31.805 ;
        RECT 17.840 31.745 18.085 32.350 ;
        RECT 18.305 32.020 18.815 32.555 ;
        RECT 16.875 31.095 17.395 31.635 ;
        RECT 6.985 30.005 12.330 30.440 ;
        RECT 12.505 30.005 16.015 31.095 ;
        RECT 16.185 30.005 17.395 31.095 ;
        RECT 17.565 31.575 18.795 31.745 ;
        RECT 17.565 30.765 17.905 31.575 ;
        RECT 18.075 31.010 18.825 31.200 ;
        RECT 17.565 30.355 18.080 30.765 ;
        RECT 18.315 30.005 18.485 30.765 ;
        RECT 18.655 30.345 18.825 31.010 ;
        RECT 18.995 31.025 19.185 32.385 ;
        RECT 19.355 31.535 19.630 32.385 ;
        RECT 19.820 32.020 20.350 32.385 ;
        RECT 20.775 32.155 21.105 32.555 ;
        RECT 20.175 31.985 20.350 32.020 ;
        RECT 19.355 31.365 19.635 31.535 ;
        RECT 19.355 31.225 19.630 31.365 ;
        RECT 19.835 31.025 20.005 31.825 ;
        RECT 18.995 30.855 20.005 31.025 ;
        RECT 20.175 31.815 21.105 31.985 ;
        RECT 21.275 31.815 21.530 32.385 ;
        RECT 20.175 30.685 20.345 31.815 ;
        RECT 20.935 31.645 21.105 31.815 ;
        RECT 19.220 30.515 20.345 30.685 ;
        RECT 20.515 31.315 20.710 31.645 ;
        RECT 20.935 31.315 21.190 31.645 ;
        RECT 20.515 30.345 20.685 31.315 ;
        RECT 21.360 31.145 21.530 31.815 ;
        RECT 21.705 31.785 24.295 32.555 ;
        RECT 24.555 32.005 24.725 32.385 ;
        RECT 24.905 32.175 25.235 32.555 ;
        RECT 24.555 31.835 25.220 32.005 ;
        RECT 25.415 31.880 25.675 32.385 ;
        RECT 25.845 32.010 31.190 32.555 ;
        RECT 21.705 31.265 22.915 31.785 ;
        RECT 18.655 30.175 20.685 30.345 ;
        RECT 20.855 30.005 21.025 31.145 ;
        RECT 21.195 30.175 21.530 31.145 ;
        RECT 23.085 31.095 24.295 31.615 ;
        RECT 24.485 31.285 24.815 31.655 ;
        RECT 25.050 31.580 25.220 31.835 ;
        RECT 25.050 31.250 25.335 31.580 ;
        RECT 25.050 31.105 25.220 31.250 ;
        RECT 21.705 30.005 24.295 31.095 ;
        RECT 24.555 30.935 25.220 31.105 ;
        RECT 25.505 31.080 25.675 31.880 ;
        RECT 27.430 31.180 27.770 32.010 ;
        RECT 31.365 31.830 31.655 32.555 ;
        RECT 31.825 32.010 37.170 32.555 ;
        RECT 24.555 30.175 24.725 30.935 ;
        RECT 24.905 30.005 25.235 30.765 ;
        RECT 25.405 30.175 25.675 31.080 ;
        RECT 29.250 30.440 29.600 31.690 ;
        RECT 33.410 31.180 33.750 32.010 ;
        RECT 37.345 31.785 39.015 32.555 ;
        RECT 39.275 32.005 39.445 32.295 ;
        RECT 39.615 32.175 39.945 32.555 ;
        RECT 39.275 31.835 39.940 32.005 ;
        RECT 25.845 30.005 31.190 30.440 ;
        RECT 31.365 30.005 31.655 31.170 ;
        RECT 35.230 30.440 35.580 31.690 ;
        RECT 37.345 31.265 38.095 31.785 ;
        RECT 38.265 31.095 39.015 31.615 ;
        RECT 31.825 30.005 37.170 30.440 ;
        RECT 37.345 30.005 39.015 31.095 ;
        RECT 39.190 31.015 39.540 31.665 ;
        RECT 39.710 30.845 39.940 31.835 ;
        RECT 39.275 30.675 39.940 30.845 ;
        RECT 39.275 30.175 39.445 30.675 ;
        RECT 39.615 30.005 39.945 30.505 ;
        RECT 40.115 30.175 40.340 32.295 ;
        RECT 40.555 32.175 40.885 32.555 ;
        RECT 41.055 32.005 41.225 32.335 ;
        RECT 41.525 32.175 42.540 32.375 ;
        RECT 40.530 31.815 41.225 32.005 ;
        RECT 40.530 30.845 40.700 31.815 ;
        RECT 40.870 31.015 41.280 31.635 ;
        RECT 41.450 31.065 41.670 31.935 ;
        RECT 41.850 31.625 42.200 31.995 ;
        RECT 42.370 31.445 42.540 32.175 ;
        RECT 42.710 32.115 43.120 32.555 ;
        RECT 43.410 31.915 43.660 32.345 ;
        RECT 43.860 32.095 44.180 32.555 ;
        RECT 44.740 32.165 45.590 32.335 ;
        RECT 42.710 31.575 43.120 31.905 ;
        RECT 43.410 31.575 43.830 31.915 ;
        RECT 42.120 31.405 42.540 31.445 ;
        RECT 42.120 31.235 43.470 31.405 ;
        RECT 40.530 30.675 41.225 30.845 ;
        RECT 41.450 30.685 41.950 31.065 ;
        RECT 40.555 30.005 40.885 30.505 ;
        RECT 41.055 30.175 41.225 30.675 ;
        RECT 42.120 30.390 42.290 31.235 ;
        RECT 43.220 31.075 43.470 31.235 ;
        RECT 42.460 30.805 42.710 31.065 ;
        RECT 43.640 30.805 43.830 31.575 ;
        RECT 42.460 30.555 43.830 30.805 ;
        RECT 44.000 31.745 45.250 31.915 ;
        RECT 44.000 30.985 44.170 31.745 ;
        RECT 44.920 31.625 45.250 31.745 ;
        RECT 44.340 31.165 44.520 31.575 ;
        RECT 45.420 31.405 45.590 32.165 ;
        RECT 45.790 32.075 46.450 32.555 ;
        RECT 46.630 31.960 46.950 32.290 ;
        RECT 45.780 31.635 46.440 31.905 ;
        RECT 45.780 31.575 46.110 31.635 ;
        RECT 46.260 31.405 46.590 31.465 ;
        RECT 44.690 31.235 46.590 31.405 ;
        RECT 44.000 30.675 44.520 30.985 ;
        RECT 44.690 30.725 44.860 31.235 ;
        RECT 46.760 31.065 46.950 31.960 ;
        RECT 45.030 30.895 46.950 31.065 ;
        RECT 46.630 30.875 46.950 30.895 ;
        RECT 47.150 31.645 47.400 32.295 ;
        RECT 47.580 32.095 47.865 32.555 ;
        RECT 48.045 32.215 48.300 32.375 ;
        RECT 48.045 32.045 48.385 32.215 ;
        RECT 48.045 31.845 48.300 32.045 ;
        RECT 47.150 31.315 47.950 31.645 ;
        RECT 44.690 30.555 45.900 30.725 ;
        RECT 41.460 30.220 42.290 30.390 ;
        RECT 42.530 30.005 42.910 30.385 ;
        RECT 43.090 30.265 43.260 30.555 ;
        RECT 44.690 30.475 44.860 30.555 ;
        RECT 43.430 30.005 43.760 30.385 ;
        RECT 44.230 30.225 44.860 30.475 ;
        RECT 45.040 30.005 45.460 30.385 ;
        RECT 45.660 30.265 45.900 30.555 ;
        RECT 46.130 30.005 46.460 30.695 ;
        RECT 46.630 30.265 46.800 30.875 ;
        RECT 47.150 30.725 47.400 31.315 ;
        RECT 48.120 30.985 48.300 31.845 ;
        RECT 47.070 30.215 47.400 30.725 ;
        RECT 47.580 30.005 47.865 30.805 ;
        RECT 48.045 30.315 48.300 30.985 ;
        RECT 48.850 31.815 49.105 32.385 ;
        RECT 49.275 32.155 49.605 32.555 ;
        RECT 50.030 32.020 50.560 32.385 ;
        RECT 50.750 32.215 51.025 32.385 ;
        RECT 50.745 32.045 51.025 32.215 ;
        RECT 50.030 31.985 50.205 32.020 ;
        RECT 49.275 31.815 50.205 31.985 ;
        RECT 48.850 31.145 49.020 31.815 ;
        RECT 49.275 31.645 49.445 31.815 ;
        RECT 49.190 31.315 49.445 31.645 ;
        RECT 49.670 31.315 49.865 31.645 ;
        RECT 48.850 30.175 49.185 31.145 ;
        RECT 49.355 30.005 49.525 31.145 ;
        RECT 49.695 30.345 49.865 31.315 ;
        RECT 50.035 30.685 50.205 31.815 ;
        RECT 50.375 31.025 50.545 31.825 ;
        RECT 50.750 31.225 51.025 32.045 ;
        RECT 51.195 31.025 51.385 32.385 ;
        RECT 51.565 32.020 52.075 32.555 ;
        RECT 52.295 31.745 52.540 32.350 ;
        RECT 51.585 31.575 52.815 31.745 ;
        RECT 53.025 31.735 53.255 32.555 ;
        RECT 53.425 31.755 53.755 32.385 ;
        RECT 50.375 30.855 51.385 31.025 ;
        RECT 51.555 31.010 52.305 31.200 ;
        RECT 50.035 30.515 51.160 30.685 ;
        RECT 51.555 30.345 51.725 31.010 ;
        RECT 52.475 30.765 52.815 31.575 ;
        RECT 53.005 31.315 53.335 31.565 ;
        RECT 53.505 31.155 53.755 31.755 ;
        RECT 53.925 31.735 54.135 32.555 ;
        RECT 54.365 31.785 56.955 32.555 ;
        RECT 57.125 31.830 57.415 32.555 ;
        RECT 57.890 31.985 58.060 32.235 ;
        RECT 57.585 31.815 58.060 31.985 ;
        RECT 58.295 31.815 58.625 32.555 ;
        RECT 58.795 31.985 58.995 32.330 ;
        RECT 59.165 32.155 59.495 32.555 ;
        RECT 59.665 31.985 59.865 32.340 ;
        RECT 60.035 32.160 60.365 32.555 ;
        RECT 60.805 32.010 66.150 32.555 ;
        RECT 58.795 31.815 60.635 31.985 ;
        RECT 54.365 31.265 55.575 31.785 ;
        RECT 49.695 30.175 51.725 30.345 ;
        RECT 51.895 30.005 52.065 30.765 ;
        RECT 52.300 30.355 52.815 30.765 ;
        RECT 53.025 30.005 53.255 31.145 ;
        RECT 53.425 30.175 53.755 31.155 ;
        RECT 53.925 30.005 54.135 31.145 ;
        RECT 55.745 31.095 56.955 31.615 ;
        RECT 54.365 30.005 56.955 31.095 ;
        RECT 57.125 30.005 57.415 31.170 ;
        RECT 57.585 30.845 57.755 31.815 ;
        RECT 57.925 31.025 58.275 31.645 ;
        RECT 58.445 31.025 58.765 31.645 ;
        RECT 58.935 31.025 59.265 31.645 ;
        RECT 59.435 31.025 59.735 31.645 ;
        RECT 59.975 30.845 60.195 31.645 ;
        RECT 57.585 30.635 60.195 30.845 ;
        RECT 58.295 30.005 58.625 30.455 ;
        RECT 60.375 30.190 60.635 31.815 ;
        RECT 62.390 31.180 62.730 32.010 ;
        RECT 66.325 31.785 68.915 32.555 ;
        RECT 69.550 31.815 69.805 32.385 ;
        RECT 69.975 32.155 70.305 32.555 ;
        RECT 70.730 32.020 71.260 32.385 ;
        RECT 70.730 31.985 70.905 32.020 ;
        RECT 69.975 31.815 70.905 31.985 ;
        RECT 64.210 30.440 64.560 31.690 ;
        RECT 66.325 31.265 67.535 31.785 ;
        RECT 67.705 31.095 68.915 31.615 ;
        RECT 60.805 30.005 66.150 30.440 ;
        RECT 66.325 30.005 68.915 31.095 ;
        RECT 69.550 31.145 69.720 31.815 ;
        RECT 69.975 31.645 70.145 31.815 ;
        RECT 69.890 31.315 70.145 31.645 ;
        RECT 70.370 31.315 70.565 31.645 ;
        RECT 69.550 30.175 69.885 31.145 ;
        RECT 70.055 30.005 70.225 31.145 ;
        RECT 70.395 30.345 70.565 31.315 ;
        RECT 70.735 30.685 70.905 31.815 ;
        RECT 71.075 31.025 71.245 31.825 ;
        RECT 71.450 31.535 71.725 32.385 ;
        RECT 71.445 31.365 71.725 31.535 ;
        RECT 71.450 31.225 71.725 31.365 ;
        RECT 71.895 31.025 72.085 32.385 ;
        RECT 72.265 32.020 72.775 32.555 ;
        RECT 72.995 31.745 73.240 32.350 ;
        RECT 73.690 32.005 73.945 32.295 ;
        RECT 74.115 32.175 74.445 32.555 ;
        RECT 73.690 31.835 74.440 32.005 ;
        RECT 72.285 31.575 73.515 31.745 ;
        RECT 71.075 30.855 72.085 31.025 ;
        RECT 72.255 31.010 73.005 31.200 ;
        RECT 70.735 30.515 71.860 30.685 ;
        RECT 72.255 30.345 72.425 31.010 ;
        RECT 73.175 30.765 73.515 31.575 ;
        RECT 73.690 31.015 74.040 31.665 ;
        RECT 74.210 30.845 74.440 31.835 ;
        RECT 70.395 30.175 72.425 30.345 ;
        RECT 72.595 30.005 72.765 30.765 ;
        RECT 73.000 30.355 73.515 30.765 ;
        RECT 73.690 30.675 74.440 30.845 ;
        RECT 73.690 30.175 73.945 30.675 ;
        RECT 74.115 30.005 74.445 30.505 ;
        RECT 74.615 30.175 74.785 32.295 ;
        RECT 75.145 32.195 75.475 32.555 ;
        RECT 75.645 32.165 76.140 32.335 ;
        RECT 76.345 32.165 77.200 32.335 ;
        RECT 75.015 30.975 75.475 32.025 ;
        RECT 74.955 30.190 75.280 30.975 ;
        RECT 75.645 30.805 75.815 32.165 ;
        RECT 75.985 31.255 76.335 31.875 ;
        RECT 76.505 31.655 76.860 31.875 ;
        RECT 76.505 31.065 76.675 31.655 ;
        RECT 77.030 31.455 77.200 32.165 ;
        RECT 78.075 32.095 78.405 32.555 ;
        RECT 78.615 32.195 78.965 32.365 ;
        RECT 77.405 31.625 78.195 31.875 ;
        RECT 78.615 31.805 78.875 32.195 ;
        RECT 79.185 32.105 80.135 32.385 ;
        RECT 80.305 32.115 80.495 32.555 ;
        RECT 80.665 32.175 81.735 32.345 ;
        RECT 78.365 31.455 78.535 31.635 ;
        RECT 75.645 30.635 76.040 30.805 ;
        RECT 76.210 30.675 76.675 31.065 ;
        RECT 76.845 31.285 78.535 31.455 ;
        RECT 75.870 30.505 76.040 30.635 ;
        RECT 76.845 30.505 77.015 31.285 ;
        RECT 78.705 31.115 78.875 31.805 ;
        RECT 77.375 30.945 78.875 31.115 ;
        RECT 79.065 31.145 79.275 31.935 ;
        RECT 79.445 31.315 79.795 31.935 ;
        RECT 79.965 31.325 80.135 32.105 ;
        RECT 80.665 31.945 80.835 32.175 ;
        RECT 80.305 31.775 80.835 31.945 ;
        RECT 80.305 31.495 80.525 31.775 ;
        RECT 81.005 31.605 81.245 32.005 ;
        RECT 79.965 31.155 80.370 31.325 ;
        RECT 80.705 31.235 81.245 31.605 ;
        RECT 81.415 31.820 81.735 32.175 ;
        RECT 81.980 32.095 82.285 32.555 ;
        RECT 82.455 31.845 82.710 32.375 ;
        RECT 81.415 31.645 81.740 31.820 ;
        RECT 81.415 31.345 82.330 31.645 ;
        RECT 81.590 31.315 82.330 31.345 ;
        RECT 79.065 30.985 79.740 31.145 ;
        RECT 80.200 31.065 80.370 31.155 ;
        RECT 79.065 30.975 80.030 30.985 ;
        RECT 78.705 30.805 78.875 30.945 ;
        RECT 75.450 30.005 75.700 30.465 ;
        RECT 75.870 30.175 76.120 30.505 ;
        RECT 76.335 30.175 77.015 30.505 ;
        RECT 77.185 30.605 78.260 30.775 ;
        RECT 78.705 30.635 79.265 30.805 ;
        RECT 79.570 30.685 80.030 30.975 ;
        RECT 80.200 30.895 81.420 31.065 ;
        RECT 77.185 30.265 77.355 30.605 ;
        RECT 77.590 30.005 77.920 30.435 ;
        RECT 78.090 30.265 78.260 30.605 ;
        RECT 78.555 30.005 78.925 30.465 ;
        RECT 79.095 30.175 79.265 30.635 ;
        RECT 80.200 30.515 80.370 30.895 ;
        RECT 81.590 30.725 81.760 31.315 ;
        RECT 82.500 31.195 82.710 31.845 ;
        RECT 82.885 31.830 83.175 32.555 ;
        RECT 79.500 30.175 80.370 30.515 ;
        RECT 80.960 30.555 81.760 30.725 ;
        RECT 80.540 30.005 80.790 30.465 ;
        RECT 80.960 30.265 81.130 30.555 ;
        RECT 81.310 30.005 81.640 30.385 ;
        RECT 81.980 30.005 82.285 31.145 ;
        RECT 82.455 30.315 82.710 31.195 ;
        RECT 84.270 31.815 84.525 32.385 ;
        RECT 84.695 32.155 85.025 32.555 ;
        RECT 85.450 32.020 85.980 32.385 ;
        RECT 86.170 32.215 86.445 32.385 ;
        RECT 86.165 32.045 86.445 32.215 ;
        RECT 85.450 31.985 85.625 32.020 ;
        RECT 84.695 31.815 85.625 31.985 ;
        RECT 82.885 30.005 83.175 31.170 ;
        RECT 84.270 31.145 84.440 31.815 ;
        RECT 84.695 31.645 84.865 31.815 ;
        RECT 84.610 31.315 84.865 31.645 ;
        RECT 85.090 31.315 85.285 31.645 ;
        RECT 84.270 30.175 84.605 31.145 ;
        RECT 84.775 30.005 84.945 31.145 ;
        RECT 85.115 30.345 85.285 31.315 ;
        RECT 85.455 30.685 85.625 31.815 ;
        RECT 85.795 31.025 85.965 31.825 ;
        RECT 86.170 31.225 86.445 32.045 ;
        RECT 86.615 31.025 86.805 32.385 ;
        RECT 86.985 32.020 87.495 32.555 ;
        RECT 87.715 31.745 87.960 32.350 ;
        RECT 88.405 31.880 88.665 32.385 ;
        RECT 88.845 32.175 89.175 32.555 ;
        RECT 89.355 32.005 89.525 32.385 ;
        RECT 87.005 31.575 88.235 31.745 ;
        RECT 85.795 30.855 86.805 31.025 ;
        RECT 86.975 31.010 87.725 31.200 ;
        RECT 85.455 30.515 86.580 30.685 ;
        RECT 86.975 30.345 87.145 31.010 ;
        RECT 87.895 30.765 88.235 31.575 ;
        RECT 85.115 30.175 87.145 30.345 ;
        RECT 87.315 30.005 87.485 30.765 ;
        RECT 87.720 30.355 88.235 30.765 ;
        RECT 88.405 31.080 88.575 31.880 ;
        RECT 88.860 31.835 89.525 32.005 ;
        RECT 88.860 31.580 89.030 31.835 ;
        RECT 90.745 31.735 90.975 32.555 ;
        RECT 91.145 31.755 91.475 32.385 ;
        RECT 88.745 31.250 89.030 31.580 ;
        RECT 89.265 31.285 89.595 31.655 ;
        RECT 90.725 31.315 91.055 31.565 ;
        RECT 88.860 31.105 89.030 31.250 ;
        RECT 91.225 31.155 91.475 31.755 ;
        RECT 91.645 31.735 91.855 32.555 ;
        RECT 92.090 32.005 92.345 32.295 ;
        RECT 92.515 32.175 92.845 32.555 ;
        RECT 92.090 31.835 92.840 32.005 ;
        RECT 88.405 30.175 88.675 31.080 ;
        RECT 88.860 30.935 89.525 31.105 ;
        RECT 88.845 30.005 89.175 30.765 ;
        RECT 89.355 30.175 89.525 30.935 ;
        RECT 90.745 30.005 90.975 31.145 ;
        RECT 91.145 30.175 91.475 31.155 ;
        RECT 91.645 30.005 91.855 31.145 ;
        RECT 92.090 31.015 92.440 31.665 ;
        RECT 92.610 30.845 92.840 31.835 ;
        RECT 92.090 30.675 92.840 30.845 ;
        RECT 92.090 30.175 92.345 30.675 ;
        RECT 92.515 30.005 92.845 30.505 ;
        RECT 93.015 30.175 93.185 32.295 ;
        RECT 93.545 32.195 93.875 32.555 ;
        RECT 94.045 32.165 94.540 32.335 ;
        RECT 94.745 32.165 95.600 32.335 ;
        RECT 93.415 30.975 93.875 32.025 ;
        RECT 93.355 30.190 93.680 30.975 ;
        RECT 94.045 30.805 94.215 32.165 ;
        RECT 94.385 31.255 94.735 31.875 ;
        RECT 94.905 31.655 95.260 31.875 ;
        RECT 94.905 31.065 95.075 31.655 ;
        RECT 95.430 31.455 95.600 32.165 ;
        RECT 96.475 32.095 96.805 32.555 ;
        RECT 97.015 32.195 97.365 32.365 ;
        RECT 95.805 31.625 96.595 31.875 ;
        RECT 97.015 31.805 97.275 32.195 ;
        RECT 97.585 32.105 98.535 32.385 ;
        RECT 98.705 32.115 98.895 32.555 ;
        RECT 99.065 32.175 100.135 32.345 ;
        RECT 96.765 31.455 96.935 31.635 ;
        RECT 94.045 30.635 94.440 30.805 ;
        RECT 94.610 30.675 95.075 31.065 ;
        RECT 95.245 31.285 96.935 31.455 ;
        RECT 94.270 30.505 94.440 30.635 ;
        RECT 95.245 30.505 95.415 31.285 ;
        RECT 97.105 31.115 97.275 31.805 ;
        RECT 95.775 30.945 97.275 31.115 ;
        RECT 97.465 31.145 97.675 31.935 ;
        RECT 97.845 31.315 98.195 31.935 ;
        RECT 98.365 31.325 98.535 32.105 ;
        RECT 99.065 31.945 99.235 32.175 ;
        RECT 98.705 31.775 99.235 31.945 ;
        RECT 98.705 31.495 98.925 31.775 ;
        RECT 99.405 31.605 99.645 32.005 ;
        RECT 98.365 31.155 98.770 31.325 ;
        RECT 99.105 31.235 99.645 31.605 ;
        RECT 99.815 31.820 100.135 32.175 ;
        RECT 100.380 32.095 100.685 32.555 ;
        RECT 100.855 31.845 101.110 32.375 ;
        RECT 99.815 31.645 100.140 31.820 ;
        RECT 99.815 31.345 100.730 31.645 ;
        RECT 99.990 31.315 100.730 31.345 ;
        RECT 97.465 30.985 98.140 31.145 ;
        RECT 98.600 31.065 98.770 31.155 ;
        RECT 97.465 30.975 98.430 30.985 ;
        RECT 97.105 30.805 97.275 30.945 ;
        RECT 93.850 30.005 94.100 30.465 ;
        RECT 94.270 30.175 94.520 30.505 ;
        RECT 94.735 30.175 95.415 30.505 ;
        RECT 95.585 30.605 96.660 30.775 ;
        RECT 97.105 30.635 97.665 30.805 ;
        RECT 97.970 30.685 98.430 30.975 ;
        RECT 98.600 30.895 99.820 31.065 ;
        RECT 95.585 30.265 95.755 30.605 ;
        RECT 95.990 30.005 96.320 30.435 ;
        RECT 96.490 30.265 96.660 30.605 ;
        RECT 96.955 30.005 97.325 30.465 ;
        RECT 97.495 30.175 97.665 30.635 ;
        RECT 98.600 30.515 98.770 30.895 ;
        RECT 99.990 30.725 100.160 31.315 ;
        RECT 100.900 31.195 101.110 31.845 ;
        RECT 101.345 31.735 101.555 32.555 ;
        RECT 101.725 31.755 102.055 32.385 ;
        RECT 97.900 30.175 98.770 30.515 ;
        RECT 99.360 30.555 100.160 30.725 ;
        RECT 98.940 30.005 99.190 30.465 ;
        RECT 99.360 30.265 99.530 30.555 ;
        RECT 99.710 30.005 100.040 30.385 ;
        RECT 100.380 30.005 100.685 31.145 ;
        RECT 100.855 30.315 101.110 31.195 ;
        RECT 101.725 31.155 101.975 31.755 ;
        RECT 102.225 31.735 102.455 32.555 ;
        RECT 102.665 32.010 108.010 32.555 ;
        RECT 102.145 31.315 102.475 31.565 ;
        RECT 104.250 31.180 104.590 32.010 ;
        RECT 108.645 31.830 108.935 32.555 ;
        RECT 109.105 31.785 111.695 32.555 ;
        RECT 112.325 31.805 113.535 32.555 ;
        RECT 101.345 30.005 101.555 31.145 ;
        RECT 101.725 30.175 102.055 31.155 ;
        RECT 102.225 30.005 102.455 31.145 ;
        RECT 106.070 30.440 106.420 31.690 ;
        RECT 109.105 31.265 110.315 31.785 ;
        RECT 102.665 30.005 108.010 30.440 ;
        RECT 108.645 30.005 108.935 31.170 ;
        RECT 110.485 31.095 111.695 31.615 ;
        RECT 109.105 30.005 111.695 31.095 ;
        RECT 112.325 31.095 112.845 31.635 ;
        RECT 113.015 31.265 113.535 31.805 ;
        RECT 112.325 30.005 113.535 31.095 ;
        RECT 5.520 29.835 113.620 30.005 ;
        RECT 5.605 28.745 6.815 29.835 ;
        RECT 6.985 28.745 8.655 29.835 ;
        RECT 9.290 29.165 9.545 29.665 ;
        RECT 9.715 29.335 10.045 29.835 ;
        RECT 9.290 28.995 10.040 29.165 ;
        RECT 5.605 28.035 6.125 28.575 ;
        RECT 6.295 28.205 6.815 28.745 ;
        RECT 6.985 28.055 7.735 28.575 ;
        RECT 7.905 28.225 8.655 28.745 ;
        RECT 9.290 28.175 9.640 28.825 ;
        RECT 5.605 27.285 6.815 28.035 ;
        RECT 6.985 27.285 8.655 28.055 ;
        RECT 9.810 28.005 10.040 28.995 ;
        RECT 9.290 27.835 10.040 28.005 ;
        RECT 9.290 27.545 9.545 27.835 ;
        RECT 9.715 27.285 10.045 27.665 ;
        RECT 10.215 27.545 10.385 29.665 ;
        RECT 10.555 28.865 10.880 29.650 ;
        RECT 11.050 29.375 11.300 29.835 ;
        RECT 11.470 29.335 11.720 29.665 ;
        RECT 11.935 29.335 12.615 29.665 ;
        RECT 11.470 29.205 11.640 29.335 ;
        RECT 11.245 29.035 11.640 29.205 ;
        RECT 10.615 27.815 11.075 28.865 ;
        RECT 11.245 27.675 11.415 29.035 ;
        RECT 11.810 28.775 12.275 29.165 ;
        RECT 11.585 27.965 11.935 28.585 ;
        RECT 12.105 28.185 12.275 28.775 ;
        RECT 12.445 28.555 12.615 29.335 ;
        RECT 12.785 29.235 12.955 29.575 ;
        RECT 13.190 29.405 13.520 29.835 ;
        RECT 13.690 29.235 13.860 29.575 ;
        RECT 14.155 29.375 14.525 29.835 ;
        RECT 12.785 29.065 13.860 29.235 ;
        RECT 14.695 29.205 14.865 29.665 ;
        RECT 15.100 29.325 15.970 29.665 ;
        RECT 16.140 29.375 16.390 29.835 ;
        RECT 14.305 29.035 14.865 29.205 ;
        RECT 14.305 28.895 14.475 29.035 ;
        RECT 12.975 28.725 14.475 28.895 ;
        RECT 15.170 28.865 15.630 29.155 ;
        RECT 12.445 28.385 14.135 28.555 ;
        RECT 12.105 27.965 12.460 28.185 ;
        RECT 12.630 27.675 12.800 28.385 ;
        RECT 13.005 27.965 13.795 28.215 ;
        RECT 13.965 28.205 14.135 28.385 ;
        RECT 14.305 28.035 14.475 28.725 ;
        RECT 10.745 27.285 11.075 27.645 ;
        RECT 11.245 27.505 11.740 27.675 ;
        RECT 11.945 27.505 12.800 27.675 ;
        RECT 13.675 27.285 14.005 27.745 ;
        RECT 14.215 27.645 14.475 28.035 ;
        RECT 14.665 28.855 15.630 28.865 ;
        RECT 15.800 28.945 15.970 29.325 ;
        RECT 16.560 29.285 16.730 29.575 ;
        RECT 16.910 29.455 17.240 29.835 ;
        RECT 16.560 29.115 17.360 29.285 ;
        RECT 14.665 28.695 15.340 28.855 ;
        RECT 15.800 28.775 17.020 28.945 ;
        RECT 14.665 27.905 14.875 28.695 ;
        RECT 15.800 28.685 15.970 28.775 ;
        RECT 15.045 27.905 15.395 28.525 ;
        RECT 15.565 28.515 15.970 28.685 ;
        RECT 15.565 27.735 15.735 28.515 ;
        RECT 15.905 28.065 16.125 28.345 ;
        RECT 16.305 28.235 16.845 28.605 ;
        RECT 17.190 28.525 17.360 29.115 ;
        RECT 17.580 28.695 17.885 29.835 ;
        RECT 18.055 28.645 18.310 29.525 ;
        RECT 18.485 28.670 18.775 29.835 ;
        RECT 18.945 28.760 19.215 29.665 ;
        RECT 19.385 29.075 19.715 29.835 ;
        RECT 19.895 28.905 20.065 29.665 ;
        RECT 17.190 28.495 17.930 28.525 ;
        RECT 15.905 27.895 16.435 28.065 ;
        RECT 14.215 27.475 14.565 27.645 ;
        RECT 14.785 27.455 15.735 27.735 ;
        RECT 15.905 27.285 16.095 27.725 ;
        RECT 16.265 27.665 16.435 27.895 ;
        RECT 16.605 27.835 16.845 28.235 ;
        RECT 17.015 28.195 17.930 28.495 ;
        RECT 17.015 28.020 17.340 28.195 ;
        RECT 17.015 27.665 17.335 28.020 ;
        RECT 18.100 27.995 18.310 28.645 ;
        RECT 16.265 27.495 17.335 27.665 ;
        RECT 17.580 27.285 17.885 27.745 ;
        RECT 18.055 27.465 18.310 27.995 ;
        RECT 18.485 27.285 18.775 28.010 ;
        RECT 18.945 27.960 19.115 28.760 ;
        RECT 19.400 28.735 20.065 28.905 ;
        RECT 20.325 28.745 21.995 29.835 ;
        RECT 19.400 28.590 19.570 28.735 ;
        RECT 19.285 28.260 19.570 28.590 ;
        RECT 19.400 28.005 19.570 28.260 ;
        RECT 19.805 28.185 20.135 28.555 ;
        RECT 20.325 28.055 21.075 28.575 ;
        RECT 21.245 28.225 21.995 28.745 ;
        RECT 22.630 28.695 22.965 29.665 ;
        RECT 23.135 28.695 23.305 29.835 ;
        RECT 23.475 29.495 25.505 29.665 ;
        RECT 18.945 27.455 19.205 27.960 ;
        RECT 19.400 27.835 20.065 28.005 ;
        RECT 19.385 27.285 19.715 27.665 ;
        RECT 19.895 27.455 20.065 27.835 ;
        RECT 20.325 27.285 21.995 28.055 ;
        RECT 22.630 28.025 22.800 28.695 ;
        RECT 23.475 28.525 23.645 29.495 ;
        RECT 22.970 28.195 23.225 28.525 ;
        RECT 23.450 28.195 23.645 28.525 ;
        RECT 23.815 29.155 24.940 29.325 ;
        RECT 23.055 28.025 23.225 28.195 ;
        RECT 23.815 28.025 23.985 29.155 ;
        RECT 22.630 27.455 22.885 28.025 ;
        RECT 23.055 27.855 23.985 28.025 ;
        RECT 24.155 28.815 25.165 28.985 ;
        RECT 24.155 28.015 24.325 28.815 ;
        RECT 24.530 28.475 24.805 28.615 ;
        RECT 24.525 28.305 24.805 28.475 ;
        RECT 23.810 27.820 23.985 27.855 ;
        RECT 23.055 27.285 23.385 27.685 ;
        RECT 23.810 27.455 24.340 27.820 ;
        RECT 24.530 27.455 24.805 28.305 ;
        RECT 24.975 27.455 25.165 28.815 ;
        RECT 25.335 28.830 25.505 29.495 ;
        RECT 25.675 29.075 25.845 29.835 ;
        RECT 26.080 29.075 26.595 29.485 ;
        RECT 25.335 28.640 26.085 28.830 ;
        RECT 26.255 28.265 26.595 29.075 ;
        RECT 26.765 28.745 30.275 29.835 ;
        RECT 25.365 28.095 26.595 28.265 ;
        RECT 25.345 27.285 25.855 27.820 ;
        RECT 26.075 27.490 26.320 28.095 ;
        RECT 26.765 28.055 28.415 28.575 ;
        RECT 28.585 28.225 30.275 28.745 ;
        RECT 30.450 28.695 30.785 29.665 ;
        RECT 30.955 28.695 31.125 29.835 ;
        RECT 31.295 29.495 33.325 29.665 ;
        RECT 26.765 27.285 30.275 28.055 ;
        RECT 30.450 28.025 30.620 28.695 ;
        RECT 31.295 28.525 31.465 29.495 ;
        RECT 30.790 28.195 31.045 28.525 ;
        RECT 31.270 28.195 31.465 28.525 ;
        RECT 31.635 29.155 32.760 29.325 ;
        RECT 30.875 28.025 31.045 28.195 ;
        RECT 31.635 28.025 31.805 29.155 ;
        RECT 30.450 27.455 30.705 28.025 ;
        RECT 30.875 27.855 31.805 28.025 ;
        RECT 31.975 28.815 32.985 28.985 ;
        RECT 31.975 28.015 32.145 28.815 ;
        RECT 32.350 28.475 32.625 28.615 ;
        RECT 32.345 28.305 32.625 28.475 ;
        RECT 31.630 27.820 31.805 27.855 ;
        RECT 30.875 27.285 31.205 27.685 ;
        RECT 31.630 27.455 32.160 27.820 ;
        RECT 32.350 27.455 32.625 28.305 ;
        RECT 32.795 27.455 32.985 28.815 ;
        RECT 33.155 28.830 33.325 29.495 ;
        RECT 33.495 29.075 33.665 29.835 ;
        RECT 33.900 29.075 34.415 29.485 ;
        RECT 33.155 28.640 33.905 28.830 ;
        RECT 34.075 28.265 34.415 29.075 ;
        RECT 34.960 28.855 35.215 29.525 ;
        RECT 35.395 29.035 35.680 29.835 ;
        RECT 35.860 29.115 36.190 29.625 ;
        RECT 34.960 28.815 35.140 28.855 ;
        RECT 34.875 28.645 35.140 28.815 ;
        RECT 33.185 28.095 34.415 28.265 ;
        RECT 33.165 27.285 33.675 27.820 ;
        RECT 33.895 27.490 34.140 28.095 ;
        RECT 34.960 27.995 35.140 28.645 ;
        RECT 35.860 28.525 36.110 29.115 ;
        RECT 36.460 28.965 36.630 29.575 ;
        RECT 36.800 29.145 37.130 29.835 ;
        RECT 37.360 29.285 37.600 29.575 ;
        RECT 37.800 29.455 38.220 29.835 ;
        RECT 38.400 29.365 39.030 29.615 ;
        RECT 39.500 29.455 39.830 29.835 ;
        RECT 38.400 29.285 38.570 29.365 ;
        RECT 40.000 29.285 40.170 29.575 ;
        RECT 40.350 29.455 40.730 29.835 ;
        RECT 40.970 29.450 41.800 29.620 ;
        RECT 37.360 29.115 38.570 29.285 ;
        RECT 35.310 28.195 36.110 28.525 ;
        RECT 34.960 27.465 35.215 27.995 ;
        RECT 35.395 27.285 35.680 27.745 ;
        RECT 35.860 27.545 36.110 28.195 ;
        RECT 36.310 28.945 36.630 28.965 ;
        RECT 36.310 28.775 38.230 28.945 ;
        RECT 36.310 27.880 36.500 28.775 ;
        RECT 38.400 28.605 38.570 29.115 ;
        RECT 38.740 28.855 39.260 29.165 ;
        RECT 36.670 28.435 38.570 28.605 ;
        RECT 36.670 28.375 37.000 28.435 ;
        RECT 37.150 28.205 37.480 28.265 ;
        RECT 36.820 27.935 37.480 28.205 ;
        RECT 36.310 27.550 36.630 27.880 ;
        RECT 36.810 27.285 37.470 27.765 ;
        RECT 37.670 27.675 37.840 28.435 ;
        RECT 38.740 28.265 38.920 28.675 ;
        RECT 38.010 28.095 38.340 28.215 ;
        RECT 39.090 28.095 39.260 28.855 ;
        RECT 38.010 27.925 39.260 28.095 ;
        RECT 39.430 29.035 40.800 29.285 ;
        RECT 39.430 28.265 39.620 29.035 ;
        RECT 40.550 28.775 40.800 29.035 ;
        RECT 39.790 28.605 40.040 28.765 ;
        RECT 40.970 28.605 41.140 29.450 ;
        RECT 42.035 29.165 42.205 29.665 ;
        RECT 42.375 29.335 42.705 29.835 ;
        RECT 41.310 28.775 41.810 29.155 ;
        RECT 42.035 28.995 42.730 29.165 ;
        RECT 39.790 28.435 41.140 28.605 ;
        RECT 40.720 28.395 41.140 28.435 ;
        RECT 39.430 27.925 39.850 28.265 ;
        RECT 40.140 27.935 40.550 28.265 ;
        RECT 37.670 27.505 38.520 27.675 ;
        RECT 39.080 27.285 39.400 27.745 ;
        RECT 39.600 27.495 39.850 27.925 ;
        RECT 40.140 27.285 40.550 27.725 ;
        RECT 40.720 27.665 40.890 28.395 ;
        RECT 41.060 27.845 41.410 28.215 ;
        RECT 41.590 27.905 41.810 28.775 ;
        RECT 41.980 28.205 42.390 28.825 ;
        RECT 42.560 28.025 42.730 28.995 ;
        RECT 42.035 27.835 42.730 28.025 ;
        RECT 40.720 27.465 41.735 27.665 ;
        RECT 42.035 27.505 42.205 27.835 ;
        RECT 42.375 27.285 42.705 27.665 ;
        RECT 42.920 27.545 43.145 29.665 ;
        RECT 43.315 29.335 43.645 29.835 ;
        RECT 43.815 29.165 43.985 29.665 ;
        RECT 43.320 28.995 43.985 29.165 ;
        RECT 43.320 28.005 43.550 28.995 ;
        RECT 43.720 28.175 44.070 28.825 ;
        RECT 44.245 28.670 44.535 29.835 ;
        RECT 44.765 28.695 44.975 29.835 ;
        RECT 45.145 28.685 45.475 29.665 ;
        RECT 45.645 28.695 45.875 29.835 ;
        RECT 46.145 28.695 46.355 29.835 ;
        RECT 46.525 28.685 46.855 29.665 ;
        RECT 47.025 28.695 47.255 29.835 ;
        RECT 47.930 29.165 48.185 29.665 ;
        RECT 48.355 29.335 48.685 29.835 ;
        RECT 47.930 28.995 48.680 29.165 ;
        RECT 43.320 27.835 43.985 28.005 ;
        RECT 43.315 27.285 43.645 27.665 ;
        RECT 43.815 27.545 43.985 27.835 ;
        RECT 44.245 27.285 44.535 28.010 ;
        RECT 44.765 27.285 44.975 28.105 ;
        RECT 45.145 28.085 45.395 28.685 ;
        RECT 45.565 28.275 45.895 28.525 ;
        RECT 45.145 27.455 45.475 28.085 ;
        RECT 45.645 27.285 45.875 28.105 ;
        RECT 46.145 27.285 46.355 28.105 ;
        RECT 46.525 28.085 46.775 28.685 ;
        RECT 46.945 28.275 47.275 28.525 ;
        RECT 47.930 28.175 48.280 28.825 ;
        RECT 46.525 27.455 46.855 28.085 ;
        RECT 47.025 27.285 47.255 28.105 ;
        RECT 48.450 28.005 48.680 28.995 ;
        RECT 47.930 27.835 48.680 28.005 ;
        RECT 47.930 27.545 48.185 27.835 ;
        RECT 48.355 27.285 48.685 27.665 ;
        RECT 48.855 27.545 49.025 29.665 ;
        RECT 49.195 28.865 49.520 29.650 ;
        RECT 49.690 29.375 49.940 29.835 ;
        RECT 50.110 29.335 50.360 29.665 ;
        RECT 50.575 29.335 51.255 29.665 ;
        RECT 50.110 29.205 50.280 29.335 ;
        RECT 49.885 29.035 50.280 29.205 ;
        RECT 49.255 27.815 49.715 28.865 ;
        RECT 49.885 27.675 50.055 29.035 ;
        RECT 50.450 28.775 50.915 29.165 ;
        RECT 50.225 27.965 50.575 28.585 ;
        RECT 50.745 28.185 50.915 28.775 ;
        RECT 51.085 28.555 51.255 29.335 ;
        RECT 51.425 29.235 51.595 29.575 ;
        RECT 51.830 29.405 52.160 29.835 ;
        RECT 52.330 29.235 52.500 29.575 ;
        RECT 52.795 29.375 53.165 29.835 ;
        RECT 51.425 29.065 52.500 29.235 ;
        RECT 53.335 29.205 53.505 29.665 ;
        RECT 53.740 29.325 54.610 29.665 ;
        RECT 54.780 29.375 55.030 29.835 ;
        RECT 52.945 29.035 53.505 29.205 ;
        RECT 52.945 28.895 53.115 29.035 ;
        RECT 51.615 28.725 53.115 28.895 ;
        RECT 53.810 28.865 54.270 29.155 ;
        RECT 51.085 28.385 52.775 28.555 ;
        RECT 50.745 27.965 51.100 28.185 ;
        RECT 51.270 27.675 51.440 28.385 ;
        RECT 51.645 27.965 52.435 28.215 ;
        RECT 52.605 28.205 52.775 28.385 ;
        RECT 52.945 28.035 53.115 28.725 ;
        RECT 49.385 27.285 49.715 27.645 ;
        RECT 49.885 27.505 50.380 27.675 ;
        RECT 50.585 27.505 51.440 27.675 ;
        RECT 52.315 27.285 52.645 27.745 ;
        RECT 52.855 27.645 53.115 28.035 ;
        RECT 53.305 28.855 54.270 28.865 ;
        RECT 54.440 28.945 54.610 29.325 ;
        RECT 55.200 29.285 55.370 29.575 ;
        RECT 55.550 29.455 55.880 29.835 ;
        RECT 55.200 29.115 56.000 29.285 ;
        RECT 53.305 28.695 53.980 28.855 ;
        RECT 54.440 28.775 55.660 28.945 ;
        RECT 53.305 27.905 53.515 28.695 ;
        RECT 54.440 28.685 54.610 28.775 ;
        RECT 53.685 27.905 54.035 28.525 ;
        RECT 54.205 28.515 54.610 28.685 ;
        RECT 54.205 27.735 54.375 28.515 ;
        RECT 54.545 28.065 54.765 28.345 ;
        RECT 54.945 28.235 55.485 28.605 ;
        RECT 55.830 28.525 56.000 29.115 ;
        RECT 56.220 28.695 56.525 29.835 ;
        RECT 56.695 28.645 56.950 29.525 ;
        RECT 55.830 28.495 56.570 28.525 ;
        RECT 54.545 27.895 55.075 28.065 ;
        RECT 52.855 27.475 53.205 27.645 ;
        RECT 53.425 27.455 54.375 27.735 ;
        RECT 54.545 27.285 54.735 27.725 ;
        RECT 54.905 27.665 55.075 27.895 ;
        RECT 55.245 27.835 55.485 28.235 ;
        RECT 55.655 28.195 56.570 28.495 ;
        RECT 55.655 28.020 55.980 28.195 ;
        RECT 55.655 27.665 55.975 28.020 ;
        RECT 56.740 27.995 56.950 28.645 ;
        RECT 54.905 27.495 55.975 27.665 ;
        RECT 56.220 27.285 56.525 27.745 ;
        RECT 56.695 27.465 56.950 27.995 ;
        RECT 57.125 29.335 57.385 29.665 ;
        RECT 57.695 29.455 58.025 29.835 ;
        RECT 57.125 28.655 57.295 29.335 ;
        RECT 58.265 29.285 58.455 29.665 ;
        RECT 58.705 29.455 59.035 29.835 ;
        RECT 59.245 29.285 59.415 29.665 ;
        RECT 59.610 29.455 59.940 29.835 ;
        RECT 60.200 29.285 60.370 29.665 ;
        RECT 60.795 29.455 61.125 29.835 ;
        RECT 57.465 28.825 57.815 29.155 ;
        RECT 58.265 29.115 59.005 29.285 ;
        RECT 58.085 28.775 58.665 28.945 ;
        RECT 58.085 28.655 58.255 28.775 ;
        RECT 57.125 28.485 58.255 28.655 ;
        RECT 58.835 28.605 59.005 29.115 ;
        RECT 57.125 27.785 57.295 28.485 ;
        RECT 58.435 28.435 59.005 28.605 ;
        RECT 59.175 29.115 61.125 29.285 ;
        RECT 57.645 28.145 58.265 28.315 ;
        RECT 57.645 27.965 57.855 28.145 ;
        RECT 58.435 27.955 58.605 28.435 ;
        RECT 59.175 28.125 59.345 29.115 ;
        RECT 59.935 28.525 60.120 28.835 ;
        RECT 60.390 28.525 60.585 28.835 ;
        RECT 57.125 27.455 57.385 27.785 ;
        RECT 57.695 27.285 58.025 27.665 ;
        RECT 58.205 27.625 58.605 27.955 ;
        RECT 58.795 27.795 59.345 28.125 ;
        RECT 59.515 27.625 59.685 28.525 ;
        RECT 58.205 27.455 59.685 27.625 ;
        RECT 59.935 28.195 60.165 28.525 ;
        RECT 60.390 28.195 60.645 28.525 ;
        RECT 60.955 28.195 61.125 29.115 ;
        RECT 59.935 27.615 60.120 28.195 ;
        RECT 60.390 27.620 60.585 28.195 ;
        RECT 60.795 27.285 61.125 27.665 ;
        RECT 61.295 27.455 61.555 29.665 ;
        RECT 61.725 29.400 67.070 29.835 ;
        RECT 63.310 27.830 63.650 28.660 ;
        RECT 65.130 28.150 65.480 29.400 ;
        RECT 67.245 28.745 68.455 29.835 ;
        RECT 67.245 28.035 67.765 28.575 ;
        RECT 67.935 28.205 68.455 28.745 ;
        RECT 68.715 28.905 68.885 29.665 ;
        RECT 69.065 29.075 69.395 29.835 ;
        RECT 68.715 28.735 69.380 28.905 ;
        RECT 69.565 28.760 69.835 29.665 ;
        RECT 69.210 28.590 69.380 28.735 ;
        RECT 68.645 28.185 68.975 28.555 ;
        RECT 69.210 28.260 69.495 28.590 ;
        RECT 61.725 27.285 67.070 27.830 ;
        RECT 67.245 27.285 68.455 28.035 ;
        RECT 69.210 28.005 69.380 28.260 ;
        RECT 68.715 27.835 69.380 28.005 ;
        RECT 69.665 27.960 69.835 28.760 ;
        RECT 70.005 28.670 70.295 29.835 ;
        RECT 70.470 29.165 70.725 29.665 ;
        RECT 70.895 29.335 71.225 29.835 ;
        RECT 70.470 28.995 71.220 29.165 ;
        RECT 70.470 28.175 70.820 28.825 ;
        RECT 68.715 27.455 68.885 27.835 ;
        RECT 69.065 27.285 69.395 27.665 ;
        RECT 69.575 27.455 69.835 27.960 ;
        RECT 70.005 27.285 70.295 28.010 ;
        RECT 70.990 28.005 71.220 28.995 ;
        RECT 70.470 27.835 71.220 28.005 ;
        RECT 70.470 27.545 70.725 27.835 ;
        RECT 70.895 27.285 71.225 27.665 ;
        RECT 71.395 27.545 71.565 29.665 ;
        RECT 71.735 28.865 72.060 29.650 ;
        RECT 72.230 29.375 72.480 29.835 ;
        RECT 72.650 29.335 72.900 29.665 ;
        RECT 73.115 29.335 73.795 29.665 ;
        RECT 72.650 29.205 72.820 29.335 ;
        RECT 72.425 29.035 72.820 29.205 ;
        RECT 71.795 27.815 72.255 28.865 ;
        RECT 72.425 27.675 72.595 29.035 ;
        RECT 72.990 28.775 73.455 29.165 ;
        RECT 72.765 27.965 73.115 28.585 ;
        RECT 73.285 28.185 73.455 28.775 ;
        RECT 73.625 28.555 73.795 29.335 ;
        RECT 73.965 29.235 74.135 29.575 ;
        RECT 74.370 29.405 74.700 29.835 ;
        RECT 74.870 29.235 75.040 29.575 ;
        RECT 75.335 29.375 75.705 29.835 ;
        RECT 73.965 29.065 75.040 29.235 ;
        RECT 75.875 29.205 76.045 29.665 ;
        RECT 76.280 29.325 77.150 29.665 ;
        RECT 77.320 29.375 77.570 29.835 ;
        RECT 75.485 29.035 76.045 29.205 ;
        RECT 75.485 28.895 75.655 29.035 ;
        RECT 74.155 28.725 75.655 28.895 ;
        RECT 76.350 28.865 76.810 29.155 ;
        RECT 73.625 28.385 75.315 28.555 ;
        RECT 73.285 27.965 73.640 28.185 ;
        RECT 73.810 27.675 73.980 28.385 ;
        RECT 74.185 27.965 74.975 28.215 ;
        RECT 75.145 28.205 75.315 28.385 ;
        RECT 75.485 28.035 75.655 28.725 ;
        RECT 71.925 27.285 72.255 27.645 ;
        RECT 72.425 27.505 72.920 27.675 ;
        RECT 73.125 27.505 73.980 27.675 ;
        RECT 74.855 27.285 75.185 27.745 ;
        RECT 75.395 27.645 75.655 28.035 ;
        RECT 75.845 28.855 76.810 28.865 ;
        RECT 76.980 28.945 77.150 29.325 ;
        RECT 77.740 29.285 77.910 29.575 ;
        RECT 78.090 29.455 78.420 29.835 ;
        RECT 77.740 29.115 78.540 29.285 ;
        RECT 75.845 28.695 76.520 28.855 ;
        RECT 76.980 28.775 78.200 28.945 ;
        RECT 75.845 27.905 76.055 28.695 ;
        RECT 76.980 28.685 77.150 28.775 ;
        RECT 76.225 27.905 76.575 28.525 ;
        RECT 76.745 28.515 77.150 28.685 ;
        RECT 76.745 27.735 76.915 28.515 ;
        RECT 77.085 28.065 77.305 28.345 ;
        RECT 77.485 28.235 78.025 28.605 ;
        RECT 78.370 28.525 78.540 29.115 ;
        RECT 78.760 28.695 79.065 29.835 ;
        RECT 79.235 28.645 79.490 29.525 ;
        RECT 78.370 28.495 79.110 28.525 ;
        RECT 77.085 27.895 77.615 28.065 ;
        RECT 75.395 27.475 75.745 27.645 ;
        RECT 75.965 27.455 76.915 27.735 ;
        RECT 77.085 27.285 77.275 27.725 ;
        RECT 77.445 27.665 77.615 27.895 ;
        RECT 77.785 27.835 78.025 28.235 ;
        RECT 78.195 28.195 79.110 28.495 ;
        RECT 78.195 28.020 78.520 28.195 ;
        RECT 78.195 27.665 78.515 28.020 ;
        RECT 79.280 27.995 79.490 28.645 ;
        RECT 77.445 27.495 78.515 27.665 ;
        RECT 78.760 27.285 79.065 27.745 ;
        RECT 79.235 27.465 79.490 27.995 ;
        RECT 79.665 28.760 79.935 29.665 ;
        RECT 80.105 29.075 80.435 29.835 ;
        RECT 80.615 28.905 80.785 29.665 ;
        RECT 79.665 27.960 79.835 28.760 ;
        RECT 80.120 28.735 80.785 28.905 ;
        RECT 80.120 28.590 80.290 28.735 ;
        RECT 81.085 28.695 81.315 29.835 ;
        RECT 81.485 28.685 81.815 29.665 ;
        RECT 81.985 28.695 82.195 29.835 ;
        RECT 82.515 28.905 82.685 29.665 ;
        RECT 82.865 29.075 83.195 29.835 ;
        RECT 82.515 28.735 83.180 28.905 ;
        RECT 83.365 28.760 83.635 29.665 ;
        RECT 80.005 28.260 80.290 28.590 ;
        RECT 80.120 28.005 80.290 28.260 ;
        RECT 80.525 28.185 80.855 28.555 ;
        RECT 81.065 28.275 81.395 28.525 ;
        RECT 79.665 27.455 79.925 27.960 ;
        RECT 80.120 27.835 80.785 28.005 ;
        RECT 80.105 27.285 80.435 27.665 ;
        RECT 80.615 27.455 80.785 27.835 ;
        RECT 81.085 27.285 81.315 28.105 ;
        RECT 81.565 28.085 81.815 28.685 ;
        RECT 83.010 28.590 83.180 28.735 ;
        RECT 82.445 28.185 82.775 28.555 ;
        RECT 83.010 28.260 83.295 28.590 ;
        RECT 81.485 27.455 81.815 28.085 ;
        RECT 81.985 27.285 82.195 28.105 ;
        RECT 83.010 28.005 83.180 28.260 ;
        RECT 82.515 27.835 83.180 28.005 ;
        RECT 83.465 27.960 83.635 28.760 ;
        RECT 83.805 28.745 85.475 29.835 ;
        RECT 86.195 29.165 86.365 29.665 ;
        RECT 86.535 29.335 86.865 29.835 ;
        RECT 86.195 28.995 86.860 29.165 ;
        RECT 82.515 27.455 82.685 27.835 ;
        RECT 82.865 27.285 83.195 27.665 ;
        RECT 83.375 27.455 83.635 27.960 ;
        RECT 83.805 28.055 84.555 28.575 ;
        RECT 84.725 28.225 85.475 28.745 ;
        RECT 86.110 28.175 86.460 28.825 ;
        RECT 83.805 27.285 85.475 28.055 ;
        RECT 86.630 28.005 86.860 28.995 ;
        RECT 86.195 27.835 86.860 28.005 ;
        RECT 86.195 27.545 86.365 27.835 ;
        RECT 86.535 27.285 86.865 27.665 ;
        RECT 87.035 27.545 87.260 29.665 ;
        RECT 87.475 29.335 87.805 29.835 ;
        RECT 87.975 29.165 88.145 29.665 ;
        RECT 88.380 29.450 89.210 29.620 ;
        RECT 89.450 29.455 89.830 29.835 ;
        RECT 87.450 28.995 88.145 29.165 ;
        RECT 87.450 28.025 87.620 28.995 ;
        RECT 87.790 28.205 88.200 28.825 ;
        RECT 88.370 28.775 88.870 29.155 ;
        RECT 87.450 27.835 88.145 28.025 ;
        RECT 88.370 27.905 88.590 28.775 ;
        RECT 89.040 28.605 89.210 29.450 ;
        RECT 90.010 29.285 90.180 29.575 ;
        RECT 90.350 29.455 90.680 29.835 ;
        RECT 91.150 29.365 91.780 29.615 ;
        RECT 91.960 29.455 92.380 29.835 ;
        RECT 91.610 29.285 91.780 29.365 ;
        RECT 92.580 29.285 92.820 29.575 ;
        RECT 89.380 29.035 90.750 29.285 ;
        RECT 89.380 28.775 89.630 29.035 ;
        RECT 90.140 28.605 90.390 28.765 ;
        RECT 89.040 28.435 90.390 28.605 ;
        RECT 89.040 28.395 89.460 28.435 ;
        RECT 88.770 27.845 89.120 28.215 ;
        RECT 87.475 27.285 87.805 27.665 ;
        RECT 87.975 27.505 88.145 27.835 ;
        RECT 89.290 27.665 89.460 28.395 ;
        RECT 90.560 28.265 90.750 29.035 ;
        RECT 89.630 27.935 90.040 28.265 ;
        RECT 90.330 27.925 90.750 28.265 ;
        RECT 90.920 28.855 91.440 29.165 ;
        RECT 91.610 29.115 92.820 29.285 ;
        RECT 93.050 29.145 93.380 29.835 ;
        RECT 90.920 28.095 91.090 28.855 ;
        RECT 91.260 28.265 91.440 28.675 ;
        RECT 91.610 28.605 91.780 29.115 ;
        RECT 93.550 28.965 93.720 29.575 ;
        RECT 93.990 29.115 94.320 29.625 ;
        RECT 93.550 28.945 93.870 28.965 ;
        RECT 91.950 28.775 93.870 28.945 ;
        RECT 91.610 28.435 93.510 28.605 ;
        RECT 91.840 28.095 92.170 28.215 ;
        RECT 90.920 27.925 92.170 28.095 ;
        RECT 88.445 27.465 89.460 27.665 ;
        RECT 89.630 27.285 90.040 27.725 ;
        RECT 90.330 27.495 90.580 27.925 ;
        RECT 90.780 27.285 91.100 27.745 ;
        RECT 92.340 27.675 92.510 28.435 ;
        RECT 93.180 28.375 93.510 28.435 ;
        RECT 92.700 28.205 93.030 28.265 ;
        RECT 92.700 27.935 93.360 28.205 ;
        RECT 93.680 27.880 93.870 28.775 ;
        RECT 91.660 27.505 92.510 27.675 ;
        RECT 92.710 27.285 93.370 27.765 ;
        RECT 93.550 27.550 93.870 27.880 ;
        RECT 94.070 28.525 94.320 29.115 ;
        RECT 94.500 29.035 94.785 29.835 ;
        RECT 94.965 29.495 95.220 29.525 ;
        RECT 94.965 29.325 95.305 29.495 ;
        RECT 94.965 28.855 95.220 29.325 ;
        RECT 94.070 28.195 94.870 28.525 ;
        RECT 94.070 27.545 94.320 28.195 ;
        RECT 95.040 27.995 95.220 28.855 ;
        RECT 95.765 28.670 96.055 29.835 ;
        RECT 96.225 29.400 101.570 29.835 ;
        RECT 101.745 29.400 107.090 29.835 ;
        RECT 94.500 27.285 94.785 27.745 ;
        RECT 94.965 27.465 95.220 27.995 ;
        RECT 95.765 27.285 96.055 28.010 ;
        RECT 97.810 27.830 98.150 28.660 ;
        RECT 99.630 28.150 99.980 29.400 ;
        RECT 103.330 27.830 103.670 28.660 ;
        RECT 105.150 28.150 105.500 29.400 ;
        RECT 107.265 28.745 110.775 29.835 ;
        RECT 110.945 28.745 112.155 29.835 ;
        RECT 107.265 28.055 108.915 28.575 ;
        RECT 109.085 28.225 110.775 28.745 ;
        RECT 96.225 27.285 101.570 27.830 ;
        RECT 101.745 27.285 107.090 27.830 ;
        RECT 107.265 27.285 110.775 28.055 ;
        RECT 110.945 28.035 111.465 28.575 ;
        RECT 111.635 28.205 112.155 28.745 ;
        RECT 112.325 28.745 113.535 29.835 ;
        RECT 112.325 28.205 112.845 28.745 ;
        RECT 113.015 28.035 113.535 28.575 ;
        RECT 110.945 27.285 112.155 28.035 ;
        RECT 112.325 27.285 113.535 28.035 ;
        RECT 5.520 27.115 113.620 27.285 ;
        RECT 5.605 26.365 6.815 27.115 ;
        RECT 6.985 26.570 12.330 27.115 ;
        RECT 5.605 25.825 6.125 26.365 ;
        RECT 6.295 25.655 6.815 26.195 ;
        RECT 8.570 25.740 8.910 26.570 ;
        RECT 12.505 26.345 16.015 27.115 ;
        RECT 5.605 24.565 6.815 25.655 ;
        RECT 10.390 25.000 10.740 26.250 ;
        RECT 12.505 25.825 14.155 26.345 ;
        RECT 16.705 26.295 16.915 27.115 ;
        RECT 17.085 26.315 17.415 26.945 ;
        RECT 14.325 25.655 16.015 26.175 ;
        RECT 17.085 25.715 17.335 26.315 ;
        RECT 17.585 26.295 17.815 27.115 ;
        RECT 18.030 26.565 18.285 26.855 ;
        RECT 18.455 26.735 18.785 27.115 ;
        RECT 18.030 26.395 18.780 26.565 ;
        RECT 17.505 25.875 17.835 26.125 ;
        RECT 6.985 24.565 12.330 25.000 ;
        RECT 12.505 24.565 16.015 25.655 ;
        RECT 16.705 24.565 16.915 25.705 ;
        RECT 17.085 24.735 17.415 25.715 ;
        RECT 17.585 24.565 17.815 25.705 ;
        RECT 18.030 25.575 18.380 26.225 ;
        RECT 18.550 25.405 18.780 26.395 ;
        RECT 18.030 25.235 18.780 25.405 ;
        RECT 18.030 24.735 18.285 25.235 ;
        RECT 18.455 24.565 18.785 25.065 ;
        RECT 18.955 24.735 19.125 26.855 ;
        RECT 19.485 26.755 19.815 27.115 ;
        RECT 19.985 26.725 20.480 26.895 ;
        RECT 20.685 26.725 21.540 26.895 ;
        RECT 19.355 25.535 19.815 26.585 ;
        RECT 19.295 24.750 19.620 25.535 ;
        RECT 19.985 25.365 20.155 26.725 ;
        RECT 20.325 25.815 20.675 26.435 ;
        RECT 20.845 26.215 21.200 26.435 ;
        RECT 20.845 25.625 21.015 26.215 ;
        RECT 21.370 26.015 21.540 26.725 ;
        RECT 22.415 26.655 22.745 27.115 ;
        RECT 22.955 26.755 23.305 26.925 ;
        RECT 21.745 26.185 22.535 26.435 ;
        RECT 22.955 26.365 23.215 26.755 ;
        RECT 23.525 26.665 24.475 26.945 ;
        RECT 24.645 26.675 24.835 27.115 ;
        RECT 25.005 26.735 26.075 26.905 ;
        RECT 22.705 26.015 22.875 26.195 ;
        RECT 19.985 25.195 20.380 25.365 ;
        RECT 20.550 25.235 21.015 25.625 ;
        RECT 21.185 25.845 22.875 26.015 ;
        RECT 20.210 25.065 20.380 25.195 ;
        RECT 21.185 25.065 21.355 25.845 ;
        RECT 23.045 25.675 23.215 26.365 ;
        RECT 21.715 25.505 23.215 25.675 ;
        RECT 23.405 25.705 23.615 26.495 ;
        RECT 23.785 25.875 24.135 26.495 ;
        RECT 24.305 25.885 24.475 26.665 ;
        RECT 25.005 26.505 25.175 26.735 ;
        RECT 24.645 26.335 25.175 26.505 ;
        RECT 24.645 26.055 24.865 26.335 ;
        RECT 25.345 26.165 25.585 26.565 ;
        RECT 24.305 25.715 24.710 25.885 ;
        RECT 25.045 25.795 25.585 26.165 ;
        RECT 25.755 26.380 26.075 26.735 ;
        RECT 26.320 26.655 26.625 27.115 ;
        RECT 26.795 26.405 27.050 26.935 ;
        RECT 25.755 26.205 26.080 26.380 ;
        RECT 25.755 25.905 26.670 26.205 ;
        RECT 25.930 25.875 26.670 25.905 ;
        RECT 23.405 25.545 24.080 25.705 ;
        RECT 24.540 25.625 24.710 25.715 ;
        RECT 23.405 25.535 24.370 25.545 ;
        RECT 23.045 25.365 23.215 25.505 ;
        RECT 19.790 24.565 20.040 25.025 ;
        RECT 20.210 24.735 20.460 25.065 ;
        RECT 20.675 24.735 21.355 25.065 ;
        RECT 21.525 25.165 22.600 25.335 ;
        RECT 23.045 25.195 23.605 25.365 ;
        RECT 23.910 25.245 24.370 25.535 ;
        RECT 24.540 25.455 25.760 25.625 ;
        RECT 21.525 24.825 21.695 25.165 ;
        RECT 21.930 24.565 22.260 24.995 ;
        RECT 22.430 24.825 22.600 25.165 ;
        RECT 22.895 24.565 23.265 25.025 ;
        RECT 23.435 24.735 23.605 25.195 ;
        RECT 24.540 25.075 24.710 25.455 ;
        RECT 25.930 25.285 26.100 25.875 ;
        RECT 26.840 25.755 27.050 26.405 ;
        RECT 27.285 26.295 27.495 27.115 ;
        RECT 27.665 26.315 27.995 26.945 ;
        RECT 23.840 24.735 24.710 25.075 ;
        RECT 25.300 25.115 26.100 25.285 ;
        RECT 24.880 24.565 25.130 25.025 ;
        RECT 25.300 24.825 25.470 25.115 ;
        RECT 25.650 24.565 25.980 24.945 ;
        RECT 26.320 24.565 26.625 25.705 ;
        RECT 26.795 24.875 27.050 25.755 ;
        RECT 27.665 25.715 27.915 26.315 ;
        RECT 28.165 26.295 28.395 27.115 ;
        RECT 28.605 26.365 29.815 27.115 ;
        RECT 30.075 26.565 30.245 26.945 ;
        RECT 30.425 26.735 30.755 27.115 ;
        RECT 30.075 26.395 30.740 26.565 ;
        RECT 30.935 26.440 31.195 26.945 ;
        RECT 28.085 25.875 28.415 26.125 ;
        RECT 28.605 25.825 29.125 26.365 ;
        RECT 27.285 24.565 27.495 25.705 ;
        RECT 27.665 24.735 27.995 25.715 ;
        RECT 28.165 24.565 28.395 25.705 ;
        RECT 29.295 25.655 29.815 26.195 ;
        RECT 30.005 25.845 30.335 26.215 ;
        RECT 30.570 26.140 30.740 26.395 ;
        RECT 30.570 25.810 30.855 26.140 ;
        RECT 30.570 25.665 30.740 25.810 ;
        RECT 28.605 24.565 29.815 25.655 ;
        RECT 30.075 25.495 30.740 25.665 ;
        RECT 31.025 25.640 31.195 26.440 ;
        RECT 31.365 26.390 31.655 27.115 ;
        RECT 31.830 26.405 32.085 26.935 ;
        RECT 32.255 26.655 32.560 27.115 ;
        RECT 32.805 26.735 33.875 26.905 ;
        RECT 31.830 25.755 32.040 26.405 ;
        RECT 32.805 26.380 33.125 26.735 ;
        RECT 32.800 26.205 33.125 26.380 ;
        RECT 32.210 25.905 33.125 26.205 ;
        RECT 33.295 26.165 33.535 26.565 ;
        RECT 33.705 26.505 33.875 26.735 ;
        RECT 34.045 26.675 34.235 27.115 ;
        RECT 34.405 26.665 35.355 26.945 ;
        RECT 35.575 26.755 35.925 26.925 ;
        RECT 33.705 26.335 34.235 26.505 ;
        RECT 32.210 25.875 32.950 25.905 ;
        RECT 30.075 24.735 30.245 25.495 ;
        RECT 30.425 24.565 30.755 25.325 ;
        RECT 30.925 24.735 31.195 25.640 ;
        RECT 31.365 24.565 31.655 25.730 ;
        RECT 31.830 24.875 32.085 25.755 ;
        RECT 32.255 24.565 32.560 25.705 ;
        RECT 32.780 25.285 32.950 25.875 ;
        RECT 33.295 25.795 33.835 26.165 ;
        RECT 34.015 26.055 34.235 26.335 ;
        RECT 34.405 25.885 34.575 26.665 ;
        RECT 34.170 25.715 34.575 25.885 ;
        RECT 34.745 25.875 35.095 26.495 ;
        RECT 34.170 25.625 34.340 25.715 ;
        RECT 35.265 25.705 35.475 26.495 ;
        RECT 33.120 25.455 34.340 25.625 ;
        RECT 34.800 25.545 35.475 25.705 ;
        RECT 32.780 25.115 33.580 25.285 ;
        RECT 32.900 24.565 33.230 24.945 ;
        RECT 33.410 24.825 33.580 25.115 ;
        RECT 34.170 25.075 34.340 25.455 ;
        RECT 34.510 25.535 35.475 25.545 ;
        RECT 35.665 26.365 35.925 26.755 ;
        RECT 36.135 26.655 36.465 27.115 ;
        RECT 37.340 26.725 38.195 26.895 ;
        RECT 38.400 26.725 38.895 26.895 ;
        RECT 39.065 26.755 39.395 27.115 ;
        RECT 35.665 25.675 35.835 26.365 ;
        RECT 36.005 26.015 36.175 26.195 ;
        RECT 36.345 26.185 37.135 26.435 ;
        RECT 37.340 26.015 37.510 26.725 ;
        RECT 37.680 26.215 38.035 26.435 ;
        RECT 36.005 25.845 37.695 26.015 ;
        RECT 34.510 25.245 34.970 25.535 ;
        RECT 35.665 25.505 37.165 25.675 ;
        RECT 35.665 25.365 35.835 25.505 ;
        RECT 35.275 25.195 35.835 25.365 ;
        RECT 33.750 24.565 34.000 25.025 ;
        RECT 34.170 24.735 35.040 25.075 ;
        RECT 35.275 24.735 35.445 25.195 ;
        RECT 36.280 25.165 37.355 25.335 ;
        RECT 35.615 24.565 35.985 25.025 ;
        RECT 36.280 24.825 36.450 25.165 ;
        RECT 36.620 24.565 36.950 24.995 ;
        RECT 37.185 24.825 37.355 25.165 ;
        RECT 37.525 25.065 37.695 25.845 ;
        RECT 37.865 25.625 38.035 26.215 ;
        RECT 38.205 25.815 38.555 26.435 ;
        RECT 37.865 25.235 38.330 25.625 ;
        RECT 38.725 25.365 38.895 26.725 ;
        RECT 39.065 25.535 39.525 26.585 ;
        RECT 38.500 25.195 38.895 25.365 ;
        RECT 38.500 25.065 38.670 25.195 ;
        RECT 37.525 24.735 38.205 25.065 ;
        RECT 38.420 24.735 38.670 25.065 ;
        RECT 38.840 24.565 39.090 25.025 ;
        RECT 39.260 24.750 39.585 25.535 ;
        RECT 39.755 24.735 39.925 26.855 ;
        RECT 40.095 26.735 40.425 27.115 ;
        RECT 40.595 26.565 40.850 26.855 ;
        RECT 40.100 26.395 40.850 26.565 ;
        RECT 41.025 26.440 41.285 26.945 ;
        RECT 41.465 26.735 41.795 27.115 ;
        RECT 41.975 26.565 42.145 26.945 ;
        RECT 42.405 26.570 47.750 27.115 ;
        RECT 47.925 26.570 53.270 27.115 ;
        RECT 40.100 25.405 40.330 26.395 ;
        RECT 40.500 25.575 40.850 26.225 ;
        RECT 41.025 25.640 41.195 26.440 ;
        RECT 41.480 26.395 42.145 26.565 ;
        RECT 41.480 26.140 41.650 26.395 ;
        RECT 41.365 25.810 41.650 26.140 ;
        RECT 41.885 25.845 42.215 26.215 ;
        RECT 41.480 25.665 41.650 25.810 ;
        RECT 43.990 25.740 44.330 26.570 ;
        RECT 40.100 25.235 40.850 25.405 ;
        RECT 40.095 24.565 40.425 25.065 ;
        RECT 40.595 24.735 40.850 25.235 ;
        RECT 41.025 24.735 41.295 25.640 ;
        RECT 41.480 25.495 42.145 25.665 ;
        RECT 41.465 24.565 41.795 25.325 ;
        RECT 41.975 24.735 42.145 25.495 ;
        RECT 45.810 25.000 46.160 26.250 ;
        RECT 49.510 25.740 49.850 26.570 ;
        RECT 53.505 26.295 53.715 27.115 ;
        RECT 53.885 26.315 54.215 26.945 ;
        RECT 51.330 25.000 51.680 26.250 ;
        RECT 53.885 25.715 54.135 26.315 ;
        RECT 54.385 26.295 54.615 27.115 ;
        RECT 54.825 26.345 56.495 27.115 ;
        RECT 57.125 26.390 57.415 27.115 ;
        RECT 57.670 26.545 57.845 26.945 ;
        RECT 58.015 26.735 58.345 27.115 ;
        RECT 58.590 26.615 58.820 26.945 ;
        RECT 57.670 26.375 58.300 26.545 ;
        RECT 54.305 25.875 54.635 26.125 ;
        RECT 54.825 25.825 55.575 26.345 ;
        RECT 58.130 26.205 58.300 26.375 ;
        RECT 42.405 24.565 47.750 25.000 ;
        RECT 47.925 24.565 53.270 25.000 ;
        RECT 53.505 24.565 53.715 25.705 ;
        RECT 53.885 24.735 54.215 25.715 ;
        RECT 54.385 24.565 54.615 25.705 ;
        RECT 55.745 25.655 56.495 26.175 ;
        RECT 54.825 24.565 56.495 25.655 ;
        RECT 57.125 24.565 57.415 25.730 ;
        RECT 57.585 25.525 57.950 26.205 ;
        RECT 58.130 25.875 58.480 26.205 ;
        RECT 58.130 25.355 58.300 25.875 ;
        RECT 57.670 25.185 58.300 25.355 ;
        RECT 58.650 25.325 58.820 26.615 ;
        RECT 59.020 25.505 59.300 26.780 ;
        RECT 59.525 26.775 59.795 26.780 ;
        RECT 59.485 26.605 59.795 26.775 ;
        RECT 60.255 26.735 60.585 27.115 ;
        RECT 60.755 26.860 61.090 26.905 ;
        RECT 59.525 25.505 59.795 26.605 ;
        RECT 59.985 25.505 60.325 26.535 ;
        RECT 60.755 26.395 61.095 26.860 ;
        RECT 60.495 25.875 60.755 26.205 ;
        RECT 60.495 25.325 60.665 25.875 ;
        RECT 60.925 25.705 61.095 26.395 ;
        RECT 57.670 24.735 57.845 25.185 ;
        RECT 58.650 25.155 60.665 25.325 ;
        RECT 58.015 24.565 58.345 25.005 ;
        RECT 58.650 24.735 58.820 25.155 ;
        RECT 59.055 24.565 59.725 24.975 ;
        RECT 59.940 24.735 60.110 25.155 ;
        RECT 60.310 24.565 60.640 24.975 ;
        RECT 60.835 24.735 61.095 25.705 ;
        RECT 61.265 26.615 61.525 26.945 ;
        RECT 61.735 26.635 62.010 27.115 ;
        RECT 61.265 25.705 61.435 26.615 ;
        RECT 62.220 26.545 62.425 26.945 ;
        RECT 62.595 26.715 62.930 27.115 ;
        RECT 63.105 26.570 68.450 27.115 ;
        RECT 61.605 25.875 61.965 26.455 ;
        RECT 62.220 26.375 62.905 26.545 ;
        RECT 62.145 25.705 62.395 26.205 ;
        RECT 61.265 25.535 62.395 25.705 ;
        RECT 61.265 24.765 61.535 25.535 ;
        RECT 62.565 25.345 62.905 26.375 ;
        RECT 64.690 25.740 65.030 26.570 ;
        RECT 68.625 26.345 72.135 27.115 ;
        RECT 61.705 24.565 62.035 25.345 ;
        RECT 62.240 25.170 62.905 25.345 ;
        RECT 62.240 24.765 62.425 25.170 ;
        RECT 66.510 25.000 66.860 26.250 ;
        RECT 68.625 25.825 70.275 26.345 ;
        RECT 72.805 26.295 73.035 27.115 ;
        RECT 73.205 26.315 73.535 26.945 ;
        RECT 70.445 25.655 72.135 26.175 ;
        RECT 72.785 25.875 73.115 26.125 ;
        RECT 73.285 25.715 73.535 26.315 ;
        RECT 73.705 26.295 73.915 27.115 ;
        RECT 74.145 26.570 79.490 27.115 ;
        RECT 75.730 25.740 76.070 26.570 ;
        RECT 79.665 26.345 82.255 27.115 ;
        RECT 82.885 26.390 83.175 27.115 ;
        RECT 83.345 26.570 88.690 27.115 ;
        RECT 88.865 26.570 94.210 27.115 ;
        RECT 94.385 26.570 99.730 27.115 ;
        RECT 99.905 26.570 105.250 27.115 ;
        RECT 62.595 24.565 62.930 24.990 ;
        RECT 63.105 24.565 68.450 25.000 ;
        RECT 68.625 24.565 72.135 25.655 ;
        RECT 72.805 24.565 73.035 25.705 ;
        RECT 73.205 24.735 73.535 25.715 ;
        RECT 73.705 24.565 73.915 25.705 ;
        RECT 77.550 25.000 77.900 26.250 ;
        RECT 79.665 25.825 80.875 26.345 ;
        RECT 81.045 25.655 82.255 26.175 ;
        RECT 84.930 25.740 85.270 26.570 ;
        RECT 74.145 24.565 79.490 25.000 ;
        RECT 79.665 24.565 82.255 25.655 ;
        RECT 82.885 24.565 83.175 25.730 ;
        RECT 86.750 25.000 87.100 26.250 ;
        RECT 90.450 25.740 90.790 26.570 ;
        RECT 92.270 25.000 92.620 26.250 ;
        RECT 95.970 25.740 96.310 26.570 ;
        RECT 97.790 25.000 98.140 26.250 ;
        RECT 101.490 25.740 101.830 26.570 ;
        RECT 105.425 26.345 108.015 27.115 ;
        RECT 108.645 26.390 108.935 27.115 ;
        RECT 109.105 26.345 111.695 27.115 ;
        RECT 112.325 26.365 113.535 27.115 ;
        RECT 103.310 25.000 103.660 26.250 ;
        RECT 105.425 25.825 106.635 26.345 ;
        RECT 106.805 25.655 108.015 26.175 ;
        RECT 109.105 25.825 110.315 26.345 ;
        RECT 83.345 24.565 88.690 25.000 ;
        RECT 88.865 24.565 94.210 25.000 ;
        RECT 94.385 24.565 99.730 25.000 ;
        RECT 99.905 24.565 105.250 25.000 ;
        RECT 105.425 24.565 108.015 25.655 ;
        RECT 108.645 24.565 108.935 25.730 ;
        RECT 110.485 25.655 111.695 26.175 ;
        RECT 109.105 24.565 111.695 25.655 ;
        RECT 112.325 25.655 112.845 26.195 ;
        RECT 113.015 25.825 113.535 26.365 ;
        RECT 112.325 24.565 113.535 25.655 ;
        RECT 5.520 24.395 113.620 24.565 ;
        RECT 5.605 23.305 6.815 24.395 ;
        RECT 6.985 23.960 12.330 24.395 ;
        RECT 12.505 23.960 17.850 24.395 ;
        RECT 5.605 22.595 6.125 23.135 ;
        RECT 6.295 22.765 6.815 23.305 ;
        RECT 5.605 21.845 6.815 22.595 ;
        RECT 8.570 22.390 8.910 23.220 ;
        RECT 10.390 22.710 10.740 23.960 ;
        RECT 14.090 22.390 14.430 23.220 ;
        RECT 15.910 22.710 16.260 23.960 ;
        RECT 18.485 23.230 18.775 24.395 ;
        RECT 18.945 23.305 20.615 24.395 ;
        RECT 18.945 22.615 19.695 23.135 ;
        RECT 19.865 22.785 20.615 23.305 ;
        RECT 20.785 23.320 21.055 24.225 ;
        RECT 21.225 23.635 21.555 24.395 ;
        RECT 21.735 23.465 21.905 24.225 ;
        RECT 22.165 23.960 27.510 24.395 ;
        RECT 6.985 21.845 12.330 22.390 ;
        RECT 12.505 21.845 17.850 22.390 ;
        RECT 18.485 21.845 18.775 22.570 ;
        RECT 18.945 21.845 20.615 22.615 ;
        RECT 20.785 22.520 20.955 23.320 ;
        RECT 21.240 23.295 21.905 23.465 ;
        RECT 21.240 23.150 21.410 23.295 ;
        RECT 21.125 22.820 21.410 23.150 ;
        RECT 21.240 22.565 21.410 22.820 ;
        RECT 21.645 22.745 21.975 23.115 ;
        RECT 20.785 22.015 21.045 22.520 ;
        RECT 21.240 22.395 21.905 22.565 ;
        RECT 21.225 21.845 21.555 22.225 ;
        RECT 21.735 22.015 21.905 22.395 ;
        RECT 23.750 22.390 24.090 23.220 ;
        RECT 25.570 22.710 25.920 23.960 ;
        RECT 27.685 23.305 31.195 24.395 ;
        RECT 31.365 23.305 32.575 24.395 ;
        RECT 27.685 22.615 29.335 23.135 ;
        RECT 29.505 22.785 31.195 23.305 ;
        RECT 22.165 21.845 27.510 22.390 ;
        RECT 27.685 21.845 31.195 22.615 ;
        RECT 31.365 22.595 31.885 23.135 ;
        RECT 32.055 22.765 32.575 23.305 ;
        RECT 32.785 23.255 33.015 24.395 ;
        RECT 33.185 23.245 33.515 24.225 ;
        RECT 33.685 23.255 33.895 24.395 ;
        RECT 34.125 23.960 39.470 24.395 ;
        RECT 32.765 22.835 33.095 23.085 ;
        RECT 31.365 21.845 32.575 22.595 ;
        RECT 32.785 21.845 33.015 22.665 ;
        RECT 33.265 22.645 33.515 23.245 ;
        RECT 33.185 22.015 33.515 22.645 ;
        RECT 33.685 21.845 33.895 22.665 ;
        RECT 35.710 22.390 36.050 23.220 ;
        RECT 37.530 22.710 37.880 23.960 ;
        RECT 39.645 23.305 43.155 24.395 ;
        RECT 39.645 22.615 41.295 23.135 ;
        RECT 41.465 22.785 43.155 23.305 ;
        RECT 44.245 23.230 44.535 24.395 ;
        RECT 44.705 23.960 50.050 24.395 ;
        RECT 34.125 21.845 39.470 22.390 ;
        RECT 39.645 21.845 43.155 22.615 ;
        RECT 44.245 21.845 44.535 22.570 ;
        RECT 46.290 22.390 46.630 23.220 ;
        RECT 48.110 22.710 48.460 23.960 ;
        RECT 50.225 23.305 53.735 24.395 ;
        RECT 50.225 22.615 51.875 23.135 ;
        RECT 52.045 22.785 53.735 23.305 ;
        RECT 53.905 23.425 54.175 24.195 ;
        RECT 54.345 23.615 54.675 24.395 ;
        RECT 54.880 23.790 55.065 24.195 ;
        RECT 55.235 23.970 55.570 24.395 ;
        RECT 54.880 23.615 55.545 23.790 ;
        RECT 53.905 23.255 55.035 23.425 ;
        RECT 44.705 21.845 50.050 22.390 ;
        RECT 50.225 21.845 53.735 22.615 ;
        RECT 53.905 22.345 54.075 23.255 ;
        RECT 54.245 22.505 54.605 23.085 ;
        RECT 54.785 22.755 55.035 23.255 ;
        RECT 55.205 22.585 55.545 23.615 ;
        RECT 55.930 23.425 56.320 23.600 ;
        RECT 56.805 23.595 57.135 24.395 ;
        RECT 57.305 23.605 57.840 24.225 ;
        RECT 55.930 23.255 57.355 23.425 ;
        RECT 54.860 22.415 55.545 22.585 ;
        RECT 55.805 22.525 56.160 23.085 ;
        RECT 53.905 22.015 54.165 22.345 ;
        RECT 54.375 21.845 54.650 22.325 ;
        RECT 54.860 22.015 55.065 22.415 ;
        RECT 56.330 22.355 56.500 23.255 ;
        RECT 56.670 22.525 56.935 23.085 ;
        RECT 57.185 22.755 57.355 23.255 ;
        RECT 57.525 22.585 57.840 23.605 ;
        RECT 58.045 23.255 58.305 24.395 ;
        RECT 58.475 23.425 58.805 24.225 ;
        RECT 58.975 23.595 59.145 24.395 ;
        RECT 59.345 23.425 59.675 24.225 ;
        RECT 59.875 23.595 60.155 24.395 ;
        RECT 58.475 23.255 59.755 23.425 ;
        RECT 58.070 22.755 58.355 23.085 ;
        RECT 58.555 22.755 58.935 23.085 ;
        RECT 59.105 22.755 59.415 23.085 ;
        RECT 55.235 21.845 55.570 22.245 ;
        RECT 55.910 21.845 56.150 22.355 ;
        RECT 56.330 22.025 56.610 22.355 ;
        RECT 56.840 21.845 57.055 22.355 ;
        RECT 57.225 22.015 57.840 22.585 ;
        RECT 58.050 21.845 58.385 22.585 ;
        RECT 58.555 22.060 58.770 22.755 ;
        RECT 59.105 22.585 59.310 22.755 ;
        RECT 59.585 22.585 59.755 23.255 ;
        RECT 59.935 22.755 60.175 23.425 ;
        RECT 60.345 23.255 60.620 24.225 ;
        RECT 60.830 23.595 61.110 24.395 ;
        RECT 61.280 23.885 62.895 24.215 ;
        RECT 61.280 23.545 62.455 23.715 ;
        RECT 61.280 23.425 61.450 23.545 ;
        RECT 60.790 23.255 61.450 23.425 ;
        RECT 58.960 22.060 59.310 22.585 ;
        RECT 59.480 22.015 60.175 22.585 ;
        RECT 60.345 22.520 60.515 23.255 ;
        RECT 60.790 23.085 60.960 23.255 ;
        RECT 61.710 23.085 61.955 23.375 ;
        RECT 62.125 23.255 62.455 23.545 ;
        RECT 62.715 23.085 62.885 23.645 ;
        RECT 63.135 23.255 63.395 24.395 ;
        RECT 63.575 23.335 63.905 24.185 ;
        RECT 60.685 22.755 60.960 23.085 ;
        RECT 61.130 22.755 61.955 23.085 ;
        RECT 62.170 22.755 62.885 23.085 ;
        RECT 63.055 22.835 63.390 23.085 ;
        RECT 60.790 22.585 60.960 22.755 ;
        RECT 62.635 22.665 62.885 22.755 ;
        RECT 60.345 22.175 60.620 22.520 ;
        RECT 60.790 22.415 62.455 22.585 ;
        RECT 60.810 21.845 61.185 22.245 ;
        RECT 61.355 22.065 61.525 22.415 ;
        RECT 61.695 21.845 62.025 22.245 ;
        RECT 62.195 22.015 62.455 22.415 ;
        RECT 62.635 22.245 62.965 22.665 ;
        RECT 63.135 21.845 63.395 22.665 ;
        RECT 63.575 22.570 63.765 23.335 ;
        RECT 64.075 23.255 64.325 24.395 ;
        RECT 64.515 23.755 64.765 24.175 ;
        RECT 64.995 23.925 65.325 24.395 ;
        RECT 65.555 23.755 65.805 24.175 ;
        RECT 64.515 23.585 65.805 23.755 ;
        RECT 65.985 23.755 66.315 24.185 ;
        RECT 65.985 23.585 66.440 23.755 ;
        RECT 64.505 23.085 64.720 23.415 ;
        RECT 63.935 22.755 64.245 23.085 ;
        RECT 64.415 22.755 64.720 23.085 ;
        RECT 64.895 22.755 65.180 23.415 ;
        RECT 65.375 22.755 65.640 23.415 ;
        RECT 65.855 22.755 66.100 23.415 ;
        RECT 64.075 22.585 64.245 22.755 ;
        RECT 66.270 22.585 66.440 23.585 ;
        RECT 66.785 23.305 69.375 24.395 ;
        RECT 63.575 22.060 63.905 22.570 ;
        RECT 64.075 22.415 66.440 22.585 ;
        RECT 66.785 22.615 67.995 23.135 ;
        RECT 68.165 22.785 69.375 23.305 ;
        RECT 70.005 23.230 70.295 24.395 ;
        RECT 70.465 23.960 75.810 24.395 ;
        RECT 64.075 21.845 64.405 22.245 ;
        RECT 65.455 22.075 65.785 22.415 ;
        RECT 65.955 21.845 66.285 22.245 ;
        RECT 66.785 21.845 69.375 22.615 ;
        RECT 70.005 21.845 70.295 22.570 ;
        RECT 72.050 22.390 72.390 23.220 ;
        RECT 73.870 22.710 74.220 23.960 ;
        RECT 75.985 23.305 77.655 24.395 ;
        RECT 75.985 22.615 76.735 23.135 ;
        RECT 76.905 22.785 77.655 23.305 ;
        RECT 78.290 23.205 78.545 24.085 ;
        RECT 78.715 23.255 79.020 24.395 ;
        RECT 79.360 24.015 79.690 24.395 ;
        RECT 79.870 23.845 80.040 24.135 ;
        RECT 80.210 23.935 80.460 24.395 ;
        RECT 79.240 23.675 80.040 23.845 ;
        RECT 80.630 23.885 81.500 24.225 ;
        RECT 70.465 21.845 75.810 22.390 ;
        RECT 75.985 21.845 77.655 22.615 ;
        RECT 78.290 22.555 78.500 23.205 ;
        RECT 79.240 23.085 79.410 23.675 ;
        RECT 80.630 23.505 80.800 23.885 ;
        RECT 81.735 23.765 81.905 24.225 ;
        RECT 82.075 23.935 82.445 24.395 ;
        RECT 82.740 23.795 82.910 24.135 ;
        RECT 83.080 23.965 83.410 24.395 ;
        RECT 83.645 23.795 83.815 24.135 ;
        RECT 79.580 23.335 80.800 23.505 ;
        RECT 80.970 23.425 81.430 23.715 ;
        RECT 81.735 23.595 82.295 23.765 ;
        RECT 82.740 23.625 83.815 23.795 ;
        RECT 83.985 23.895 84.665 24.225 ;
        RECT 84.880 23.895 85.130 24.225 ;
        RECT 85.300 23.935 85.550 24.395 ;
        RECT 82.125 23.455 82.295 23.595 ;
        RECT 80.970 23.415 81.935 23.425 ;
        RECT 80.630 23.245 80.800 23.335 ;
        RECT 81.260 23.255 81.935 23.415 ;
        RECT 78.670 23.055 79.410 23.085 ;
        RECT 78.670 22.755 79.585 23.055 ;
        RECT 79.260 22.580 79.585 22.755 ;
        RECT 78.290 22.025 78.545 22.555 ;
        RECT 78.715 21.845 79.020 22.305 ;
        RECT 79.265 22.225 79.585 22.580 ;
        RECT 79.755 22.795 80.295 23.165 ;
        RECT 80.630 23.075 81.035 23.245 ;
        RECT 79.755 22.395 79.995 22.795 ;
        RECT 80.475 22.625 80.695 22.905 ;
        RECT 80.165 22.455 80.695 22.625 ;
        RECT 80.165 22.225 80.335 22.455 ;
        RECT 80.865 22.295 81.035 23.075 ;
        RECT 81.205 22.465 81.555 23.085 ;
        RECT 81.725 22.465 81.935 23.255 ;
        RECT 82.125 23.285 83.625 23.455 ;
        RECT 82.125 22.595 82.295 23.285 ;
        RECT 83.985 23.115 84.155 23.895 ;
        RECT 84.960 23.765 85.130 23.895 ;
        RECT 82.465 22.945 84.155 23.115 ;
        RECT 84.325 23.335 84.790 23.725 ;
        RECT 84.960 23.595 85.355 23.765 ;
        RECT 82.465 22.765 82.635 22.945 ;
        RECT 79.265 22.055 80.335 22.225 ;
        RECT 80.505 21.845 80.695 22.285 ;
        RECT 80.865 22.015 81.815 22.295 ;
        RECT 82.125 22.205 82.385 22.595 ;
        RECT 82.805 22.525 83.595 22.775 ;
        RECT 82.035 22.035 82.385 22.205 ;
        RECT 82.595 21.845 82.925 22.305 ;
        RECT 83.800 22.235 83.970 22.945 ;
        RECT 84.325 22.745 84.495 23.335 ;
        RECT 84.140 22.525 84.495 22.745 ;
        RECT 84.665 22.525 85.015 23.145 ;
        RECT 85.185 22.235 85.355 23.595 ;
        RECT 85.720 23.425 86.045 24.210 ;
        RECT 85.525 22.375 85.985 23.425 ;
        RECT 83.800 22.065 84.655 22.235 ;
        RECT 84.860 22.065 85.355 22.235 ;
        RECT 85.525 21.845 85.855 22.205 ;
        RECT 86.215 22.105 86.385 24.225 ;
        RECT 86.555 23.895 86.885 24.395 ;
        RECT 87.055 23.725 87.310 24.225 ;
        RECT 87.485 23.960 92.830 24.395 ;
        RECT 86.560 23.555 87.310 23.725 ;
        RECT 86.560 22.565 86.790 23.555 ;
        RECT 86.960 22.735 87.310 23.385 ;
        RECT 86.560 22.395 87.310 22.565 ;
        RECT 86.555 21.845 86.885 22.225 ;
        RECT 87.055 22.105 87.310 22.395 ;
        RECT 89.070 22.390 89.410 23.220 ;
        RECT 90.890 22.710 91.240 23.960 ;
        RECT 93.005 23.305 95.595 24.395 ;
        RECT 93.005 22.615 94.215 23.135 ;
        RECT 94.385 22.785 95.595 23.305 ;
        RECT 95.765 23.230 96.055 24.395 ;
        RECT 96.225 23.960 101.570 24.395 ;
        RECT 101.745 23.960 107.090 24.395 ;
        RECT 87.485 21.845 92.830 22.390 ;
        RECT 93.005 21.845 95.595 22.615 ;
        RECT 95.765 21.845 96.055 22.570 ;
        RECT 97.810 22.390 98.150 23.220 ;
        RECT 99.630 22.710 99.980 23.960 ;
        RECT 103.330 22.390 103.670 23.220 ;
        RECT 105.150 22.710 105.500 23.960 ;
        RECT 107.265 23.305 110.775 24.395 ;
        RECT 110.945 23.305 112.155 24.395 ;
        RECT 107.265 22.615 108.915 23.135 ;
        RECT 109.085 22.785 110.775 23.305 ;
        RECT 96.225 21.845 101.570 22.390 ;
        RECT 101.745 21.845 107.090 22.390 ;
        RECT 107.265 21.845 110.775 22.615 ;
        RECT 110.945 22.595 111.465 23.135 ;
        RECT 111.635 22.765 112.155 23.305 ;
        RECT 112.325 23.305 113.535 24.395 ;
        RECT 112.325 22.765 112.845 23.305 ;
        RECT 113.015 22.595 113.535 23.135 ;
        RECT 110.945 21.845 112.155 22.595 ;
        RECT 112.325 21.845 113.535 22.595 ;
        RECT 5.520 21.675 113.620 21.845 ;
        RECT 5.605 20.925 6.815 21.675 ;
        RECT 6.985 21.130 12.330 21.675 ;
        RECT 12.505 21.130 17.850 21.675 ;
        RECT 18.025 21.130 23.370 21.675 ;
        RECT 23.545 21.130 28.890 21.675 ;
        RECT 5.605 20.385 6.125 20.925 ;
        RECT 6.295 20.215 6.815 20.755 ;
        RECT 8.570 20.300 8.910 21.130 ;
        RECT 5.605 19.125 6.815 20.215 ;
        RECT 10.390 19.560 10.740 20.810 ;
        RECT 14.090 20.300 14.430 21.130 ;
        RECT 15.910 19.560 16.260 20.810 ;
        RECT 19.610 20.300 19.950 21.130 ;
        RECT 21.430 19.560 21.780 20.810 ;
        RECT 25.130 20.300 25.470 21.130 ;
        RECT 29.065 20.905 30.735 21.675 ;
        RECT 31.365 20.950 31.655 21.675 ;
        RECT 31.825 21.130 37.170 21.675 ;
        RECT 37.345 21.130 42.690 21.675 ;
        RECT 42.865 21.130 48.210 21.675 ;
        RECT 26.950 19.560 27.300 20.810 ;
        RECT 29.065 20.385 29.815 20.905 ;
        RECT 29.985 20.215 30.735 20.735 ;
        RECT 33.410 20.300 33.750 21.130 ;
        RECT 6.985 19.125 12.330 19.560 ;
        RECT 12.505 19.125 17.850 19.560 ;
        RECT 18.025 19.125 23.370 19.560 ;
        RECT 23.545 19.125 28.890 19.560 ;
        RECT 29.065 19.125 30.735 20.215 ;
        RECT 31.365 19.125 31.655 20.290 ;
        RECT 35.230 19.560 35.580 20.810 ;
        RECT 38.930 20.300 39.270 21.130 ;
        RECT 40.750 19.560 41.100 20.810 ;
        RECT 44.450 20.300 44.790 21.130 ;
        RECT 48.385 20.925 49.595 21.675 ;
        RECT 49.765 21.000 50.025 21.505 ;
        RECT 50.205 21.295 50.535 21.675 ;
        RECT 50.715 21.125 50.885 21.505 ;
        RECT 46.270 19.560 46.620 20.810 ;
        RECT 48.385 20.385 48.905 20.925 ;
        RECT 49.075 20.215 49.595 20.755 ;
        RECT 31.825 19.125 37.170 19.560 ;
        RECT 37.345 19.125 42.690 19.560 ;
        RECT 42.865 19.125 48.210 19.560 ;
        RECT 48.385 19.125 49.595 20.215 ;
        RECT 49.765 20.200 49.935 21.000 ;
        RECT 50.220 20.955 50.885 21.125 ;
        RECT 50.220 20.700 50.390 20.955 ;
        RECT 51.150 20.835 51.410 21.675 ;
        RECT 51.585 20.930 51.840 21.505 ;
        RECT 52.010 21.295 52.340 21.675 ;
        RECT 52.555 21.125 52.725 21.505 ;
        RECT 52.010 20.955 52.725 21.125 ;
        RECT 50.105 20.370 50.390 20.700 ;
        RECT 50.625 20.405 50.955 20.775 ;
        RECT 50.220 20.225 50.390 20.370 ;
        RECT 49.765 19.295 50.035 20.200 ;
        RECT 50.220 20.055 50.885 20.225 ;
        RECT 50.205 19.125 50.535 19.885 ;
        RECT 50.715 19.295 50.885 20.055 ;
        RECT 51.150 19.125 51.410 20.275 ;
        RECT 51.585 20.200 51.755 20.930 ;
        RECT 52.010 20.765 52.180 20.955 ;
        RECT 52.985 20.935 53.305 21.415 ;
        RECT 53.475 21.105 53.705 21.505 ;
        RECT 53.875 21.285 54.225 21.675 ;
        RECT 53.475 21.025 53.985 21.105 ;
        RECT 54.395 21.025 54.725 21.505 ;
        RECT 53.475 20.935 54.725 21.025 ;
        RECT 51.925 20.435 52.180 20.765 ;
        RECT 52.010 20.225 52.180 20.435 ;
        RECT 52.460 20.405 52.815 20.775 ;
        RECT 51.585 19.295 51.840 20.200 ;
        RECT 52.010 20.055 52.725 20.225 ;
        RECT 52.010 19.125 52.340 19.885 ;
        RECT 52.555 19.295 52.725 20.055 ;
        RECT 52.985 20.005 53.155 20.935 ;
        RECT 53.815 20.855 54.725 20.935 ;
        RECT 54.895 20.855 55.065 21.675 ;
        RECT 55.570 20.935 56.035 21.480 ;
        RECT 57.125 20.950 57.415 21.675 ;
        RECT 53.325 20.345 53.495 20.765 ;
        RECT 53.725 20.515 54.325 20.685 ;
        RECT 53.325 20.175 53.985 20.345 ;
        RECT 52.985 19.805 53.645 20.005 ;
        RECT 53.815 19.975 53.985 20.175 ;
        RECT 54.155 20.315 54.325 20.515 ;
        RECT 54.495 20.485 55.190 20.685 ;
        RECT 55.450 20.315 55.695 20.765 ;
        RECT 54.155 20.145 55.695 20.315 ;
        RECT 55.865 19.975 56.035 20.935 ;
        RECT 57.585 20.875 58.280 21.505 ;
        RECT 58.485 20.875 58.795 21.675 ;
        RECT 58.965 21.000 59.240 21.345 ;
        RECT 59.430 21.275 59.805 21.675 ;
        RECT 59.975 21.105 60.145 21.455 ;
        RECT 60.315 21.275 60.645 21.675 ;
        RECT 60.815 21.105 61.075 21.505 ;
        RECT 57.605 20.435 57.940 20.685 ;
        RECT 58.110 20.315 58.280 20.875 ;
        RECT 58.450 20.435 58.785 20.705 ;
        RECT 53.815 19.805 56.035 19.975 ;
        RECT 53.475 19.635 53.645 19.805 ;
        RECT 53.005 19.125 53.305 19.635 ;
        RECT 53.475 19.465 53.855 19.635 ;
        RECT 54.435 19.125 55.065 19.635 ;
        RECT 55.235 19.295 55.565 19.805 ;
        RECT 55.735 19.125 56.035 19.635 ;
        RECT 57.125 19.125 57.415 20.290 ;
        RECT 58.105 20.275 58.280 20.315 ;
        RECT 57.585 19.125 57.845 20.265 ;
        RECT 58.015 19.295 58.345 20.275 ;
        RECT 58.965 20.265 59.135 21.000 ;
        RECT 59.410 20.935 61.075 21.105 ;
        RECT 59.410 20.765 59.580 20.935 ;
        RECT 61.255 20.855 61.585 21.275 ;
        RECT 61.755 20.855 62.015 21.675 ;
        RECT 62.185 20.935 62.650 21.480 ;
        RECT 61.255 20.765 61.505 20.855 ;
        RECT 59.305 20.435 59.580 20.765 ;
        RECT 59.750 20.435 60.575 20.765 ;
        RECT 60.790 20.435 61.505 20.765 ;
        RECT 61.675 20.435 62.010 20.685 ;
        RECT 59.410 20.265 59.580 20.435 ;
        RECT 58.515 19.125 58.795 20.265 ;
        RECT 58.965 19.295 59.240 20.265 ;
        RECT 59.410 20.095 60.070 20.265 ;
        RECT 60.330 20.145 60.575 20.435 ;
        RECT 59.900 19.975 60.070 20.095 ;
        RECT 60.745 19.975 61.075 20.265 ;
        RECT 59.450 19.125 59.730 19.925 ;
        RECT 59.900 19.805 61.075 19.975 ;
        RECT 61.335 19.875 61.505 20.435 ;
        RECT 59.900 19.305 61.515 19.635 ;
        RECT 61.755 19.125 62.015 20.265 ;
        RECT 62.185 19.975 62.355 20.935 ;
        RECT 63.155 20.855 63.325 21.675 ;
        RECT 63.495 21.025 63.825 21.505 ;
        RECT 63.995 21.285 64.345 21.675 ;
        RECT 64.515 21.105 64.745 21.505 ;
        RECT 64.235 21.025 64.745 21.105 ;
        RECT 63.495 20.935 64.745 21.025 ;
        RECT 64.915 20.935 65.235 21.415 ;
        RECT 65.410 21.125 65.665 21.415 ;
        RECT 65.835 21.295 66.165 21.675 ;
        RECT 65.410 20.955 66.160 21.125 ;
        RECT 63.495 20.855 64.405 20.935 ;
        RECT 62.525 20.315 62.770 20.765 ;
        RECT 63.030 20.485 63.725 20.685 ;
        RECT 63.895 20.515 64.495 20.685 ;
        RECT 63.895 20.315 64.065 20.515 ;
        RECT 64.725 20.345 64.895 20.765 ;
        RECT 62.525 20.145 64.065 20.315 ;
        RECT 64.235 20.175 64.895 20.345 ;
        RECT 64.235 19.975 64.405 20.175 ;
        RECT 65.065 20.005 65.235 20.935 ;
        RECT 65.410 20.135 65.760 20.785 ;
        RECT 62.185 19.805 64.405 19.975 ;
        RECT 64.575 19.805 65.235 20.005 ;
        RECT 65.930 19.965 66.160 20.955 ;
        RECT 62.185 19.125 62.485 19.635 ;
        RECT 62.655 19.295 62.985 19.805 ;
        RECT 64.575 19.635 64.745 19.805 ;
        RECT 65.410 19.795 66.160 19.965 ;
        RECT 63.155 19.125 63.785 19.635 ;
        RECT 64.365 19.465 64.745 19.635 ;
        RECT 64.915 19.125 65.215 19.635 ;
        RECT 65.410 19.295 65.665 19.795 ;
        RECT 65.835 19.125 66.165 19.625 ;
        RECT 66.335 19.295 66.505 21.415 ;
        RECT 66.865 21.315 67.195 21.675 ;
        RECT 67.365 21.285 67.860 21.455 ;
        RECT 68.065 21.285 68.920 21.455 ;
        RECT 66.735 20.095 67.195 21.145 ;
        RECT 66.675 19.310 67.000 20.095 ;
        RECT 67.365 19.925 67.535 21.285 ;
        RECT 67.705 20.375 68.055 20.995 ;
        RECT 68.225 20.775 68.580 20.995 ;
        RECT 68.225 20.185 68.395 20.775 ;
        RECT 68.750 20.575 68.920 21.285 ;
        RECT 69.795 21.215 70.125 21.675 ;
        RECT 70.335 21.315 70.685 21.485 ;
        RECT 69.125 20.745 69.915 20.995 ;
        RECT 70.335 20.925 70.595 21.315 ;
        RECT 70.905 21.225 71.855 21.505 ;
        RECT 72.025 21.235 72.215 21.675 ;
        RECT 72.385 21.295 73.455 21.465 ;
        RECT 70.085 20.575 70.255 20.755 ;
        RECT 67.365 19.755 67.760 19.925 ;
        RECT 67.930 19.795 68.395 20.185 ;
        RECT 68.565 20.405 70.255 20.575 ;
        RECT 67.590 19.625 67.760 19.755 ;
        RECT 68.565 19.625 68.735 20.405 ;
        RECT 70.425 20.235 70.595 20.925 ;
        RECT 69.095 20.065 70.595 20.235 ;
        RECT 70.785 20.265 70.995 21.055 ;
        RECT 71.165 20.435 71.515 21.055 ;
        RECT 71.685 20.445 71.855 21.225 ;
        RECT 72.385 21.065 72.555 21.295 ;
        RECT 72.025 20.895 72.555 21.065 ;
        RECT 72.025 20.615 72.245 20.895 ;
        RECT 72.725 20.725 72.965 21.125 ;
        RECT 71.685 20.275 72.090 20.445 ;
        RECT 72.425 20.355 72.965 20.725 ;
        RECT 73.135 20.940 73.455 21.295 ;
        RECT 73.700 21.215 74.005 21.675 ;
        RECT 74.175 20.965 74.425 21.495 ;
        RECT 73.135 20.765 73.460 20.940 ;
        RECT 73.135 20.465 74.050 20.765 ;
        RECT 73.310 20.435 74.050 20.465 ;
        RECT 70.785 20.105 71.460 20.265 ;
        RECT 71.920 20.185 72.090 20.275 ;
        RECT 70.785 20.095 71.750 20.105 ;
        RECT 70.425 19.925 70.595 20.065 ;
        RECT 67.170 19.125 67.420 19.585 ;
        RECT 67.590 19.295 67.840 19.625 ;
        RECT 68.055 19.295 68.735 19.625 ;
        RECT 68.905 19.725 69.980 19.895 ;
        RECT 70.425 19.755 70.985 19.925 ;
        RECT 71.290 19.805 71.750 20.095 ;
        RECT 71.920 20.015 73.140 20.185 ;
        RECT 68.905 19.385 69.075 19.725 ;
        RECT 69.310 19.125 69.640 19.555 ;
        RECT 69.810 19.385 69.980 19.725 ;
        RECT 70.275 19.125 70.645 19.585 ;
        RECT 70.815 19.295 70.985 19.755 ;
        RECT 71.920 19.635 72.090 20.015 ;
        RECT 73.310 19.845 73.480 20.435 ;
        RECT 74.220 20.315 74.425 20.965 ;
        RECT 74.595 20.920 74.845 21.675 ;
        RECT 75.065 21.130 80.410 21.675 ;
        RECT 71.220 19.295 72.090 19.635 ;
        RECT 72.680 19.675 73.480 19.845 ;
        RECT 72.260 19.125 72.510 19.585 ;
        RECT 72.680 19.385 72.850 19.675 ;
        RECT 73.030 19.125 73.360 19.505 ;
        RECT 73.700 19.125 74.005 20.265 ;
        RECT 74.175 19.435 74.425 20.315 ;
        RECT 76.650 20.300 76.990 21.130 ;
        RECT 80.585 20.905 82.255 21.675 ;
        RECT 82.885 20.950 83.175 21.675 ;
        RECT 83.345 21.130 88.690 21.675 ;
        RECT 88.865 21.130 94.210 21.675 ;
        RECT 94.385 21.130 99.730 21.675 ;
        RECT 99.905 21.130 105.250 21.675 ;
        RECT 74.595 19.125 74.845 20.265 ;
        RECT 78.470 19.560 78.820 20.810 ;
        RECT 80.585 20.385 81.335 20.905 ;
        RECT 81.505 20.215 82.255 20.735 ;
        RECT 84.930 20.300 85.270 21.130 ;
        RECT 75.065 19.125 80.410 19.560 ;
        RECT 80.585 19.125 82.255 20.215 ;
        RECT 82.885 19.125 83.175 20.290 ;
        RECT 86.750 19.560 87.100 20.810 ;
        RECT 90.450 20.300 90.790 21.130 ;
        RECT 92.270 19.560 92.620 20.810 ;
        RECT 95.970 20.300 96.310 21.130 ;
        RECT 97.790 19.560 98.140 20.810 ;
        RECT 101.490 20.300 101.830 21.130 ;
        RECT 105.425 20.905 108.015 21.675 ;
        RECT 108.645 20.950 108.935 21.675 ;
        RECT 109.105 20.905 111.695 21.675 ;
        RECT 112.325 20.925 113.535 21.675 ;
        RECT 103.310 19.560 103.660 20.810 ;
        RECT 105.425 20.385 106.635 20.905 ;
        RECT 106.805 20.215 108.015 20.735 ;
        RECT 109.105 20.385 110.315 20.905 ;
        RECT 83.345 19.125 88.690 19.560 ;
        RECT 88.865 19.125 94.210 19.560 ;
        RECT 94.385 19.125 99.730 19.560 ;
        RECT 99.905 19.125 105.250 19.560 ;
        RECT 105.425 19.125 108.015 20.215 ;
        RECT 108.645 19.125 108.935 20.290 ;
        RECT 110.485 20.215 111.695 20.735 ;
        RECT 109.105 19.125 111.695 20.215 ;
        RECT 112.325 20.215 112.845 20.755 ;
        RECT 113.015 20.385 113.535 20.925 ;
        RECT 112.325 19.125 113.535 20.215 ;
        RECT 5.520 18.955 113.620 19.125 ;
        RECT 5.605 17.865 6.815 18.955 ;
        RECT 6.985 18.520 12.330 18.955 ;
        RECT 12.505 18.520 17.850 18.955 ;
        RECT 5.605 17.155 6.125 17.695 ;
        RECT 6.295 17.325 6.815 17.865 ;
        RECT 5.605 16.405 6.815 17.155 ;
        RECT 8.570 16.950 8.910 17.780 ;
        RECT 10.390 17.270 10.740 18.520 ;
        RECT 14.090 16.950 14.430 17.780 ;
        RECT 15.910 17.270 16.260 18.520 ;
        RECT 18.485 17.790 18.775 18.955 ;
        RECT 18.945 18.520 24.290 18.955 ;
        RECT 24.465 18.520 29.810 18.955 ;
        RECT 29.985 18.520 35.330 18.955 ;
        RECT 35.505 18.520 40.850 18.955 ;
        RECT 6.985 16.405 12.330 16.950 ;
        RECT 12.505 16.405 17.850 16.950 ;
        RECT 18.485 16.405 18.775 17.130 ;
        RECT 20.530 16.950 20.870 17.780 ;
        RECT 22.350 17.270 22.700 18.520 ;
        RECT 26.050 16.950 26.390 17.780 ;
        RECT 27.870 17.270 28.220 18.520 ;
        RECT 31.570 16.950 31.910 17.780 ;
        RECT 33.390 17.270 33.740 18.520 ;
        RECT 37.090 16.950 37.430 17.780 ;
        RECT 38.910 17.270 39.260 18.520 ;
        RECT 41.025 17.865 43.615 18.955 ;
        RECT 41.025 17.175 42.235 17.695 ;
        RECT 42.405 17.345 43.615 17.865 ;
        RECT 44.245 17.790 44.535 18.955 ;
        RECT 44.705 17.865 46.375 18.955 ;
        RECT 44.705 17.175 45.455 17.695 ;
        RECT 45.625 17.345 46.375 17.865 ;
        RECT 46.585 17.815 46.815 18.955 ;
        RECT 46.985 17.805 47.315 18.785 ;
        RECT 47.485 17.815 47.695 18.955 ;
        RECT 47.930 18.285 48.185 18.785 ;
        RECT 48.355 18.455 48.685 18.955 ;
        RECT 47.930 18.115 48.680 18.285 ;
        RECT 46.565 17.395 46.895 17.645 ;
        RECT 18.945 16.405 24.290 16.950 ;
        RECT 24.465 16.405 29.810 16.950 ;
        RECT 29.985 16.405 35.330 16.950 ;
        RECT 35.505 16.405 40.850 16.950 ;
        RECT 41.025 16.405 43.615 17.175 ;
        RECT 44.245 16.405 44.535 17.130 ;
        RECT 44.705 16.405 46.375 17.175 ;
        RECT 46.585 16.405 46.815 17.225 ;
        RECT 47.065 17.205 47.315 17.805 ;
        RECT 47.930 17.295 48.280 17.945 ;
        RECT 46.985 16.575 47.315 17.205 ;
        RECT 47.485 16.405 47.695 17.225 ;
        RECT 48.450 17.125 48.680 18.115 ;
        RECT 47.930 16.955 48.680 17.125 ;
        RECT 47.930 16.665 48.185 16.955 ;
        RECT 48.355 16.405 48.685 16.785 ;
        RECT 48.855 16.665 49.025 18.785 ;
        RECT 49.195 17.985 49.520 18.770 ;
        RECT 49.690 18.495 49.940 18.955 ;
        RECT 50.110 18.455 50.360 18.785 ;
        RECT 50.575 18.455 51.255 18.785 ;
        RECT 50.110 18.325 50.280 18.455 ;
        RECT 49.885 18.155 50.280 18.325 ;
        RECT 49.255 16.935 49.715 17.985 ;
        RECT 49.885 16.795 50.055 18.155 ;
        RECT 50.450 17.895 50.915 18.285 ;
        RECT 50.225 17.085 50.575 17.705 ;
        RECT 50.745 17.305 50.915 17.895 ;
        RECT 51.085 17.675 51.255 18.455 ;
        RECT 51.425 18.355 51.595 18.695 ;
        RECT 51.830 18.525 52.160 18.955 ;
        RECT 52.330 18.355 52.500 18.695 ;
        RECT 52.795 18.495 53.165 18.955 ;
        RECT 51.425 18.185 52.500 18.355 ;
        RECT 53.335 18.325 53.505 18.785 ;
        RECT 53.740 18.445 54.610 18.785 ;
        RECT 54.780 18.495 55.030 18.955 ;
        RECT 52.945 18.155 53.505 18.325 ;
        RECT 52.945 18.015 53.115 18.155 ;
        RECT 51.615 17.845 53.115 18.015 ;
        RECT 53.810 17.985 54.270 18.275 ;
        RECT 51.085 17.505 52.775 17.675 ;
        RECT 50.745 17.085 51.100 17.305 ;
        RECT 51.270 16.795 51.440 17.505 ;
        RECT 51.645 17.085 52.435 17.335 ;
        RECT 52.605 17.325 52.775 17.505 ;
        RECT 52.945 17.155 53.115 17.845 ;
        RECT 49.385 16.405 49.715 16.765 ;
        RECT 49.885 16.625 50.380 16.795 ;
        RECT 50.585 16.625 51.440 16.795 ;
        RECT 52.315 16.405 52.645 16.865 ;
        RECT 52.855 16.765 53.115 17.155 ;
        RECT 53.305 17.975 54.270 17.985 ;
        RECT 54.440 18.065 54.610 18.445 ;
        RECT 55.200 18.405 55.370 18.695 ;
        RECT 55.550 18.575 55.880 18.955 ;
        RECT 55.200 18.235 56.000 18.405 ;
        RECT 53.305 17.815 53.980 17.975 ;
        RECT 54.440 17.895 55.660 18.065 ;
        RECT 53.305 17.025 53.515 17.815 ;
        RECT 54.440 17.805 54.610 17.895 ;
        RECT 53.685 17.025 54.035 17.645 ;
        RECT 54.205 17.635 54.610 17.805 ;
        RECT 54.205 16.855 54.375 17.635 ;
        RECT 54.545 17.185 54.765 17.465 ;
        RECT 54.945 17.355 55.485 17.725 ;
        RECT 55.830 17.645 56.000 18.235 ;
        RECT 56.220 17.815 56.525 18.955 ;
        RECT 56.695 17.765 56.950 18.645 ;
        RECT 55.830 17.615 56.570 17.645 ;
        RECT 54.545 17.015 55.075 17.185 ;
        RECT 52.855 16.595 53.205 16.765 ;
        RECT 53.425 16.575 54.375 16.855 ;
        RECT 54.545 16.405 54.735 16.845 ;
        RECT 54.905 16.785 55.075 17.015 ;
        RECT 55.245 16.955 55.485 17.355 ;
        RECT 55.655 17.315 56.570 17.615 ;
        RECT 55.655 17.140 55.980 17.315 ;
        RECT 55.655 16.785 55.975 17.140 ;
        RECT 56.740 17.115 56.950 17.765 ;
        RECT 54.905 16.615 55.975 16.785 ;
        RECT 56.220 16.405 56.525 16.865 ;
        RECT 56.695 16.585 56.950 17.115 ;
        RECT 57.125 18.085 57.400 18.785 ;
        RECT 57.570 18.410 57.825 18.955 ;
        RECT 57.995 18.445 58.475 18.785 ;
        RECT 58.650 18.400 59.255 18.955 ;
        RECT 58.640 18.300 59.255 18.400 ;
        RECT 58.640 18.275 58.825 18.300 ;
        RECT 57.125 17.055 57.295 18.085 ;
        RECT 57.570 17.955 58.325 18.205 ;
        RECT 58.495 18.030 58.825 18.275 ;
        RECT 59.430 18.285 59.685 18.785 ;
        RECT 59.855 18.455 60.185 18.955 ;
        RECT 57.570 17.920 58.340 17.955 ;
        RECT 57.570 17.910 58.355 17.920 ;
        RECT 57.465 17.895 58.360 17.910 ;
        RECT 57.465 17.880 58.380 17.895 ;
        RECT 57.465 17.870 58.400 17.880 ;
        RECT 57.465 17.860 58.425 17.870 ;
        RECT 57.465 17.830 58.495 17.860 ;
        RECT 57.465 17.800 58.515 17.830 ;
        RECT 57.465 17.770 58.535 17.800 ;
        RECT 57.465 17.745 58.565 17.770 ;
        RECT 57.465 17.710 58.600 17.745 ;
        RECT 57.465 17.705 58.630 17.710 ;
        RECT 57.465 17.310 57.695 17.705 ;
        RECT 58.240 17.700 58.630 17.705 ;
        RECT 58.265 17.690 58.630 17.700 ;
        RECT 58.280 17.685 58.630 17.690 ;
        RECT 58.295 17.680 58.630 17.685 ;
        RECT 58.995 17.680 59.255 18.130 ;
        RECT 59.430 18.115 60.180 18.285 ;
        RECT 58.295 17.675 59.255 17.680 ;
        RECT 58.305 17.665 59.255 17.675 ;
        RECT 58.315 17.660 59.255 17.665 ;
        RECT 58.325 17.650 59.255 17.660 ;
        RECT 58.330 17.640 59.255 17.650 ;
        RECT 58.335 17.635 59.255 17.640 ;
        RECT 58.345 17.620 59.255 17.635 ;
        RECT 58.350 17.605 59.255 17.620 ;
        RECT 58.360 17.580 59.255 17.605 ;
        RECT 57.865 17.110 58.195 17.535 ;
        RECT 57.125 16.575 57.385 17.055 ;
        RECT 57.555 16.405 57.805 16.945 ;
        RECT 57.975 16.625 58.195 17.110 ;
        RECT 58.365 17.510 59.255 17.580 ;
        RECT 58.365 16.785 58.535 17.510 ;
        RECT 58.705 16.955 59.255 17.340 ;
        RECT 59.430 17.295 59.780 17.945 ;
        RECT 59.950 17.125 60.180 18.115 ;
        RECT 59.430 16.955 60.180 17.125 ;
        RECT 58.365 16.615 59.255 16.785 ;
        RECT 59.430 16.665 59.685 16.955 ;
        RECT 59.855 16.405 60.185 16.785 ;
        RECT 60.355 16.665 60.525 18.785 ;
        RECT 60.695 17.985 61.020 18.770 ;
        RECT 61.190 18.495 61.440 18.955 ;
        RECT 61.610 18.455 61.860 18.785 ;
        RECT 62.075 18.455 62.755 18.785 ;
        RECT 61.610 18.325 61.780 18.455 ;
        RECT 61.385 18.155 61.780 18.325 ;
        RECT 60.755 16.935 61.215 17.985 ;
        RECT 61.385 16.795 61.555 18.155 ;
        RECT 61.950 17.895 62.415 18.285 ;
        RECT 61.725 17.085 62.075 17.705 ;
        RECT 62.245 17.305 62.415 17.895 ;
        RECT 62.585 17.675 62.755 18.455 ;
        RECT 62.925 18.355 63.095 18.695 ;
        RECT 63.330 18.525 63.660 18.955 ;
        RECT 63.830 18.355 64.000 18.695 ;
        RECT 64.295 18.495 64.665 18.955 ;
        RECT 62.925 18.185 64.000 18.355 ;
        RECT 64.835 18.325 65.005 18.785 ;
        RECT 65.240 18.445 66.110 18.785 ;
        RECT 66.280 18.495 66.530 18.955 ;
        RECT 64.445 18.155 65.005 18.325 ;
        RECT 64.445 18.015 64.615 18.155 ;
        RECT 63.115 17.845 64.615 18.015 ;
        RECT 65.310 17.985 65.770 18.275 ;
        RECT 62.585 17.505 64.275 17.675 ;
        RECT 62.245 17.085 62.600 17.305 ;
        RECT 62.770 16.795 62.940 17.505 ;
        RECT 63.145 17.085 63.935 17.335 ;
        RECT 64.105 17.325 64.275 17.505 ;
        RECT 64.445 17.155 64.615 17.845 ;
        RECT 60.885 16.405 61.215 16.765 ;
        RECT 61.385 16.625 61.880 16.795 ;
        RECT 62.085 16.625 62.940 16.795 ;
        RECT 63.815 16.405 64.145 16.865 ;
        RECT 64.355 16.765 64.615 17.155 ;
        RECT 64.805 17.975 65.770 17.985 ;
        RECT 65.940 18.065 66.110 18.445 ;
        RECT 66.700 18.405 66.870 18.695 ;
        RECT 67.050 18.575 67.380 18.955 ;
        RECT 66.700 18.235 67.500 18.405 ;
        RECT 64.805 17.815 65.480 17.975 ;
        RECT 65.940 17.895 67.160 18.065 ;
        RECT 64.805 17.025 65.015 17.815 ;
        RECT 65.940 17.805 66.110 17.895 ;
        RECT 65.185 17.025 65.535 17.645 ;
        RECT 65.705 17.635 66.110 17.805 ;
        RECT 65.705 16.855 65.875 17.635 ;
        RECT 66.045 17.185 66.265 17.465 ;
        RECT 66.445 17.355 66.985 17.725 ;
        RECT 67.330 17.615 67.500 18.235 ;
        RECT 67.675 17.895 67.845 18.955 ;
        RECT 68.055 17.945 68.345 18.785 ;
        RECT 68.515 18.115 68.685 18.955 ;
        RECT 68.895 17.945 69.145 18.785 ;
        RECT 69.355 18.115 69.525 18.955 ;
        RECT 68.055 17.775 69.780 17.945 ;
        RECT 70.005 17.790 70.295 18.955 ;
        RECT 70.525 17.815 70.735 18.955 ;
        RECT 70.905 17.805 71.235 18.785 ;
        RECT 71.405 17.815 71.635 18.955 ;
        RECT 71.885 17.815 72.115 18.955 ;
        RECT 72.285 17.805 72.615 18.785 ;
        RECT 72.785 17.815 72.995 18.955 ;
        RECT 73.225 18.520 78.570 18.955 ;
        RECT 78.745 18.520 84.090 18.955 ;
        RECT 84.265 18.520 89.610 18.955 ;
        RECT 89.785 18.520 95.130 18.955 ;
        RECT 66.045 17.015 66.575 17.185 ;
        RECT 64.355 16.595 64.705 16.765 ;
        RECT 64.925 16.575 65.875 16.855 ;
        RECT 66.045 16.405 66.235 16.845 ;
        RECT 66.405 16.785 66.575 17.015 ;
        RECT 66.745 16.955 66.985 17.355 ;
        RECT 67.155 17.605 67.500 17.615 ;
        RECT 67.155 17.395 69.185 17.605 ;
        RECT 67.155 17.140 67.480 17.395 ;
        RECT 69.370 17.225 69.780 17.775 ;
        RECT 67.155 16.785 67.475 17.140 ;
        RECT 66.405 16.615 67.475 16.785 ;
        RECT 67.675 16.405 67.845 17.215 ;
        RECT 68.015 17.055 69.780 17.225 ;
        RECT 68.015 16.575 68.345 17.055 ;
        RECT 68.515 16.405 68.685 16.875 ;
        RECT 68.855 16.575 69.185 17.055 ;
        RECT 69.355 16.405 69.525 16.875 ;
        RECT 70.005 16.405 70.295 17.130 ;
        RECT 70.525 16.405 70.735 17.225 ;
        RECT 70.905 17.205 71.155 17.805 ;
        RECT 71.325 17.395 71.655 17.645 ;
        RECT 71.865 17.395 72.195 17.645 ;
        RECT 70.905 16.575 71.235 17.205 ;
        RECT 71.405 16.405 71.635 17.225 ;
        RECT 71.885 16.405 72.115 17.225 ;
        RECT 72.365 17.205 72.615 17.805 ;
        RECT 72.285 16.575 72.615 17.205 ;
        RECT 72.785 16.405 72.995 17.225 ;
        RECT 74.810 16.950 75.150 17.780 ;
        RECT 76.630 17.270 76.980 18.520 ;
        RECT 80.330 16.950 80.670 17.780 ;
        RECT 82.150 17.270 82.500 18.520 ;
        RECT 85.850 16.950 86.190 17.780 ;
        RECT 87.670 17.270 88.020 18.520 ;
        RECT 91.370 16.950 91.710 17.780 ;
        RECT 93.190 17.270 93.540 18.520 ;
        RECT 95.765 17.790 96.055 18.955 ;
        RECT 96.225 18.520 101.570 18.955 ;
        RECT 101.745 18.520 107.090 18.955 ;
        RECT 73.225 16.405 78.570 16.950 ;
        RECT 78.745 16.405 84.090 16.950 ;
        RECT 84.265 16.405 89.610 16.950 ;
        RECT 89.785 16.405 95.130 16.950 ;
        RECT 95.765 16.405 96.055 17.130 ;
        RECT 97.810 16.950 98.150 17.780 ;
        RECT 99.630 17.270 99.980 18.520 ;
        RECT 103.330 16.950 103.670 17.780 ;
        RECT 105.150 17.270 105.500 18.520 ;
        RECT 107.265 17.865 110.775 18.955 ;
        RECT 110.945 17.865 112.155 18.955 ;
        RECT 107.265 17.175 108.915 17.695 ;
        RECT 109.085 17.345 110.775 17.865 ;
        RECT 96.225 16.405 101.570 16.950 ;
        RECT 101.745 16.405 107.090 16.950 ;
        RECT 107.265 16.405 110.775 17.175 ;
        RECT 110.945 17.155 111.465 17.695 ;
        RECT 111.635 17.325 112.155 17.865 ;
        RECT 112.325 17.865 113.535 18.955 ;
        RECT 112.325 17.325 112.845 17.865 ;
        RECT 113.015 17.155 113.535 17.695 ;
        RECT 110.945 16.405 112.155 17.155 ;
        RECT 112.325 16.405 113.535 17.155 ;
        RECT 5.520 16.235 113.620 16.405 ;
        RECT 5.605 15.485 6.815 16.235 ;
        RECT 6.985 15.690 12.330 16.235 ;
        RECT 12.505 15.690 17.850 16.235 ;
        RECT 18.025 15.690 23.370 16.235 ;
        RECT 23.545 15.690 28.890 16.235 ;
        RECT 5.605 14.945 6.125 15.485 ;
        RECT 6.295 14.775 6.815 15.315 ;
        RECT 8.570 14.860 8.910 15.690 ;
        RECT 5.605 13.685 6.815 14.775 ;
        RECT 10.390 14.120 10.740 15.370 ;
        RECT 14.090 14.860 14.430 15.690 ;
        RECT 15.910 14.120 16.260 15.370 ;
        RECT 19.610 14.860 19.950 15.690 ;
        RECT 21.430 14.120 21.780 15.370 ;
        RECT 25.130 14.860 25.470 15.690 ;
        RECT 29.065 15.465 30.735 16.235 ;
        RECT 31.365 15.510 31.655 16.235 ;
        RECT 31.825 15.690 37.170 16.235 ;
        RECT 37.345 15.690 42.690 16.235 ;
        RECT 26.950 14.120 27.300 15.370 ;
        RECT 29.065 14.945 29.815 15.465 ;
        RECT 29.985 14.775 30.735 15.295 ;
        RECT 33.410 14.860 33.750 15.690 ;
        RECT 6.985 13.685 12.330 14.120 ;
        RECT 12.505 13.685 17.850 14.120 ;
        RECT 18.025 13.685 23.370 14.120 ;
        RECT 23.545 13.685 28.890 14.120 ;
        RECT 29.065 13.685 30.735 14.775 ;
        RECT 31.365 13.685 31.655 14.850 ;
        RECT 35.230 14.120 35.580 15.370 ;
        RECT 38.930 14.860 39.270 15.690 ;
        RECT 42.865 15.465 45.455 16.235 ;
        RECT 46.090 15.685 46.345 15.975 ;
        RECT 46.515 15.855 46.845 16.235 ;
        RECT 46.090 15.515 46.840 15.685 ;
        RECT 40.750 14.120 41.100 15.370 ;
        RECT 42.865 14.945 44.075 15.465 ;
        RECT 44.245 14.775 45.455 15.295 ;
        RECT 31.825 13.685 37.170 14.120 ;
        RECT 37.345 13.685 42.690 14.120 ;
        RECT 42.865 13.685 45.455 14.775 ;
        RECT 46.090 14.695 46.440 15.345 ;
        RECT 46.610 14.525 46.840 15.515 ;
        RECT 46.090 14.355 46.840 14.525 ;
        RECT 46.090 13.855 46.345 14.355 ;
        RECT 46.515 13.685 46.845 14.185 ;
        RECT 47.015 13.855 47.185 15.975 ;
        RECT 47.545 15.875 47.875 16.235 ;
        RECT 48.045 15.845 48.540 16.015 ;
        RECT 48.745 15.845 49.600 16.015 ;
        RECT 47.415 14.655 47.875 15.705 ;
        RECT 47.355 13.870 47.680 14.655 ;
        RECT 48.045 14.485 48.215 15.845 ;
        RECT 48.385 14.935 48.735 15.555 ;
        RECT 48.905 15.335 49.260 15.555 ;
        RECT 48.905 14.745 49.075 15.335 ;
        RECT 49.430 15.135 49.600 15.845 ;
        RECT 50.475 15.775 50.805 16.235 ;
        RECT 51.015 15.875 51.365 16.045 ;
        RECT 49.805 15.305 50.595 15.555 ;
        RECT 51.015 15.485 51.275 15.875 ;
        RECT 51.585 15.785 52.535 16.065 ;
        RECT 52.705 15.795 52.895 16.235 ;
        RECT 53.065 15.855 54.135 16.025 ;
        RECT 50.765 15.135 50.935 15.315 ;
        RECT 48.045 14.315 48.440 14.485 ;
        RECT 48.610 14.355 49.075 14.745 ;
        RECT 49.245 14.965 50.935 15.135 ;
        RECT 48.270 14.185 48.440 14.315 ;
        RECT 49.245 14.185 49.415 14.965 ;
        RECT 51.105 14.795 51.275 15.485 ;
        RECT 49.775 14.625 51.275 14.795 ;
        RECT 51.465 14.825 51.675 15.615 ;
        RECT 51.845 14.995 52.195 15.615 ;
        RECT 52.365 15.005 52.535 15.785 ;
        RECT 53.065 15.625 53.235 15.855 ;
        RECT 52.705 15.455 53.235 15.625 ;
        RECT 52.705 15.175 52.925 15.455 ;
        RECT 53.405 15.285 53.645 15.685 ;
        RECT 52.365 14.835 52.770 15.005 ;
        RECT 53.105 14.915 53.645 15.285 ;
        RECT 53.815 15.500 54.135 15.855 ;
        RECT 54.380 15.775 54.685 16.235 ;
        RECT 54.855 15.525 55.110 16.055 ;
        RECT 53.815 15.325 54.140 15.500 ;
        RECT 53.815 15.025 54.730 15.325 ;
        RECT 53.990 14.995 54.730 15.025 ;
        RECT 51.465 14.665 52.140 14.825 ;
        RECT 52.600 14.745 52.770 14.835 ;
        RECT 51.465 14.655 52.430 14.665 ;
        RECT 51.105 14.485 51.275 14.625 ;
        RECT 47.850 13.685 48.100 14.145 ;
        RECT 48.270 13.855 48.520 14.185 ;
        RECT 48.735 13.855 49.415 14.185 ;
        RECT 49.585 14.285 50.660 14.455 ;
        RECT 51.105 14.315 51.665 14.485 ;
        RECT 51.970 14.365 52.430 14.655 ;
        RECT 52.600 14.575 53.820 14.745 ;
        RECT 49.585 13.945 49.755 14.285 ;
        RECT 49.990 13.685 50.320 14.115 ;
        RECT 50.490 13.945 50.660 14.285 ;
        RECT 50.955 13.685 51.325 14.145 ;
        RECT 51.495 13.855 51.665 14.315 ;
        RECT 52.600 14.195 52.770 14.575 ;
        RECT 53.990 14.405 54.160 14.995 ;
        RECT 54.900 14.875 55.110 15.525 ;
        RECT 55.345 15.415 55.555 16.235 ;
        RECT 55.725 15.435 56.055 16.065 ;
        RECT 51.900 13.855 52.770 14.195 ;
        RECT 53.360 14.235 54.160 14.405 ;
        RECT 52.940 13.685 53.190 14.145 ;
        RECT 53.360 13.945 53.530 14.235 ;
        RECT 53.710 13.685 54.040 14.065 ;
        RECT 54.380 13.685 54.685 14.825 ;
        RECT 54.855 13.995 55.110 14.875 ;
        RECT 55.725 14.835 55.975 15.435 ;
        RECT 56.225 15.415 56.455 16.235 ;
        RECT 57.125 15.510 57.415 16.235 ;
        RECT 57.585 15.465 60.175 16.235 ;
        RECT 60.345 15.855 61.235 16.025 ;
        RECT 56.145 14.995 56.475 15.245 ;
        RECT 57.585 14.945 58.795 15.465 ;
        RECT 60.345 15.300 60.895 15.685 ;
        RECT 55.345 13.685 55.555 14.825 ;
        RECT 55.725 13.855 56.055 14.835 ;
        RECT 56.225 13.685 56.455 14.825 ;
        RECT 57.125 13.685 57.415 14.850 ;
        RECT 58.965 14.775 60.175 15.295 ;
        RECT 61.065 15.130 61.235 15.855 ;
        RECT 57.585 13.685 60.175 14.775 ;
        RECT 60.345 15.060 61.235 15.130 ;
        RECT 61.405 15.555 61.625 16.015 ;
        RECT 61.795 15.695 62.045 16.235 ;
        RECT 62.215 15.585 62.475 16.065 ;
        RECT 61.405 15.530 61.655 15.555 ;
        RECT 61.405 15.105 61.735 15.530 ;
        RECT 60.345 15.035 61.240 15.060 ;
        RECT 60.345 15.020 61.250 15.035 ;
        RECT 60.345 15.005 61.255 15.020 ;
        RECT 60.345 15.000 61.265 15.005 ;
        RECT 60.345 14.990 61.270 15.000 ;
        RECT 60.345 14.980 61.275 14.990 ;
        RECT 60.345 14.975 61.285 14.980 ;
        RECT 60.345 14.965 61.295 14.975 ;
        RECT 60.345 14.960 61.305 14.965 ;
        RECT 60.345 14.510 60.605 14.960 ;
        RECT 60.970 14.955 61.305 14.960 ;
        RECT 60.970 14.950 61.320 14.955 ;
        RECT 60.970 14.940 61.335 14.950 ;
        RECT 60.970 14.935 61.360 14.940 ;
        RECT 61.905 14.935 62.135 15.330 ;
        RECT 60.970 14.930 62.135 14.935 ;
        RECT 61.000 14.895 62.135 14.930 ;
        RECT 61.035 14.870 62.135 14.895 ;
        RECT 61.065 14.840 62.135 14.870 ;
        RECT 61.085 14.810 62.135 14.840 ;
        RECT 61.105 14.780 62.135 14.810 ;
        RECT 61.175 14.770 62.135 14.780 ;
        RECT 61.200 14.760 62.135 14.770 ;
        RECT 61.220 14.745 62.135 14.760 ;
        RECT 61.240 14.730 62.135 14.745 ;
        RECT 61.245 14.720 62.030 14.730 ;
        RECT 61.260 14.685 62.030 14.720 ;
        RECT 60.775 14.365 61.105 14.610 ;
        RECT 61.275 14.435 62.030 14.685 ;
        RECT 62.305 14.555 62.475 15.585 ;
        RECT 60.775 14.340 60.960 14.365 ;
        RECT 60.345 14.240 60.960 14.340 ;
        RECT 60.345 13.685 60.950 14.240 ;
        RECT 61.125 13.855 61.605 14.195 ;
        RECT 61.775 13.685 62.030 14.230 ;
        RECT 62.200 13.855 62.475 14.555 ;
        RECT 62.645 15.560 62.905 16.065 ;
        RECT 63.085 15.855 63.415 16.235 ;
        RECT 63.595 15.685 63.765 16.065 ;
        RECT 64.025 15.690 69.370 16.235 ;
        RECT 69.545 15.690 74.890 16.235 ;
        RECT 75.065 15.690 80.410 16.235 ;
        RECT 62.645 14.760 62.815 15.560 ;
        RECT 63.100 15.515 63.765 15.685 ;
        RECT 63.100 15.260 63.270 15.515 ;
        RECT 62.985 14.930 63.270 15.260 ;
        RECT 63.505 14.965 63.835 15.335 ;
        RECT 63.100 14.785 63.270 14.930 ;
        RECT 65.610 14.860 65.950 15.690 ;
        RECT 62.645 13.855 62.915 14.760 ;
        RECT 63.100 14.615 63.765 14.785 ;
        RECT 63.085 13.685 63.415 14.445 ;
        RECT 63.595 13.855 63.765 14.615 ;
        RECT 67.430 14.120 67.780 15.370 ;
        RECT 71.130 14.860 71.470 15.690 ;
        RECT 72.950 14.120 73.300 15.370 ;
        RECT 76.650 14.860 76.990 15.690 ;
        RECT 80.585 15.465 82.255 16.235 ;
        RECT 82.885 15.510 83.175 16.235 ;
        RECT 83.345 15.690 88.690 16.235 ;
        RECT 88.865 15.690 94.210 16.235 ;
        RECT 94.385 15.690 99.730 16.235 ;
        RECT 99.905 15.690 105.250 16.235 ;
        RECT 78.470 14.120 78.820 15.370 ;
        RECT 80.585 14.945 81.335 15.465 ;
        RECT 81.505 14.775 82.255 15.295 ;
        RECT 84.930 14.860 85.270 15.690 ;
        RECT 64.025 13.685 69.370 14.120 ;
        RECT 69.545 13.685 74.890 14.120 ;
        RECT 75.065 13.685 80.410 14.120 ;
        RECT 80.585 13.685 82.255 14.775 ;
        RECT 82.885 13.685 83.175 14.850 ;
        RECT 86.750 14.120 87.100 15.370 ;
        RECT 90.450 14.860 90.790 15.690 ;
        RECT 92.270 14.120 92.620 15.370 ;
        RECT 95.970 14.860 96.310 15.690 ;
        RECT 97.790 14.120 98.140 15.370 ;
        RECT 101.490 14.860 101.830 15.690 ;
        RECT 105.425 15.465 108.015 16.235 ;
        RECT 108.645 15.510 108.935 16.235 ;
        RECT 109.105 15.465 111.695 16.235 ;
        RECT 112.325 15.485 113.535 16.235 ;
        RECT 103.310 14.120 103.660 15.370 ;
        RECT 105.425 14.945 106.635 15.465 ;
        RECT 106.805 14.775 108.015 15.295 ;
        RECT 109.105 14.945 110.315 15.465 ;
        RECT 83.345 13.685 88.690 14.120 ;
        RECT 88.865 13.685 94.210 14.120 ;
        RECT 94.385 13.685 99.730 14.120 ;
        RECT 99.905 13.685 105.250 14.120 ;
        RECT 105.425 13.685 108.015 14.775 ;
        RECT 108.645 13.685 108.935 14.850 ;
        RECT 110.485 14.775 111.695 15.295 ;
        RECT 109.105 13.685 111.695 14.775 ;
        RECT 112.325 14.775 112.845 15.315 ;
        RECT 113.015 14.945 113.535 15.485 ;
        RECT 112.325 13.685 113.535 14.775 ;
        RECT 5.520 13.515 113.620 13.685 ;
        RECT 5.605 12.425 6.815 13.515 ;
        RECT 6.985 13.080 12.330 13.515 ;
        RECT 12.505 13.080 17.850 13.515 ;
        RECT 5.605 11.715 6.125 12.255 ;
        RECT 6.295 11.885 6.815 12.425 ;
        RECT 5.605 10.965 6.815 11.715 ;
        RECT 8.570 11.510 8.910 12.340 ;
        RECT 10.390 11.830 10.740 13.080 ;
        RECT 14.090 11.510 14.430 12.340 ;
        RECT 15.910 11.830 16.260 13.080 ;
        RECT 18.485 12.350 18.775 13.515 ;
        RECT 18.945 13.080 24.290 13.515 ;
        RECT 24.465 13.080 29.810 13.515 ;
        RECT 6.985 10.965 12.330 11.510 ;
        RECT 12.505 10.965 17.850 11.510 ;
        RECT 18.485 10.965 18.775 11.690 ;
        RECT 20.530 11.510 20.870 12.340 ;
        RECT 22.350 11.830 22.700 13.080 ;
        RECT 26.050 11.510 26.390 12.340 ;
        RECT 27.870 11.830 28.220 13.080 ;
        RECT 29.985 12.425 31.195 13.515 ;
        RECT 29.985 11.715 30.505 12.255 ;
        RECT 30.675 11.885 31.195 12.425 ;
        RECT 31.365 12.350 31.655 13.515 ;
        RECT 31.825 13.080 37.170 13.515 ;
        RECT 37.345 13.080 42.690 13.515 ;
        RECT 18.945 10.965 24.290 11.510 ;
        RECT 24.465 10.965 29.810 11.510 ;
        RECT 29.985 10.965 31.195 11.715 ;
        RECT 31.365 10.965 31.655 11.690 ;
        RECT 33.410 11.510 33.750 12.340 ;
        RECT 35.230 11.830 35.580 13.080 ;
        RECT 38.930 11.510 39.270 12.340 ;
        RECT 40.750 11.830 41.100 13.080 ;
        RECT 42.865 12.425 44.075 13.515 ;
        RECT 42.865 11.715 43.385 12.255 ;
        RECT 43.555 11.885 44.075 12.425 ;
        RECT 44.245 12.350 44.535 13.515 ;
        RECT 44.705 13.080 50.050 13.515 ;
        RECT 50.225 13.080 55.570 13.515 ;
        RECT 31.825 10.965 37.170 11.510 ;
        RECT 37.345 10.965 42.690 11.510 ;
        RECT 42.865 10.965 44.075 11.715 ;
        RECT 44.245 10.965 44.535 11.690 ;
        RECT 46.290 11.510 46.630 12.340 ;
        RECT 48.110 11.830 48.460 13.080 ;
        RECT 51.810 11.510 52.150 12.340 ;
        RECT 53.630 11.830 53.980 13.080 ;
        RECT 55.745 12.425 56.955 13.515 ;
        RECT 55.745 11.715 56.265 12.255 ;
        RECT 56.435 11.885 56.955 12.425 ;
        RECT 57.125 12.350 57.415 13.515 ;
        RECT 57.585 13.080 62.930 13.515 ;
        RECT 63.105 13.080 68.450 13.515 ;
        RECT 44.705 10.965 50.050 11.510 ;
        RECT 50.225 10.965 55.570 11.510 ;
        RECT 55.745 10.965 56.955 11.715 ;
        RECT 57.125 10.965 57.415 11.690 ;
        RECT 59.170 11.510 59.510 12.340 ;
        RECT 60.990 11.830 61.340 13.080 ;
        RECT 64.690 11.510 65.030 12.340 ;
        RECT 66.510 11.830 66.860 13.080 ;
        RECT 68.625 12.425 69.835 13.515 ;
        RECT 68.625 11.715 69.145 12.255 ;
        RECT 69.315 11.885 69.835 12.425 ;
        RECT 70.005 12.350 70.295 13.515 ;
        RECT 70.465 13.080 75.810 13.515 ;
        RECT 75.985 13.080 81.330 13.515 ;
        RECT 57.585 10.965 62.930 11.510 ;
        RECT 63.105 10.965 68.450 11.510 ;
        RECT 68.625 10.965 69.835 11.715 ;
        RECT 70.005 10.965 70.295 11.690 ;
        RECT 72.050 11.510 72.390 12.340 ;
        RECT 73.870 11.830 74.220 13.080 ;
        RECT 77.570 11.510 77.910 12.340 ;
        RECT 79.390 11.830 79.740 13.080 ;
        RECT 81.505 12.425 82.715 13.515 ;
        RECT 81.505 11.715 82.025 12.255 ;
        RECT 82.195 11.885 82.715 12.425 ;
        RECT 82.885 12.350 83.175 13.515 ;
        RECT 83.345 13.080 88.690 13.515 ;
        RECT 88.865 13.080 94.210 13.515 ;
        RECT 70.465 10.965 75.810 11.510 ;
        RECT 75.985 10.965 81.330 11.510 ;
        RECT 81.505 10.965 82.715 11.715 ;
        RECT 82.885 10.965 83.175 11.690 ;
        RECT 84.930 11.510 85.270 12.340 ;
        RECT 86.750 11.830 87.100 13.080 ;
        RECT 90.450 11.510 90.790 12.340 ;
        RECT 92.270 11.830 92.620 13.080 ;
        RECT 94.385 12.425 95.595 13.515 ;
        RECT 94.385 11.715 94.905 12.255 ;
        RECT 95.075 11.885 95.595 12.425 ;
        RECT 95.765 12.350 96.055 13.515 ;
        RECT 96.225 13.080 101.570 13.515 ;
        RECT 101.745 13.080 107.090 13.515 ;
        RECT 83.345 10.965 88.690 11.510 ;
        RECT 88.865 10.965 94.210 11.510 ;
        RECT 94.385 10.965 95.595 11.715 ;
        RECT 95.765 10.965 96.055 11.690 ;
        RECT 97.810 11.510 98.150 12.340 ;
        RECT 99.630 11.830 99.980 13.080 ;
        RECT 103.330 11.510 103.670 12.340 ;
        RECT 105.150 11.830 105.500 13.080 ;
        RECT 107.265 12.425 108.475 13.515 ;
        RECT 107.265 11.715 107.785 12.255 ;
        RECT 107.955 11.885 108.475 12.425 ;
        RECT 108.645 12.350 108.935 13.515 ;
        RECT 109.105 12.425 111.695 13.515 ;
        RECT 109.105 11.735 110.315 12.255 ;
        RECT 110.485 11.905 111.695 12.425 ;
        RECT 112.325 12.425 113.535 13.515 ;
        RECT 112.325 11.885 112.845 12.425 ;
        RECT 96.225 10.965 101.570 11.510 ;
        RECT 101.745 10.965 107.090 11.510 ;
        RECT 107.265 10.965 108.475 11.715 ;
        RECT 108.645 10.965 108.935 11.690 ;
        RECT 109.105 10.965 111.695 11.735 ;
        RECT 113.015 11.715 113.535 12.255 ;
        RECT 112.325 10.965 113.535 11.715 ;
        RECT 5.520 10.795 113.620 10.965 ;
      LAYER met1 ;
        RECT 5.520 116.720 113.620 117.200 ;
        RECT 31.825 116.520 32.115 116.565 ;
        RECT 32.730 116.520 33.050 116.580 ;
        RECT 31.825 116.380 33.050 116.520 ;
        RECT 31.825 116.335 32.115 116.380 ;
        RECT 32.730 116.320 33.050 116.380 ;
        RECT 108.185 116.520 108.475 116.565 ;
        RECT 116.450 116.520 116.770 116.580 ;
        RECT 108.185 116.380 116.770 116.520 ;
        RECT 108.185 116.335 108.475 116.380 ;
        RECT 116.450 116.320 116.770 116.380 ;
        RECT 34.685 116.180 34.975 116.225 ;
        RECT 37.805 116.180 38.095 116.225 ;
        RECT 39.695 116.180 39.985 116.225 ;
        RECT 34.685 116.040 39.985 116.180 ;
        RECT 34.685 115.995 34.975 116.040 ;
        RECT 37.805 115.995 38.095 116.040 ;
        RECT 39.695 115.995 39.985 116.040 ;
        RECT 100.315 116.180 100.605 116.225 ;
        RECT 102.205 116.180 102.495 116.225 ;
        RECT 105.325 116.180 105.615 116.225 ;
        RECT 100.315 116.040 105.615 116.180 ;
        RECT 100.315 115.995 100.605 116.040 ;
        RECT 102.205 115.995 102.495 116.040 ;
        RECT 105.325 115.995 105.615 116.040 ;
        RECT 35.490 115.840 35.810 115.900 ;
        RECT 39.185 115.840 39.475 115.885 ;
        RECT 104.490 115.840 104.810 115.900 ;
        RECT 35.490 115.700 39.475 115.840 ;
        RECT 35.490 115.640 35.810 115.700 ;
        RECT 39.185 115.655 39.475 115.700 ;
        RECT 97.220 115.700 104.810 115.840 ;
        RECT 1.910 115.500 2.230 115.560 ;
        RECT 6.985 115.500 7.275 115.545 ;
        RECT 33.650 115.520 33.970 115.560 ;
        RECT 1.910 115.360 7.275 115.500 ;
        RECT 1.910 115.300 2.230 115.360 ;
        RECT 6.985 115.315 7.275 115.360 ;
        RECT 33.605 115.300 33.970 115.520 ;
        RECT 34.685 115.500 34.975 115.545 ;
        RECT 38.265 115.500 38.555 115.545 ;
        RECT 40.100 115.500 40.390 115.545 ;
        RECT 34.685 115.360 40.390 115.500 ;
        RECT 34.685 115.315 34.975 115.360 ;
        RECT 38.265 115.315 38.555 115.360 ;
        RECT 40.100 115.315 40.390 115.360 ;
        RECT 40.565 115.500 40.855 115.545 ;
        RECT 41.930 115.500 42.250 115.560 ;
        RECT 40.565 115.360 42.250 115.500 ;
        RECT 40.565 115.315 40.855 115.360 ;
        RECT 41.930 115.300 42.250 115.360 ;
        RECT 51.130 115.500 51.450 115.560 ;
        RECT 52.985 115.500 53.275 115.545 ;
        RECT 51.130 115.360 53.275 115.500 ;
        RECT 51.130 115.300 51.450 115.360 ;
        RECT 52.985 115.315 53.275 115.360 ;
        RECT 81.490 115.500 81.810 115.560 ;
        RECT 97.220 115.545 97.360 115.700 ;
        RECT 104.490 115.640 104.810 115.700 ;
        RECT 84.725 115.500 85.015 115.545 ;
        RECT 90.705 115.500 90.995 115.545 ;
        RECT 97.145 115.500 97.435 115.545 ;
        RECT 81.490 115.360 97.435 115.500 ;
        RECT 81.490 115.300 81.810 115.360 ;
        RECT 84.725 115.315 85.015 115.360 ;
        RECT 90.705 115.315 90.995 115.360 ;
        RECT 97.145 115.315 97.435 115.360 ;
        RECT 97.590 115.500 97.910 115.560 ;
        RECT 99.445 115.500 99.735 115.545 ;
        RECT 97.590 115.360 99.735 115.500 ;
        RECT 97.590 115.300 97.910 115.360 ;
        RECT 99.445 115.315 99.735 115.360 ;
        RECT 99.910 115.500 100.200 115.545 ;
        RECT 101.745 115.500 102.035 115.545 ;
        RECT 105.325 115.500 105.615 115.545 ;
        RECT 99.910 115.360 105.615 115.500 ;
        RECT 99.910 115.315 100.200 115.360 ;
        RECT 101.745 115.315 102.035 115.360 ;
        RECT 105.325 115.315 105.615 115.360 ;
        RECT 33.605 115.205 33.895 115.300 ;
        RECT 33.305 115.160 33.895 115.205 ;
        RECT 36.545 115.160 37.195 115.205 ;
        RECT 57.110 115.160 57.430 115.220 ;
        RECT 33.305 115.020 37.195 115.160 ;
        RECT 33.305 114.975 33.595 115.020 ;
        RECT 36.545 114.975 37.195 115.020 ;
        RECT 45.240 115.020 57.430 115.160 ;
        RECT 7.905 114.820 8.195 114.865 ;
        RECT 45.240 114.820 45.380 115.020 ;
        RECT 57.110 114.960 57.430 115.020 ;
        RECT 100.810 114.960 101.130 115.220 ;
        RECT 106.405 115.205 106.695 115.520 ;
        RECT 103.105 115.160 103.755 115.205 ;
        RECT 106.405 115.160 106.995 115.205 ;
        RECT 107.250 115.160 107.570 115.220 ;
        RECT 103.105 115.020 107.570 115.160 ;
        RECT 103.105 114.975 103.755 115.020 ;
        RECT 106.705 114.975 106.995 115.020 ;
        RECT 107.250 114.960 107.570 115.020 ;
        RECT 7.905 114.680 45.380 114.820 ;
        RECT 7.905 114.635 8.195 114.680 ;
        RECT 51.590 114.620 51.910 114.880 ;
        RECT 52.970 114.820 53.290 114.880 ;
        RECT 53.445 114.820 53.735 114.865 ;
        RECT 52.970 114.680 53.735 114.820 ;
        RECT 52.970 114.620 53.290 114.680 ;
        RECT 53.445 114.635 53.735 114.680 ;
        RECT 85.185 114.820 85.475 114.865 ;
        RECT 87.010 114.820 87.330 114.880 ;
        RECT 85.185 114.680 87.330 114.820 ;
        RECT 85.185 114.635 85.475 114.680 ;
        RECT 87.010 114.620 87.330 114.680 ;
        RECT 90.690 114.820 91.010 114.880 ;
        RECT 91.165 114.820 91.455 114.865 ;
        RECT 90.690 114.680 91.455 114.820 ;
        RECT 90.690 114.620 91.010 114.680 ;
        RECT 91.165 114.635 91.455 114.680 ;
        RECT 97.130 114.820 97.450 114.880 ;
        RECT 97.605 114.820 97.895 114.865 ;
        RECT 97.130 114.680 97.895 114.820 ;
        RECT 97.130 114.620 97.450 114.680 ;
        RECT 97.605 114.635 97.895 114.680 ;
        RECT 5.520 114.000 113.620 114.480 ;
        RECT 10.205 113.800 10.495 113.845 ;
        RECT 14.330 113.800 14.650 113.860 ;
        RECT 10.205 113.660 14.650 113.800 ;
        RECT 10.205 113.615 10.495 113.660 ;
        RECT 14.330 113.600 14.650 113.660 ;
        RECT 26.750 113.800 27.070 113.860 ;
        RECT 29.985 113.800 30.275 113.845 ;
        RECT 26.750 113.660 30.275 113.800 ;
        RECT 26.750 113.600 27.070 113.660 ;
        RECT 29.985 113.615 30.275 113.660 ;
        RECT 44.230 113.800 44.550 113.860 ;
        RECT 47.005 113.800 47.295 113.845 ;
        RECT 44.230 113.660 47.295 113.800 ;
        RECT 44.230 113.600 44.550 113.660 ;
        RECT 47.005 113.615 47.295 113.660 ;
        RECT 56.650 113.600 56.970 113.860 ;
        RECT 68.610 113.800 68.930 113.860 ;
        RECT 70.925 113.800 71.215 113.845 ;
        RECT 68.610 113.660 71.215 113.800 ;
        RECT 68.610 113.600 68.930 113.660 ;
        RECT 70.925 113.615 71.215 113.660 ;
        RECT 74.590 113.800 74.910 113.860 ;
        RECT 80.125 113.800 80.415 113.845 ;
        RECT 74.590 113.660 80.415 113.800 ;
        RECT 74.590 113.600 74.910 113.660 ;
        RECT 80.125 113.615 80.415 113.660 ;
        RECT 86.550 113.800 86.870 113.860 ;
        RECT 92.085 113.800 92.375 113.845 ;
        RECT 86.550 113.660 92.375 113.800 ;
        RECT 86.550 113.600 86.870 113.660 ;
        RECT 92.085 113.615 92.375 113.660 ;
        RECT 100.810 113.800 101.130 113.860 ;
        RECT 101.745 113.800 102.035 113.845 ;
        RECT 100.810 113.660 102.035 113.800 ;
        RECT 100.810 113.600 101.130 113.660 ;
        RECT 101.745 113.615 102.035 113.660 ;
        RECT 107.250 113.600 107.570 113.860 ;
        RECT 11.685 113.460 11.975 113.505 ;
        RECT 14.925 113.460 15.575 113.505 ;
        RECT 18.010 113.460 18.330 113.520 ;
        RECT 11.685 113.320 18.330 113.460 ;
        RECT 11.685 113.275 12.275 113.320 ;
        RECT 14.925 113.275 15.575 113.320 ;
        RECT 11.985 112.960 12.275 113.275 ;
        RECT 18.010 113.260 18.330 113.320 ;
        RECT 24.905 113.460 25.555 113.505 ;
        RECT 28.505 113.460 28.795 113.505 ;
        RECT 29.510 113.460 29.830 113.520 ;
        RECT 24.905 113.320 29.830 113.460 ;
        RECT 24.905 113.275 25.555 113.320 ;
        RECT 28.205 113.275 28.795 113.320 ;
        RECT 13.065 113.120 13.355 113.165 ;
        RECT 16.645 113.120 16.935 113.165 ;
        RECT 18.480 113.120 18.770 113.165 ;
        RECT 13.065 112.980 18.770 113.120 ;
        RECT 13.065 112.935 13.355 112.980 ;
        RECT 16.645 112.935 16.935 112.980 ;
        RECT 18.480 112.935 18.770 112.980 ;
        RECT 21.710 113.120 22.000 113.165 ;
        RECT 23.545 113.120 23.835 113.165 ;
        RECT 27.125 113.120 27.415 113.165 ;
        RECT 21.710 112.980 27.415 113.120 ;
        RECT 21.710 112.935 22.000 112.980 ;
        RECT 23.545 112.935 23.835 112.980 ;
        RECT 27.125 112.935 27.415 112.980 ;
        RECT 28.205 112.960 28.495 113.275 ;
        RECT 29.510 113.260 29.830 113.320 ;
        RECT 41.925 113.460 42.575 113.505 ;
        RECT 44.690 113.460 45.010 113.520 ;
        RECT 45.525 113.460 45.815 113.505 ;
        RECT 41.925 113.320 45.815 113.460 ;
        RECT 41.925 113.275 42.575 113.320 ;
        RECT 44.690 113.260 45.010 113.320 ;
        RECT 45.225 113.275 45.815 113.320 ;
        RECT 51.585 113.460 52.235 113.505 ;
        RECT 52.970 113.460 53.290 113.520 ;
        RECT 55.185 113.460 55.475 113.505 ;
        RECT 51.585 113.320 55.475 113.460 ;
        RECT 51.585 113.275 52.235 113.320 ;
        RECT 38.730 113.120 39.020 113.165 ;
        RECT 40.565 113.120 40.855 113.165 ;
        RECT 44.145 113.120 44.435 113.165 ;
        RECT 38.730 112.980 44.435 113.120 ;
        RECT 38.730 112.935 39.020 112.980 ;
        RECT 40.565 112.935 40.855 112.980 ;
        RECT 44.145 112.935 44.435 112.980 ;
        RECT 45.225 112.960 45.515 113.275 ;
        RECT 52.970 113.260 53.290 113.320 ;
        RECT 54.885 113.275 55.475 113.320 ;
        RECT 65.845 113.460 66.495 113.505 ;
        RECT 69.445 113.460 69.735 113.505 ;
        RECT 65.845 113.320 69.735 113.460 ;
        RECT 65.845 113.275 66.495 113.320 ;
        RECT 69.145 113.275 69.735 113.320 ;
        RECT 75.045 113.460 75.695 113.505 ;
        RECT 75.970 113.460 76.290 113.520 ;
        RECT 87.010 113.505 87.330 113.520 ;
        RECT 78.645 113.460 78.935 113.505 ;
        RECT 75.045 113.320 78.935 113.460 ;
        RECT 75.045 113.275 75.695 113.320 ;
        RECT 48.390 113.120 48.680 113.165 ;
        RECT 50.225 113.120 50.515 113.165 ;
        RECT 53.805 113.120 54.095 113.165 ;
        RECT 48.390 112.980 54.095 113.120 ;
        RECT 48.390 112.935 48.680 112.980 ;
        RECT 50.225 112.935 50.515 112.980 ;
        RECT 53.805 112.935 54.095 112.980 ;
        RECT 54.885 112.960 55.175 113.275 ;
        RECT 69.145 113.180 69.435 113.275 ;
        RECT 75.970 113.260 76.290 113.320 ;
        RECT 78.345 113.275 78.935 113.320 ;
        RECT 87.005 113.460 87.655 113.505 ;
        RECT 90.605 113.460 90.895 113.505 ;
        RECT 87.005 113.320 90.895 113.460 ;
        RECT 87.005 113.275 87.655 113.320 ;
        RECT 90.305 113.275 90.895 113.320 ;
        RECT 96.205 113.460 96.855 113.505 ;
        RECT 97.130 113.460 97.450 113.520 ;
        RECT 99.805 113.460 100.095 113.505 ;
        RECT 96.205 113.320 100.095 113.460 ;
        RECT 96.205 113.275 96.855 113.320 ;
        RECT 62.650 113.120 62.940 113.165 ;
        RECT 64.485 113.120 64.775 113.165 ;
        RECT 68.065 113.120 68.355 113.165 ;
        RECT 62.650 112.980 68.355 113.120 ;
        RECT 62.650 112.935 62.940 112.980 ;
        RECT 64.485 112.935 64.775 112.980 ;
        RECT 68.065 112.935 68.355 112.980 ;
        RECT 69.070 112.960 69.435 113.180 ;
        RECT 71.850 113.120 72.140 113.165 ;
        RECT 73.685 113.120 73.975 113.165 ;
        RECT 77.265 113.120 77.555 113.165 ;
        RECT 71.850 112.980 77.555 113.120 ;
        RECT 69.070 112.920 69.390 112.960 ;
        RECT 71.850 112.935 72.140 112.980 ;
        RECT 73.685 112.935 73.975 112.980 ;
        RECT 77.265 112.935 77.555 112.980 ;
        RECT 78.345 112.960 78.635 113.275 ;
        RECT 87.010 113.260 87.330 113.275 ;
        RECT 81.490 112.920 81.810 113.180 ;
        RECT 83.810 113.120 84.100 113.165 ;
        RECT 85.645 113.120 85.935 113.165 ;
        RECT 89.225 113.120 89.515 113.165 ;
        RECT 83.810 112.980 89.515 113.120 ;
        RECT 83.810 112.935 84.100 112.980 ;
        RECT 85.645 112.935 85.935 112.980 ;
        RECT 89.225 112.935 89.515 112.980 ;
        RECT 90.305 112.960 90.595 113.275 ;
        RECT 97.130 113.260 97.450 113.320 ;
        RECT 99.505 113.275 100.095 113.320 ;
        RECT 93.010 113.120 93.300 113.165 ;
        RECT 94.845 113.120 95.135 113.165 ;
        RECT 98.425 113.120 98.715 113.165 ;
        RECT 93.010 112.980 98.715 113.120 ;
        RECT 93.010 112.935 93.300 112.980 ;
        RECT 94.845 112.935 95.135 112.980 ;
        RECT 98.425 112.935 98.715 112.980 ;
        RECT 99.505 112.960 99.795 113.275 ;
        RECT 102.650 112.920 102.970 113.180 ;
        RECT 104.045 113.120 104.335 113.165 ;
        RECT 104.490 113.120 104.810 113.180 ;
        RECT 106.805 113.120 107.095 113.165 ;
        RECT 104.045 112.980 107.095 113.120 ;
        RECT 104.045 112.935 104.335 112.980 ;
        RECT 104.490 112.920 104.810 112.980 ;
        RECT 106.805 112.935 107.095 112.980 ;
        RECT 17.550 112.580 17.870 112.840 ;
        RECT 18.945 112.780 19.235 112.825 ;
        RECT 20.770 112.780 21.090 112.840 ;
        RECT 21.245 112.780 21.535 112.825 ;
        RECT 18.945 112.640 21.535 112.780 ;
        RECT 18.945 112.595 19.235 112.640 ;
        RECT 20.770 112.580 21.090 112.640 ;
        RECT 21.245 112.595 21.535 112.640 ;
        RECT 22.610 112.580 22.930 112.840 ;
        RECT 38.265 112.780 38.555 112.825 ;
        RECT 39.645 112.780 39.935 112.825 ;
        RECT 42.390 112.780 42.710 112.840 ;
        RECT 38.265 112.640 38.940 112.780 ;
        RECT 38.265 112.595 38.555 112.640 ;
        RECT 13.065 112.440 13.355 112.485 ;
        RECT 16.185 112.440 16.475 112.485 ;
        RECT 18.075 112.440 18.365 112.485 ;
        RECT 13.065 112.300 18.365 112.440 ;
        RECT 13.065 112.255 13.355 112.300 ;
        RECT 16.185 112.255 16.475 112.300 ;
        RECT 18.075 112.255 18.365 112.300 ;
        RECT 22.115 112.440 22.405 112.485 ;
        RECT 24.005 112.440 24.295 112.485 ;
        RECT 27.125 112.440 27.415 112.485 ;
        RECT 22.115 112.300 27.415 112.440 ;
        RECT 22.115 112.255 22.405 112.300 ;
        RECT 24.005 112.255 24.295 112.300 ;
        RECT 27.125 112.255 27.415 112.300 ;
        RECT 38.800 112.100 38.940 112.640 ;
        RECT 39.645 112.640 42.710 112.780 ;
        RECT 39.645 112.595 39.935 112.640 ;
        RECT 42.390 112.580 42.710 112.640 ;
        RECT 46.990 112.780 47.310 112.840 ;
        RECT 47.925 112.780 48.215 112.825 ;
        RECT 46.990 112.640 48.215 112.780 ;
        RECT 46.990 112.580 47.310 112.640 ;
        RECT 47.925 112.595 48.215 112.640 ;
        RECT 49.290 112.580 49.610 112.840 ;
        RECT 62.185 112.595 62.475 112.825 ;
        RECT 39.135 112.440 39.425 112.485 ;
        RECT 41.025 112.440 41.315 112.485 ;
        RECT 44.145 112.440 44.435 112.485 ;
        RECT 39.135 112.300 44.435 112.440 ;
        RECT 39.135 112.255 39.425 112.300 ;
        RECT 41.025 112.255 41.315 112.300 ;
        RECT 44.145 112.255 44.435 112.300 ;
        RECT 48.795 112.440 49.085 112.485 ;
        RECT 50.685 112.440 50.975 112.485 ;
        RECT 53.805 112.440 54.095 112.485 ;
        RECT 48.795 112.300 54.095 112.440 ;
        RECT 48.795 112.255 49.085 112.300 ;
        RECT 50.685 112.255 50.975 112.300 ;
        RECT 53.805 112.255 54.095 112.300 ;
        RECT 62.260 112.160 62.400 112.595 ;
        RECT 63.550 112.580 63.870 112.840 ;
        RECT 71.385 112.595 71.675 112.825 ;
        RECT 63.055 112.440 63.345 112.485 ;
        RECT 64.945 112.440 65.235 112.485 ;
        RECT 68.065 112.440 68.355 112.485 ;
        RECT 71.460 112.440 71.600 112.595 ;
        RECT 72.750 112.580 73.070 112.840 ;
        RECT 83.345 112.780 83.635 112.825 ;
        RECT 77.900 112.640 83.635 112.780 ;
        RECT 63.055 112.300 68.355 112.440 ;
        RECT 63.055 112.255 63.345 112.300 ;
        RECT 64.945 112.255 65.235 112.300 ;
        RECT 68.065 112.255 68.355 112.300 ;
        RECT 68.700 112.300 71.600 112.440 ;
        RECT 41.930 112.100 42.250 112.160 ;
        RECT 38.800 111.960 42.250 112.100 ;
        RECT 41.930 111.900 42.250 111.960 ;
        RECT 62.170 112.100 62.490 112.160 ;
        RECT 68.700 112.100 68.840 112.300 ;
        RECT 62.170 111.960 68.840 112.100 ;
        RECT 71.460 112.100 71.600 112.300 ;
        RECT 72.255 112.440 72.545 112.485 ;
        RECT 74.145 112.440 74.435 112.485 ;
        RECT 77.265 112.440 77.555 112.485 ;
        RECT 72.255 112.300 77.555 112.440 ;
        RECT 72.255 112.255 72.545 112.300 ;
        RECT 74.145 112.255 74.435 112.300 ;
        RECT 77.265 112.255 77.555 112.300 ;
        RECT 73.210 112.100 73.530 112.160 ;
        RECT 77.900 112.100 78.040 112.640 ;
        RECT 83.345 112.595 83.635 112.640 ;
        RECT 84.710 112.580 85.030 112.840 ;
        RECT 92.545 112.780 92.835 112.825 ;
        RECT 92.545 112.640 93.220 112.780 ;
        RECT 92.545 112.595 92.835 112.640 ;
        RECT 84.215 112.440 84.505 112.485 ;
        RECT 86.105 112.440 86.395 112.485 ;
        RECT 89.225 112.440 89.515 112.485 ;
        RECT 84.215 112.300 89.515 112.440 ;
        RECT 84.215 112.255 84.505 112.300 ;
        RECT 86.105 112.255 86.395 112.300 ;
        RECT 89.225 112.255 89.515 112.300 ;
        RECT 71.460 111.960 78.040 112.100 ;
        RECT 62.170 111.900 62.490 111.960 ;
        RECT 73.210 111.900 73.530 111.960 ;
        RECT 81.030 111.900 81.350 112.160 ;
        RECT 93.080 112.100 93.220 112.640 ;
        RECT 93.910 112.580 94.230 112.840 ;
        RECT 93.415 112.440 93.705 112.485 ;
        RECT 95.305 112.440 95.595 112.485 ;
        RECT 98.425 112.440 98.715 112.485 ;
        RECT 93.415 112.300 98.715 112.440 ;
        RECT 93.415 112.255 93.705 112.300 ;
        RECT 95.305 112.255 95.595 112.300 ;
        RECT 98.425 112.255 98.715 112.300 ;
        RECT 98.970 112.440 99.290 112.500 ;
        RECT 101.285 112.440 101.575 112.485 ;
        RECT 98.970 112.300 101.575 112.440 ;
        RECT 98.970 112.240 99.290 112.300 ;
        RECT 101.285 112.255 101.575 112.300 ;
        RECT 97.590 112.100 97.910 112.160 ;
        RECT 93.080 111.960 97.910 112.100 ;
        RECT 97.590 111.900 97.910 111.960 ;
        RECT 103.585 112.100 103.875 112.145 ;
        RECT 104.030 112.100 104.350 112.160 ;
        RECT 103.585 111.960 104.350 112.100 ;
        RECT 103.585 111.915 103.875 111.960 ;
        RECT 104.030 111.900 104.350 111.960 ;
        RECT 5.520 111.280 113.620 111.760 ;
        RECT 63.550 111.080 63.870 111.140 ;
        RECT 68.165 111.080 68.455 111.125 ;
        RECT 63.550 110.940 68.455 111.080 ;
        RECT 63.550 110.880 63.870 110.940 ;
        RECT 68.165 110.895 68.455 110.940 ;
        RECT 69.070 111.080 69.390 111.140 ;
        RECT 70.925 111.080 71.215 111.125 ;
        RECT 69.070 110.940 71.215 111.080 ;
        RECT 69.070 110.880 69.390 110.940 ;
        RECT 70.925 110.895 71.215 110.940 ;
        RECT 72.750 110.880 73.070 111.140 ;
        RECT 73.670 111.080 73.990 111.140 ;
        RECT 81.490 111.080 81.810 111.140 ;
        RECT 73.300 110.940 81.810 111.080 ;
        RECT 11.225 110.740 11.515 110.785 ;
        RECT 14.345 110.740 14.635 110.785 ;
        RECT 16.235 110.740 16.525 110.785 ;
        RECT 11.225 110.600 16.525 110.740 ;
        RECT 11.225 110.555 11.515 110.600 ;
        RECT 14.345 110.555 14.635 110.600 ;
        RECT 16.235 110.555 16.525 110.600 ;
        RECT 22.725 110.740 23.015 110.785 ;
        RECT 25.845 110.740 26.135 110.785 ;
        RECT 27.735 110.740 28.025 110.785 ;
        RECT 22.725 110.600 28.025 110.740 ;
        RECT 22.725 110.555 23.015 110.600 ;
        RECT 25.845 110.555 26.135 110.600 ;
        RECT 27.735 110.555 28.025 110.600 ;
        RECT 35.455 110.740 35.745 110.785 ;
        RECT 37.345 110.740 37.635 110.785 ;
        RECT 40.465 110.740 40.755 110.785 ;
        RECT 35.455 110.600 40.755 110.740 ;
        RECT 35.455 110.555 35.745 110.600 ;
        RECT 37.345 110.555 37.635 110.600 ;
        RECT 40.465 110.555 40.755 110.600 ;
        RECT 47.875 110.740 48.165 110.785 ;
        RECT 49.765 110.740 50.055 110.785 ;
        RECT 52.885 110.740 53.175 110.785 ;
        RECT 47.875 110.600 53.175 110.740 ;
        RECT 47.875 110.555 48.165 110.600 ;
        RECT 49.765 110.555 50.055 110.600 ;
        RECT 52.885 110.555 53.175 110.600 ;
        RECT 59.835 110.740 60.125 110.785 ;
        RECT 61.725 110.740 62.015 110.785 ;
        RECT 64.845 110.740 65.135 110.785 ;
        RECT 73.300 110.740 73.440 110.940 ;
        RECT 73.670 110.880 73.990 110.940 ;
        RECT 81.490 110.880 81.810 110.940 ;
        RECT 84.265 111.080 84.555 111.125 ;
        RECT 84.710 111.080 85.030 111.140 ;
        RECT 84.265 110.940 85.030 111.080 ;
        RECT 84.265 110.895 84.555 110.940 ;
        RECT 84.710 110.880 85.030 110.940 ;
        RECT 93.910 111.080 94.230 111.140 ;
        RECT 96.225 111.080 96.515 111.125 ;
        RECT 93.910 110.940 96.515 111.080 ;
        RECT 93.910 110.880 94.230 110.940 ;
        RECT 96.225 110.895 96.515 110.940 ;
        RECT 99.430 111.080 99.750 111.140 ;
        RECT 102.650 111.080 102.970 111.140 ;
        RECT 99.430 110.940 102.970 111.080 ;
        RECT 99.430 110.880 99.750 110.940 ;
        RECT 102.650 110.880 102.970 110.940 ;
        RECT 59.835 110.600 65.135 110.740 ;
        RECT 59.835 110.555 60.125 110.600 ;
        RECT 61.725 110.555 62.015 110.600 ;
        RECT 64.845 110.555 65.135 110.600 ;
        RECT 71.460 110.600 73.440 110.740 ;
        RECT 75.015 110.740 75.305 110.785 ;
        RECT 76.905 110.740 77.195 110.785 ;
        RECT 80.025 110.740 80.315 110.785 ;
        RECT 75.015 110.600 80.315 110.740 ;
        RECT 2.830 110.400 3.150 110.460 ;
        RECT 8.365 110.400 8.655 110.445 ;
        RECT 2.830 110.260 8.655 110.400 ;
        RECT 2.830 110.200 3.150 110.260 ;
        RECT 8.365 110.215 8.655 110.260 ;
        RECT 13.410 110.400 13.730 110.460 ;
        RECT 17.105 110.400 17.395 110.445 ;
        RECT 20.770 110.400 21.090 110.460 ;
        RECT 28.605 110.400 28.895 110.445 ;
        RECT 13.410 110.260 28.895 110.400 ;
        RECT 13.410 110.200 13.730 110.260 ;
        RECT 17.105 110.215 17.395 110.260 ;
        RECT 20.770 110.200 21.090 110.260 ;
        RECT 28.605 110.215 28.895 110.260 ;
        RECT 29.510 110.200 29.830 110.460 ;
        RECT 30.060 110.260 33.420 110.400 ;
        RECT 30.060 110.105 30.200 110.260 ;
        RECT 33.280 110.120 33.420 110.260 ;
        RECT 33.650 110.200 33.970 110.460 ;
        RECT 34.585 110.400 34.875 110.445 ;
        RECT 41.930 110.400 42.250 110.460 ;
        RECT 46.990 110.400 47.310 110.460 ;
        RECT 34.585 110.260 47.310 110.400 ;
        RECT 34.585 110.215 34.875 110.260 ;
        RECT 41.930 110.200 42.250 110.260 ;
        RECT 46.990 110.200 47.310 110.260 ;
        RECT 50.670 110.400 50.990 110.460 ;
        RECT 55.745 110.400 56.035 110.445 ;
        RECT 50.670 110.260 56.035 110.400 ;
        RECT 50.670 110.200 50.990 110.260 ;
        RECT 55.745 110.215 56.035 110.260 ;
        RECT 58.965 110.400 59.255 110.445 ;
        RECT 62.170 110.400 62.490 110.460 ;
        RECT 58.965 110.260 62.490 110.400 ;
        RECT 58.965 110.215 59.255 110.260 ;
        RECT 62.170 110.200 62.490 110.260 ;
        RECT 62.630 110.400 62.950 110.460 ;
        RECT 67.705 110.400 67.995 110.445 ;
        RECT 62.630 110.260 67.995 110.400 ;
        RECT 62.630 110.200 62.950 110.260 ;
        RECT 67.705 110.215 67.995 110.260 ;
        RECT 10.145 109.765 10.435 110.080 ;
        RECT 11.225 110.060 11.515 110.105 ;
        RECT 14.805 110.060 15.095 110.105 ;
        RECT 16.640 110.060 16.930 110.105 ;
        RECT 11.225 109.920 16.930 110.060 ;
        RECT 11.225 109.875 11.515 109.920 ;
        RECT 14.805 109.875 15.095 109.920 ;
        RECT 16.640 109.875 16.930 109.920 ;
        RECT 9.845 109.720 10.435 109.765 ;
        RECT 13.085 109.720 13.735 109.765 ;
        RECT 14.330 109.720 14.650 109.780 ;
        RECT 9.845 109.580 14.650 109.720 ;
        RECT 9.845 109.535 10.135 109.580 ;
        RECT 13.085 109.535 13.735 109.580 ;
        RECT 14.330 109.520 14.650 109.580 ;
        RECT 15.710 109.520 16.030 109.780 ;
        RECT 21.645 109.765 21.935 110.080 ;
        RECT 22.725 110.060 23.015 110.105 ;
        RECT 26.305 110.060 26.595 110.105 ;
        RECT 28.140 110.060 28.430 110.105 ;
        RECT 22.725 109.920 28.430 110.060 ;
        RECT 22.725 109.875 23.015 109.920 ;
        RECT 26.305 109.875 26.595 109.920 ;
        RECT 28.140 109.875 28.430 109.920 ;
        RECT 29.985 109.875 30.275 110.105 ;
        RECT 31.825 110.060 32.115 110.105 ;
        RECT 32.730 110.060 33.050 110.120 ;
        RECT 31.825 109.920 33.050 110.060 ;
        RECT 31.825 109.875 32.115 109.920 ;
        RECT 32.730 109.860 33.050 109.920 ;
        RECT 33.190 109.860 33.510 110.120 ;
        RECT 35.050 110.060 35.340 110.105 ;
        RECT 36.885 110.060 37.175 110.105 ;
        RECT 40.465 110.060 40.755 110.105 ;
        RECT 35.050 109.920 40.755 110.060 ;
        RECT 35.050 109.875 35.340 109.920 ;
        RECT 36.885 109.875 37.175 109.920 ;
        RECT 40.465 109.875 40.755 109.920 ;
        RECT 21.345 109.720 21.935 109.765 ;
        RECT 24.585 109.720 25.235 109.765 ;
        RECT 26.750 109.720 27.070 109.780 ;
        RECT 21.345 109.580 27.070 109.720 ;
        RECT 21.345 109.535 21.635 109.580 ;
        RECT 24.585 109.535 25.235 109.580 ;
        RECT 26.750 109.520 27.070 109.580 ;
        RECT 27.210 109.520 27.530 109.780 ;
        RECT 35.950 109.520 36.270 109.780 ;
        RECT 38.245 109.720 38.895 109.765 ;
        RECT 41.010 109.720 41.330 109.780 ;
        RECT 41.545 109.765 41.835 110.080 ;
        RECT 45.150 110.060 45.470 110.120 ;
        RECT 45.625 110.060 45.915 110.105 ;
        RECT 45.150 109.920 45.915 110.060 ;
        RECT 45.150 109.860 45.470 109.920 ;
        RECT 45.625 109.875 45.915 109.920 ;
        RECT 47.470 110.060 47.760 110.105 ;
        RECT 49.305 110.060 49.595 110.105 ;
        RECT 52.885 110.060 53.175 110.105 ;
        RECT 47.470 109.920 53.175 110.060 ;
        RECT 47.470 109.875 47.760 109.920 ;
        RECT 49.305 109.875 49.595 109.920 ;
        RECT 52.885 109.875 53.175 109.920 ;
        RECT 41.545 109.720 42.135 109.765 ;
        RECT 48.385 109.720 48.675 109.765 ;
        RECT 38.245 109.580 42.135 109.720 ;
        RECT 38.245 109.535 38.895 109.580 ;
        RECT 41.010 109.520 41.330 109.580 ;
        RECT 41.845 109.535 42.135 109.580 ;
        RECT 46.620 109.580 48.675 109.720 ;
        RECT 19.865 109.380 20.155 109.425 ;
        RECT 20.770 109.380 21.090 109.440 ;
        RECT 19.865 109.240 21.090 109.380 ;
        RECT 19.865 109.195 20.155 109.240 ;
        RECT 20.770 109.180 21.090 109.240 ;
        RECT 32.745 109.380 33.035 109.425 ;
        RECT 35.490 109.380 35.810 109.440 ;
        RECT 32.745 109.240 35.810 109.380 ;
        RECT 32.745 109.195 33.035 109.240 ;
        RECT 35.490 109.180 35.810 109.240 ;
        RECT 39.170 109.380 39.490 109.440 ;
        RECT 46.620 109.425 46.760 109.580 ;
        RECT 48.385 109.535 48.675 109.580 ;
        RECT 50.665 109.720 51.315 109.765 ;
        RECT 51.590 109.720 51.910 109.780 ;
        RECT 53.965 109.765 54.255 110.080 ;
        RECT 56.205 110.060 56.495 110.105 ;
        RECT 57.110 110.060 57.430 110.120 ;
        RECT 56.205 109.920 57.430 110.060 ;
        RECT 56.205 109.875 56.495 109.920 ;
        RECT 57.110 109.860 57.430 109.920 ;
        RECT 59.430 110.060 59.720 110.105 ;
        RECT 61.265 110.060 61.555 110.105 ;
        RECT 64.845 110.060 65.135 110.105 ;
        RECT 59.430 109.920 65.135 110.060 ;
        RECT 59.430 109.875 59.720 109.920 ;
        RECT 61.265 109.875 61.555 109.920 ;
        RECT 64.845 109.875 65.135 109.920 ;
        RECT 65.850 110.080 66.170 110.120 ;
        RECT 65.850 109.860 66.215 110.080 ;
        RECT 69.070 109.860 69.390 110.120 ;
        RECT 69.530 110.060 69.850 110.120 ;
        RECT 71.460 110.105 71.600 110.600 ;
        RECT 75.015 110.555 75.305 110.600 ;
        RECT 76.905 110.555 77.195 110.600 ;
        RECT 80.025 110.555 80.315 110.600 ;
        RECT 86.515 110.740 86.805 110.785 ;
        RECT 88.405 110.740 88.695 110.785 ;
        RECT 91.525 110.740 91.815 110.785 ;
        RECT 86.515 110.600 91.815 110.740 ;
        RECT 86.515 110.555 86.805 110.600 ;
        RECT 88.405 110.555 88.695 110.600 ;
        RECT 91.525 110.555 91.815 110.600 ;
        RECT 98.475 110.740 98.765 110.785 ;
        RECT 100.365 110.740 100.655 110.785 ;
        RECT 103.485 110.740 103.775 110.785 ;
        RECT 98.475 110.600 103.775 110.740 ;
        RECT 98.475 110.555 98.765 110.600 ;
        RECT 100.365 110.555 100.655 110.600 ;
        RECT 103.485 110.555 103.775 110.600 ;
        RECT 73.210 110.400 73.530 110.460 ;
        RECT 74.145 110.400 74.435 110.445 ;
        RECT 73.210 110.260 74.435 110.400 ;
        RECT 73.210 110.200 73.530 110.260 ;
        RECT 74.145 110.215 74.435 110.260 ;
        RECT 80.570 110.400 80.890 110.460 ;
        RECT 82.885 110.400 83.175 110.445 ;
        RECT 97.590 110.400 97.910 110.460 ;
        RECT 80.570 110.260 83.175 110.400 ;
        RECT 80.570 110.200 80.890 110.260 ;
        RECT 82.885 110.215 83.175 110.260 ;
        RECT 85.720 110.260 97.910 110.400 ;
        RECT 71.385 110.060 71.675 110.105 ;
        RECT 69.530 109.920 71.675 110.060 ;
        RECT 69.530 109.860 69.850 109.920 ;
        RECT 71.385 109.875 71.675 109.920 ;
        RECT 73.685 109.875 73.975 110.105 ;
        RECT 74.610 110.060 74.900 110.105 ;
        RECT 76.445 110.060 76.735 110.105 ;
        RECT 80.025 110.060 80.315 110.105 ;
        RECT 74.610 109.920 80.315 110.060 ;
        RECT 74.610 109.875 74.900 109.920 ;
        RECT 76.445 109.875 76.735 109.920 ;
        RECT 80.025 109.875 80.315 109.920 ;
        RECT 81.030 110.080 81.350 110.120 ;
        RECT 65.925 109.765 66.215 109.860 ;
        RECT 53.965 109.720 54.555 109.765 ;
        RECT 50.665 109.580 54.555 109.720 ;
        RECT 50.665 109.535 51.315 109.580 ;
        RECT 51.590 109.520 51.910 109.580 ;
        RECT 54.265 109.535 54.555 109.580 ;
        RECT 60.345 109.720 60.635 109.765 ;
        RECT 62.625 109.720 63.275 109.765 ;
        RECT 65.925 109.720 66.515 109.765 ;
        RECT 60.345 109.580 62.400 109.720 ;
        RECT 60.345 109.535 60.635 109.580 ;
        RECT 62.260 109.440 62.400 109.580 ;
        RECT 62.625 109.580 66.515 109.720 ;
        RECT 62.625 109.535 63.275 109.580 ;
        RECT 66.225 109.535 66.515 109.580 ;
        RECT 43.325 109.380 43.615 109.425 ;
        RECT 39.170 109.240 43.615 109.380 ;
        RECT 39.170 109.180 39.490 109.240 ;
        RECT 43.325 109.195 43.615 109.240 ;
        RECT 46.545 109.195 46.835 109.425 ;
        RECT 56.665 109.380 56.955 109.425 ;
        RECT 61.710 109.380 62.030 109.440 ;
        RECT 56.665 109.240 62.030 109.380 ;
        RECT 56.665 109.195 56.955 109.240 ;
        RECT 61.710 109.180 62.030 109.240 ;
        RECT 62.170 109.180 62.490 109.440 ;
        RECT 73.760 109.380 73.900 109.875 ;
        RECT 81.030 109.860 81.395 110.080 ;
        RECT 83.330 109.860 83.650 110.120 ;
        RECT 85.720 110.105 85.860 110.260 ;
        RECT 97.590 110.200 97.910 110.260 ;
        RECT 105.870 110.400 106.190 110.460 ;
        RECT 106.345 110.400 106.635 110.445 ;
        RECT 105.870 110.260 106.635 110.400 ;
        RECT 105.870 110.200 106.190 110.260 ;
        RECT 106.345 110.215 106.635 110.260 ;
        RECT 85.645 109.875 85.935 110.105 ;
        RECT 86.110 110.060 86.400 110.105 ;
        RECT 87.945 110.060 88.235 110.105 ;
        RECT 91.525 110.060 91.815 110.105 ;
        RECT 86.110 109.920 91.815 110.060 ;
        RECT 86.110 109.875 86.400 109.920 ;
        RECT 87.945 109.875 88.235 109.920 ;
        RECT 91.525 109.875 91.815 109.920 ;
        RECT 75.525 109.720 75.815 109.765 ;
        RECT 76.890 109.720 77.210 109.780 ;
        RECT 81.105 109.765 81.395 109.860 ;
        RECT 75.525 109.580 77.210 109.720 ;
        RECT 75.525 109.535 75.815 109.580 ;
        RECT 76.890 109.520 77.210 109.580 ;
        RECT 77.805 109.720 78.455 109.765 ;
        RECT 81.105 109.720 81.695 109.765 ;
        RECT 77.805 109.580 81.695 109.720 ;
        RECT 85.720 109.720 85.860 109.875 ;
        RECT 86.550 109.720 86.870 109.780 ;
        RECT 85.720 109.580 86.870 109.720 ;
        RECT 77.805 109.535 78.455 109.580 ;
        RECT 81.405 109.535 81.695 109.580 ;
        RECT 86.550 109.520 86.870 109.580 ;
        RECT 87.010 109.520 87.330 109.780 ;
        RECT 89.305 109.720 89.955 109.765 ;
        RECT 90.690 109.720 91.010 109.780 ;
        RECT 92.605 109.765 92.895 110.080 ;
        RECT 97.145 109.875 97.435 110.105 ;
        RECT 98.070 110.060 98.360 110.105 ;
        RECT 99.905 110.060 100.195 110.105 ;
        RECT 103.485 110.060 103.775 110.105 ;
        RECT 98.070 109.920 103.775 110.060 ;
        RECT 98.070 109.875 98.360 109.920 ;
        RECT 99.905 109.875 100.195 109.920 ;
        RECT 103.485 109.875 103.775 109.920 ;
        RECT 92.605 109.720 93.195 109.765 ;
        RECT 89.305 109.580 93.195 109.720 ;
        RECT 89.305 109.535 89.955 109.580 ;
        RECT 90.690 109.520 91.010 109.580 ;
        RECT 92.905 109.535 93.195 109.580 ;
        RECT 77.350 109.380 77.670 109.440 ;
        RECT 73.760 109.240 77.670 109.380 ;
        RECT 77.350 109.180 77.670 109.240 ;
        RECT 92.070 109.380 92.390 109.440 ;
        RECT 94.385 109.380 94.675 109.425 ;
        RECT 92.070 109.240 94.675 109.380 ;
        RECT 97.220 109.380 97.360 109.875 ;
        RECT 98.970 109.520 99.290 109.780 ;
        RECT 101.265 109.720 101.915 109.765 ;
        RECT 104.030 109.720 104.350 109.780 ;
        RECT 104.565 109.765 104.855 110.080 ;
        RECT 104.565 109.720 105.155 109.765 ;
        RECT 101.265 109.580 105.155 109.720 ;
        RECT 101.265 109.535 101.915 109.580 ;
        RECT 104.030 109.520 104.350 109.580 ;
        RECT 104.865 109.535 105.155 109.580 ;
        RECT 98.050 109.380 98.370 109.440 ;
        RECT 97.220 109.240 98.370 109.380 ;
        RECT 92.070 109.180 92.390 109.240 ;
        RECT 94.385 109.195 94.675 109.240 ;
        RECT 98.050 109.180 98.370 109.240 ;
        RECT 5.520 108.560 113.620 109.040 ;
        RECT 8.810 108.360 9.130 108.420 ;
        RECT 15.725 108.360 16.015 108.405 ;
        RECT 8.810 108.220 16.015 108.360 ;
        RECT 8.810 108.160 9.130 108.220 ;
        RECT 15.725 108.175 16.015 108.220 ;
        RECT 18.010 108.160 18.330 108.420 ;
        RECT 22.610 108.360 22.930 108.420 ;
        RECT 24.465 108.360 24.755 108.405 ;
        RECT 22.610 108.220 24.755 108.360 ;
        RECT 22.610 108.160 22.930 108.220 ;
        RECT 24.465 108.175 24.755 108.220 ;
        RECT 26.305 108.360 26.595 108.405 ;
        RECT 26.750 108.360 27.070 108.420 ;
        RECT 26.305 108.220 27.070 108.360 ;
        RECT 26.305 108.175 26.595 108.220 ;
        RECT 26.750 108.160 27.070 108.220 ;
        RECT 35.950 108.360 36.270 108.420 ;
        RECT 39.185 108.360 39.475 108.405 ;
        RECT 35.950 108.220 39.475 108.360 ;
        RECT 35.950 108.160 36.270 108.220 ;
        RECT 39.185 108.175 39.475 108.220 ;
        RECT 41.010 108.160 41.330 108.420 ;
        RECT 42.390 108.160 42.710 108.420 ;
        RECT 44.245 108.360 44.535 108.405 ;
        RECT 44.690 108.360 45.010 108.420 ;
        RECT 44.245 108.220 45.010 108.360 ;
        RECT 44.245 108.175 44.535 108.220 ;
        RECT 44.690 108.160 45.010 108.220 ;
        RECT 49.290 108.360 49.610 108.420 ;
        RECT 52.525 108.360 52.815 108.405 ;
        RECT 49.290 108.220 52.815 108.360 ;
        RECT 49.290 108.160 49.610 108.220 ;
        RECT 52.525 108.175 52.815 108.220 ;
        RECT 62.170 108.360 62.490 108.420 ;
        RECT 62.645 108.360 62.935 108.405 ;
        RECT 62.170 108.220 62.935 108.360 ;
        RECT 62.170 108.160 62.490 108.220 ;
        RECT 62.645 108.175 62.935 108.220 ;
        RECT 65.850 108.360 66.170 108.420 ;
        RECT 66.325 108.360 66.615 108.405 ;
        RECT 65.850 108.220 66.615 108.360 ;
        RECT 65.850 108.160 66.170 108.220 ;
        RECT 66.325 108.175 66.615 108.220 ;
        RECT 73.685 108.360 73.975 108.405 ;
        RECT 75.970 108.360 76.290 108.420 ;
        RECT 73.685 108.220 76.290 108.360 ;
        RECT 73.685 108.175 73.975 108.220 ;
        RECT 75.970 108.160 76.290 108.220 ;
        RECT 76.890 108.360 77.210 108.420 ;
        RECT 78.285 108.360 78.575 108.405 ;
        RECT 76.890 108.220 78.575 108.360 ;
        RECT 76.890 108.160 77.210 108.220 ;
        RECT 78.285 108.175 78.575 108.220 ;
        RECT 87.010 108.160 87.330 108.420 ;
        RECT 97.145 108.360 97.435 108.405 ;
        RECT 98.970 108.360 99.290 108.420 ;
        RECT 97.145 108.220 99.290 108.360 ;
        RECT 97.145 108.175 97.435 108.220 ;
        RECT 98.970 108.160 99.290 108.220 ;
        RECT 107.265 108.360 107.555 108.405 ;
        RECT 110.470 108.360 110.790 108.420 ;
        RECT 107.265 108.220 110.790 108.360 ;
        RECT 107.265 108.175 107.555 108.220 ;
        RECT 110.470 108.160 110.790 108.220 ;
        RECT 10.645 108.020 11.295 108.065 ;
        RECT 14.245 108.020 14.535 108.065 ;
        RECT 16.645 108.020 16.935 108.065 ;
        RECT 33.190 108.020 33.510 108.080 ;
        RECT 50.685 108.020 50.975 108.065 ;
        RECT 51.130 108.020 51.450 108.080 ;
        RECT 68.150 108.020 68.470 108.080 ;
        RECT 10.645 107.880 16.935 108.020 ;
        RECT 10.645 107.835 11.295 107.880 ;
        RECT 13.945 107.835 14.535 107.880 ;
        RECT 16.645 107.835 16.935 107.880 ;
        RECT 18.560 107.880 26.980 108.020 ;
        RECT 7.450 107.680 7.740 107.725 ;
        RECT 9.285 107.680 9.575 107.725 ;
        RECT 12.865 107.680 13.155 107.725 ;
        RECT 7.450 107.540 13.155 107.680 ;
        RECT 7.450 107.495 7.740 107.540 ;
        RECT 9.285 107.495 9.575 107.540 ;
        RECT 12.865 107.495 13.155 107.540 ;
        RECT 13.945 107.520 14.235 107.835 ;
        RECT 15.250 107.680 15.570 107.740 ;
        RECT 18.560 107.725 18.700 107.880 ;
        RECT 17.105 107.680 17.395 107.725 ;
        RECT 18.485 107.680 18.775 107.725 ;
        RECT 15.250 107.540 18.775 107.680 ;
        RECT 15.250 107.480 15.570 107.540 ;
        RECT 17.105 107.495 17.395 107.540 ;
        RECT 18.485 107.495 18.775 107.540 ;
        RECT 20.785 107.495 21.075 107.725 ;
        RECT 6.970 107.140 7.290 107.400 ;
        RECT 8.350 107.140 8.670 107.400 ;
        RECT 7.855 107.000 8.145 107.045 ;
        RECT 9.745 107.000 10.035 107.045 ;
        RECT 12.865 107.000 13.155 107.045 ;
        RECT 7.855 106.860 13.155 107.000 ;
        RECT 7.855 106.815 8.145 106.860 ;
        RECT 9.745 106.815 10.035 106.860 ;
        RECT 12.865 106.815 13.155 106.860 ;
        RECT 17.550 107.000 17.870 107.060 ;
        RECT 19.865 107.000 20.155 107.045 ;
        RECT 17.550 106.860 20.155 107.000 ;
        RECT 17.550 106.800 17.870 106.860 ;
        RECT 19.865 106.815 20.155 106.860 ;
        RECT 20.860 106.660 21.000 107.495 ;
        RECT 23.530 107.480 23.850 107.740 ;
        RECT 26.840 107.725 26.980 107.880 ;
        RECT 33.190 107.880 44.920 108.020 ;
        RECT 33.190 107.820 33.510 107.880 ;
        RECT 25.385 107.495 25.675 107.725 ;
        RECT 26.765 107.680 27.055 107.725 ;
        RECT 33.280 107.680 33.420 107.820 ;
        RECT 41.560 107.725 41.700 107.880 ;
        RECT 44.780 107.725 44.920 107.880 ;
        RECT 50.685 107.880 51.450 108.020 ;
        RECT 50.685 107.835 50.975 107.880 ;
        RECT 26.765 107.540 33.420 107.680 ;
        RECT 26.765 107.495 27.055 107.540 ;
        RECT 40.105 107.495 40.395 107.725 ;
        RECT 41.485 107.495 41.775 107.725 ;
        RECT 43.325 107.495 43.615 107.725 ;
        RECT 44.705 107.680 44.995 107.725 ;
        RECT 50.760 107.680 50.900 107.835 ;
        RECT 51.130 107.820 51.450 107.880 ;
        RECT 63.640 107.880 68.470 108.020 ;
        RECT 44.705 107.540 50.900 107.680 ;
        RECT 44.705 107.495 44.995 107.540 ;
        RECT 52.065 107.495 52.355 107.725 ;
        RECT 52.970 107.680 53.290 107.740 ;
        RECT 63.640 107.725 63.780 107.880 ;
        RECT 68.150 107.820 68.470 107.880 ;
        RECT 69.070 108.020 69.390 108.080 ;
        RECT 76.430 108.020 76.750 108.080 ;
        RECT 69.070 107.880 76.750 108.020 ;
        RECT 69.070 107.820 69.390 107.880 ;
        RECT 76.430 107.820 76.750 107.880 ;
        RECT 102.185 108.020 102.835 108.065 ;
        RECT 104.950 108.020 105.270 108.080 ;
        RECT 105.785 108.020 106.075 108.065 ;
        RECT 102.185 107.880 106.075 108.020 ;
        RECT 102.185 107.835 102.835 107.880 ;
        RECT 104.950 107.820 105.270 107.880 ;
        RECT 105.485 107.835 106.075 107.880 ;
        RECT 53.445 107.680 53.735 107.725 ;
        RECT 52.970 107.540 53.735 107.680 ;
        RECT 21.690 107.340 22.010 107.400 ;
        RECT 25.460 107.340 25.600 107.495 ;
        RECT 21.690 107.200 25.600 107.340 ;
        RECT 21.690 107.140 22.010 107.200 ;
        RECT 22.625 107.000 22.915 107.045 ;
        RECT 27.210 107.000 27.530 107.060 ;
        RECT 22.625 106.860 27.530 107.000 ;
        RECT 22.625 106.815 22.915 106.860 ;
        RECT 27.210 106.800 27.530 106.860 ;
        RECT 29.510 106.660 29.830 106.720 ;
        RECT 20.860 106.520 29.830 106.660 ;
        RECT 40.180 106.660 40.320 107.495 ;
        RECT 43.400 107.000 43.540 107.495 ;
        RECT 52.140 107.340 52.280 107.495 ;
        RECT 52.970 107.480 53.290 107.540 ;
        RECT 53.445 107.495 53.735 107.540 ;
        RECT 63.565 107.495 63.855 107.725 ;
        RECT 66.785 107.680 67.075 107.725 ;
        RECT 69.530 107.680 69.850 107.740 ;
        RECT 66.785 107.540 69.850 107.680 ;
        RECT 66.785 107.495 67.075 107.540 ;
        RECT 69.530 107.480 69.850 107.540 ;
        RECT 70.925 107.495 71.215 107.725 ;
        RECT 73.225 107.680 73.515 107.725 ;
        RECT 73.670 107.680 73.990 107.740 ;
        RECT 73.225 107.540 73.990 107.680 ;
        RECT 73.225 107.495 73.515 107.540 ;
        RECT 64.470 107.340 64.790 107.400 ;
        RECT 71.000 107.340 71.140 107.495 ;
        RECT 73.670 107.480 73.990 107.540 ;
        RECT 79.190 107.480 79.510 107.740 ;
        RECT 87.930 107.480 88.250 107.740 ;
        RECT 95.750 107.680 96.070 107.740 ;
        RECT 96.225 107.680 96.515 107.725 ;
        RECT 95.750 107.540 96.515 107.680 ;
        RECT 95.750 107.480 96.070 107.540 ;
        RECT 96.225 107.495 96.515 107.540 ;
        RECT 97.590 107.680 97.910 107.740 ;
        RECT 98.525 107.680 98.815 107.725 ;
        RECT 97.590 107.540 98.815 107.680 ;
        RECT 97.590 107.480 97.910 107.540 ;
        RECT 98.525 107.495 98.815 107.540 ;
        RECT 98.990 107.680 99.280 107.725 ;
        RECT 100.825 107.680 101.115 107.725 ;
        RECT 104.405 107.680 104.695 107.725 ;
        RECT 98.990 107.540 104.695 107.680 ;
        RECT 98.990 107.495 99.280 107.540 ;
        RECT 100.825 107.495 101.115 107.540 ;
        RECT 104.405 107.495 104.695 107.540 ;
        RECT 105.485 107.520 105.775 107.835 ;
        RECT 99.905 107.340 100.195 107.385 ;
        RECT 52.140 107.200 71.140 107.340 ;
        RECT 98.600 107.200 100.195 107.340 ;
        RECT 64.470 107.140 64.790 107.200 ;
        RECT 98.600 107.060 98.740 107.200 ;
        RECT 99.905 107.155 100.195 107.200 ;
        RECT 57.110 107.000 57.430 107.060 ;
        RECT 43.400 106.860 57.430 107.000 ;
        RECT 57.110 106.800 57.430 106.860 ;
        RECT 98.510 106.800 98.830 107.060 ;
        RECT 99.395 107.000 99.685 107.045 ;
        RECT 101.285 107.000 101.575 107.045 ;
        RECT 104.405 107.000 104.695 107.045 ;
        RECT 99.395 106.860 104.695 107.000 ;
        RECT 99.395 106.815 99.685 106.860 ;
        RECT 101.285 106.815 101.575 106.860 ;
        RECT 104.405 106.815 104.695 106.860 ;
        RECT 48.830 106.660 49.150 106.720 ;
        RECT 40.180 106.520 49.150 106.660 ;
        RECT 29.510 106.460 29.830 106.520 ;
        RECT 48.830 106.460 49.150 106.520 ;
        RECT 5.520 105.840 113.620 106.320 ;
        RECT 8.350 105.640 8.670 105.700 ;
        RECT 9.745 105.640 10.035 105.685 ;
        RECT 8.350 105.500 10.035 105.640 ;
        RECT 8.350 105.440 8.670 105.500 ;
        RECT 9.745 105.455 10.035 105.500 ;
        RECT 12.045 105.640 12.335 105.685 ;
        RECT 15.710 105.640 16.030 105.700 ;
        RECT 12.045 105.500 16.030 105.640 ;
        RECT 12.045 105.455 12.335 105.500 ;
        RECT 15.710 105.440 16.030 105.500 ;
        RECT 98.510 105.440 98.830 105.700 ;
        RECT 104.505 105.640 104.795 105.685 ;
        RECT 104.950 105.640 105.270 105.700 ;
        RECT 104.505 105.500 105.270 105.640 ;
        RECT 104.505 105.455 104.795 105.500 ;
        RECT 104.950 105.440 105.270 105.500 ;
        RECT 14.330 105.300 14.650 105.360 ;
        RECT 14.805 105.300 15.095 105.345 ;
        RECT 14.330 105.160 15.095 105.300 ;
        RECT 14.330 105.100 14.650 105.160 ;
        RECT 14.805 105.115 15.095 105.160 ;
        RECT 30.430 104.960 30.750 105.020 ;
        RECT 13.040 104.820 30.750 104.960 ;
        RECT 13.040 104.665 13.180 104.820 ;
        RECT 30.430 104.760 30.750 104.820 ;
        RECT 47.910 104.960 48.230 105.020 ;
        RECT 48.845 104.960 49.135 105.005 ;
        RECT 47.910 104.820 49.135 104.960 ;
        RECT 47.910 104.760 48.230 104.820 ;
        RECT 48.845 104.775 49.135 104.820 ;
        RECT 69.530 104.960 69.850 105.020 ;
        RECT 73.225 104.960 73.515 105.005 ;
        RECT 69.530 104.820 73.515 104.960 ;
        RECT 69.530 104.760 69.850 104.820 ;
        RECT 73.225 104.775 73.515 104.820 ;
        RECT 10.665 104.435 10.955 104.665 ;
        RECT 12.965 104.435 13.255 104.665 ;
        RECT 10.740 104.280 10.880 104.435 ;
        RECT 15.250 104.420 15.570 104.680 ;
        RECT 36.425 104.620 36.715 104.665 ;
        RECT 42.850 104.620 43.170 104.680 ;
        RECT 36.425 104.480 43.170 104.620 ;
        RECT 36.425 104.435 36.715 104.480 ;
        RECT 42.850 104.420 43.170 104.480 ;
        RECT 64.470 104.620 64.790 104.680 ;
        RECT 75.510 104.620 75.830 104.680 ;
        RECT 64.470 104.480 75.830 104.620 ;
        RECT 64.470 104.420 64.790 104.480 ;
        RECT 75.510 104.420 75.830 104.480 ;
        RECT 97.130 104.420 97.450 104.680 ;
        RECT 97.590 104.420 97.910 104.680 ;
        RECT 104.490 104.620 104.810 104.680 ;
        RECT 104.965 104.620 105.255 104.665 ;
        RECT 104.490 104.480 105.255 104.620 ;
        RECT 104.490 104.420 104.810 104.480 ;
        RECT 104.965 104.435 105.255 104.480 ;
        RECT 18.010 104.280 18.330 104.340 ;
        RECT 10.740 104.140 18.330 104.280 ;
        RECT 18.010 104.080 18.330 104.140 ;
        RECT 47.925 104.280 48.215 104.325 ;
        RECT 51.590 104.280 51.910 104.340 ;
        RECT 47.925 104.140 51.910 104.280 ;
        RECT 47.925 104.095 48.215 104.140 ;
        RECT 51.590 104.080 51.910 104.140 ;
        RECT 35.490 103.940 35.810 104.000 ;
        RECT 35.965 103.940 36.255 103.985 ;
        RECT 35.490 103.800 36.255 103.940 ;
        RECT 35.490 103.740 35.810 103.800 ;
        RECT 35.965 103.755 36.255 103.800 ;
        RECT 46.085 103.940 46.375 103.985 ;
        RECT 46.530 103.940 46.850 104.000 ;
        RECT 46.085 103.800 46.850 103.940 ;
        RECT 46.085 103.755 46.375 103.800 ;
        RECT 46.530 103.740 46.850 103.800 ;
        RECT 47.450 103.940 47.770 104.000 ;
        RECT 48.385 103.940 48.675 103.985 ;
        RECT 47.450 103.800 48.675 103.940 ;
        RECT 47.450 103.740 47.770 103.800 ;
        RECT 48.385 103.755 48.675 103.800 ;
        RECT 69.070 103.940 69.390 104.000 ;
        RECT 70.465 103.940 70.755 103.985 ;
        RECT 69.070 103.800 70.755 103.940 ;
        RECT 69.070 103.740 69.390 103.800 ;
        RECT 70.465 103.755 70.755 103.800 ;
        RECT 72.290 103.740 72.610 104.000 ;
        RECT 72.765 103.940 73.055 103.985 ;
        RECT 73.670 103.940 73.990 104.000 ;
        RECT 72.765 103.800 73.990 103.940 ;
        RECT 72.765 103.755 73.055 103.800 ;
        RECT 73.670 103.740 73.990 103.800 ;
        RECT 75.050 103.740 75.370 104.000 ;
        RECT 96.670 103.740 96.990 104.000 ;
        RECT 5.520 103.120 113.620 103.600 ;
        RECT 63.565 102.920 63.855 102.965 ;
        RECT 73.670 102.920 73.990 102.980 ;
        RECT 97.130 102.920 97.450 102.980 ;
        RECT 63.565 102.780 73.990 102.920 ;
        RECT 63.565 102.735 63.855 102.780 ;
        RECT 73.670 102.720 73.990 102.780 ;
        RECT 81.580 102.780 97.450 102.920 ;
        RECT 23.070 102.625 23.390 102.640 ;
        RECT 17.110 102.580 17.400 102.625 ;
        RECT 18.970 102.580 19.260 102.625 ;
        RECT 17.110 102.440 19.260 102.580 ;
        RECT 17.110 102.395 17.400 102.440 ;
        RECT 18.970 102.395 19.260 102.440 ;
        RECT 19.890 102.580 20.180 102.625 ;
        RECT 23.070 102.580 23.440 102.625 ;
        RECT 19.890 102.440 23.440 102.580 ;
        RECT 19.890 102.395 20.180 102.440 ;
        RECT 23.070 102.395 23.440 102.440 ;
        RECT 34.060 102.580 34.350 102.625 ;
        RECT 35.490 102.580 35.810 102.640 ;
        RECT 37.320 102.580 37.610 102.625 ;
        RECT 34.060 102.440 37.610 102.580 ;
        RECT 34.060 102.395 34.350 102.440 ;
        RECT 19.045 102.240 19.260 102.395 ;
        RECT 23.070 102.380 23.390 102.395 ;
        RECT 35.490 102.380 35.810 102.440 ;
        RECT 37.320 102.395 37.610 102.440 ;
        RECT 38.240 102.580 38.530 102.625 ;
        RECT 40.100 102.580 40.390 102.625 ;
        RECT 38.240 102.440 40.390 102.580 ;
        RECT 38.240 102.395 38.530 102.440 ;
        RECT 40.100 102.395 40.390 102.440 ;
        RECT 44.710 102.580 45.000 102.625 ;
        RECT 46.570 102.580 46.860 102.625 ;
        RECT 44.710 102.440 46.860 102.580 ;
        RECT 44.710 102.395 45.000 102.440 ;
        RECT 46.570 102.395 46.860 102.440 ;
        RECT 47.490 102.580 47.780 102.625 ;
        RECT 49.290 102.580 49.610 102.640 ;
        RECT 50.750 102.580 51.040 102.625 ;
        RECT 47.490 102.440 51.040 102.580 ;
        RECT 47.490 102.395 47.780 102.440 ;
        RECT 21.290 102.240 21.580 102.285 ;
        RECT 19.045 102.100 21.580 102.240 ;
        RECT 21.290 102.055 21.580 102.100 ;
        RECT 26.750 102.240 27.070 102.300 ;
        RECT 27.685 102.240 27.975 102.285 ;
        RECT 26.750 102.100 27.975 102.240 ;
        RECT 26.750 102.040 27.070 102.100 ;
        RECT 27.685 102.055 27.975 102.100 ;
        RECT 35.920 102.240 36.210 102.285 ;
        RECT 38.240 102.240 38.455 102.395 ;
        RECT 35.920 102.100 38.455 102.240 ;
        RECT 42.405 102.240 42.695 102.285 ;
        RECT 42.850 102.240 43.170 102.300 ;
        RECT 42.405 102.100 43.170 102.240 ;
        RECT 46.645 102.240 46.860 102.395 ;
        RECT 49.290 102.380 49.610 102.440 ;
        RECT 50.750 102.395 51.040 102.440 ;
        RECT 66.790 102.580 67.080 102.625 ;
        RECT 68.650 102.580 68.940 102.625 ;
        RECT 66.790 102.440 68.940 102.580 ;
        RECT 66.790 102.395 67.080 102.440 ;
        RECT 68.650 102.395 68.940 102.440 ;
        RECT 69.570 102.580 69.860 102.625 ;
        RECT 72.830 102.580 73.120 102.625 ;
        RECT 75.050 102.580 75.370 102.640 ;
        RECT 69.570 102.440 75.370 102.580 ;
        RECT 69.570 102.395 69.860 102.440 ;
        RECT 72.830 102.395 73.120 102.440 ;
        RECT 48.890 102.240 49.180 102.285 ;
        RECT 46.645 102.100 49.180 102.240 ;
        RECT 35.920 102.055 36.210 102.100 ;
        RECT 42.405 102.055 42.695 102.100 ;
        RECT 42.850 102.040 43.170 102.100 ;
        RECT 48.890 102.055 49.180 102.100 ;
        RECT 53.445 102.240 53.735 102.285 ;
        RECT 53.890 102.240 54.210 102.300 ;
        RECT 53.445 102.100 54.210 102.240 ;
        RECT 53.445 102.055 53.735 102.100 ;
        RECT 53.890 102.040 54.210 102.100 ;
        RECT 60.345 102.240 60.635 102.285 ;
        RECT 64.470 102.240 64.790 102.300 ;
        RECT 60.345 102.100 64.790 102.240 ;
        RECT 60.345 102.055 60.635 102.100 ;
        RECT 64.470 102.040 64.790 102.100 ;
        RECT 65.865 102.240 66.155 102.285 ;
        RECT 68.725 102.240 68.940 102.395 ;
        RECT 75.050 102.380 75.370 102.440 ;
        RECT 76.905 102.580 77.195 102.625 ;
        RECT 81.580 102.580 81.720 102.780 ;
        RECT 97.130 102.720 97.450 102.780 ;
        RECT 76.905 102.440 81.720 102.580 ;
        RECT 76.905 102.395 77.195 102.440 ;
        RECT 70.970 102.240 71.260 102.285 ;
        RECT 65.865 102.100 68.380 102.240 ;
        RECT 68.725 102.100 71.260 102.240 ;
        RECT 65.865 102.055 66.155 102.100 ;
        RECT 13.410 101.900 13.730 101.960 ;
        RECT 16.185 101.900 16.475 101.945 ;
        RECT 13.410 101.760 16.475 101.900 ;
        RECT 13.410 101.700 13.730 101.760 ;
        RECT 16.185 101.715 16.475 101.760 ;
        RECT 17.550 101.900 17.870 101.960 ;
        RECT 18.025 101.900 18.315 101.945 ;
        RECT 39.185 101.900 39.475 101.945 ;
        RECT 17.550 101.760 18.315 101.900 ;
        RECT 17.550 101.700 17.870 101.760 ;
        RECT 18.025 101.715 18.315 101.760 ;
        RECT 28.680 101.760 39.475 101.900 ;
        RECT 28.680 101.605 28.820 101.760 ;
        RECT 39.185 101.715 39.475 101.760 ;
        RECT 41.025 101.900 41.315 101.945 ;
        RECT 41.930 101.900 42.250 101.960 ;
        RECT 43.785 101.900 44.075 101.945 ;
        RECT 41.025 101.760 44.075 101.900 ;
        RECT 41.025 101.715 41.315 101.760 ;
        RECT 41.930 101.700 42.250 101.760 ;
        RECT 43.785 101.715 44.075 101.760 ;
        RECT 45.610 101.700 45.930 101.960 ;
        RECT 62.630 101.900 62.950 101.960 ;
        RECT 64.025 101.900 64.315 101.945 ;
        RECT 62.630 101.760 64.315 101.900 ;
        RECT 62.630 101.700 62.950 101.760 ;
        RECT 64.025 101.715 64.315 101.760 ;
        RECT 64.945 101.900 65.235 101.945 ;
        RECT 64.945 101.760 66.080 101.900 ;
        RECT 64.945 101.715 65.235 101.760 ;
        RECT 16.650 101.560 16.940 101.605 ;
        RECT 18.510 101.560 18.800 101.605 ;
        RECT 21.290 101.560 21.580 101.605 ;
        RECT 16.650 101.420 21.580 101.560 ;
        RECT 16.650 101.375 16.940 101.420 ;
        RECT 18.510 101.375 18.800 101.420 ;
        RECT 21.290 101.375 21.580 101.420 ;
        RECT 28.605 101.375 28.895 101.605 ;
        RECT 35.920 101.560 36.210 101.605 ;
        RECT 38.700 101.560 38.990 101.605 ;
        RECT 40.560 101.560 40.850 101.605 ;
        RECT 35.920 101.420 40.850 101.560 ;
        RECT 35.920 101.375 36.210 101.420 ;
        RECT 38.700 101.375 38.990 101.420 ;
        RECT 40.560 101.375 40.850 101.420 ;
        RECT 44.250 101.560 44.540 101.605 ;
        RECT 46.110 101.560 46.400 101.605 ;
        RECT 48.890 101.560 49.180 101.605 ;
        RECT 44.250 101.420 49.180 101.560 ;
        RECT 44.250 101.375 44.540 101.420 ;
        RECT 46.110 101.375 46.400 101.420 ;
        RECT 48.890 101.375 49.180 101.420 ;
        RECT 22.610 101.220 22.930 101.280 ;
        RECT 25.155 101.220 25.445 101.265 ;
        RECT 22.610 101.080 25.445 101.220 ;
        RECT 22.610 101.020 22.930 101.080 ;
        RECT 25.155 101.035 25.445 101.080 ;
        RECT 29.970 101.220 30.290 101.280 ;
        RECT 32.055 101.220 32.345 101.265 ;
        RECT 33.650 101.220 33.970 101.280 ;
        RECT 29.970 101.080 33.970 101.220 ;
        RECT 29.970 101.020 30.290 101.080 ;
        RECT 32.055 101.035 32.345 101.080 ;
        RECT 33.650 101.020 33.970 101.080 ;
        RECT 39.170 101.220 39.490 101.280 ;
        RECT 41.945 101.220 42.235 101.265 ;
        RECT 39.170 101.080 42.235 101.220 ;
        RECT 39.170 101.020 39.490 101.080 ;
        RECT 41.945 101.035 42.235 101.080 ;
        RECT 51.590 101.220 51.910 101.280 ;
        RECT 52.755 101.220 53.045 101.265 ;
        RECT 51.590 101.080 53.045 101.220 ;
        RECT 51.590 101.020 51.910 101.080 ;
        RECT 52.755 101.035 53.045 101.080 ;
        RECT 54.350 101.020 54.670 101.280 ;
        RECT 60.330 101.220 60.650 101.280 ;
        RECT 60.805 101.220 61.095 101.265 ;
        RECT 60.330 101.080 61.095 101.220 ;
        RECT 60.330 101.020 60.650 101.080 ;
        RECT 60.805 101.035 61.095 101.080 ;
        RECT 61.710 101.020 62.030 101.280 ;
        RECT 65.940 101.220 66.080 101.760 ;
        RECT 67.690 101.700 68.010 101.960 ;
        RECT 68.240 101.900 68.380 102.100 ;
        RECT 70.970 102.055 71.260 102.100 ;
        RECT 75.510 102.040 75.830 102.300 ;
        RECT 79.650 102.040 79.970 102.300 ;
        RECT 81.580 102.285 81.720 102.440 ;
        RECT 87.030 102.580 87.320 102.625 ;
        RECT 88.890 102.580 89.180 102.625 ;
        RECT 87.030 102.440 89.180 102.580 ;
        RECT 87.030 102.395 87.320 102.440 ;
        RECT 88.890 102.395 89.180 102.440 ;
        RECT 89.810 102.580 90.100 102.625 ;
        RECT 93.070 102.580 93.360 102.625 ;
        RECT 96.670 102.580 96.990 102.640 ;
        RECT 89.810 102.440 96.990 102.580 ;
        RECT 97.220 102.580 97.360 102.720 ;
        RECT 102.190 102.580 102.510 102.640 ;
        RECT 97.220 102.440 107.020 102.580 ;
        RECT 89.810 102.395 90.100 102.440 ;
        RECT 93.070 102.395 93.360 102.440 ;
        RECT 81.505 102.055 81.795 102.285 ;
        RECT 83.790 102.240 84.110 102.300 ;
        RECT 84.725 102.240 85.015 102.285 ;
        RECT 83.790 102.100 85.015 102.240 ;
        RECT 83.790 102.040 84.110 102.100 ;
        RECT 84.725 102.055 85.015 102.100 ;
        RECT 86.105 102.240 86.395 102.285 ;
        RECT 86.550 102.240 86.870 102.300 ;
        RECT 86.105 102.100 86.870 102.240 ;
        RECT 88.965 102.240 89.180 102.395 ;
        RECT 96.670 102.380 96.990 102.440 ;
        RECT 102.190 102.380 102.510 102.440 ;
        RECT 91.210 102.240 91.500 102.285 ;
        RECT 88.965 102.100 91.500 102.240 ;
        RECT 86.105 102.055 86.395 102.100 ;
        RECT 86.550 102.040 86.870 102.100 ;
        RECT 91.210 102.055 91.500 102.100 ;
        RECT 96.210 102.040 96.530 102.300 ;
        RECT 106.330 102.040 106.650 102.300 ;
        RECT 106.880 102.285 107.020 102.440 ;
        RECT 106.805 102.055 107.095 102.285 ;
        RECT 73.210 101.900 73.530 101.960 ;
        RECT 87.945 101.900 88.235 101.945 ;
        RECT 68.240 101.760 73.530 101.900 ;
        RECT 73.210 101.700 73.530 101.760 ;
        RECT 85.720 101.760 88.235 101.900 ;
        RECT 85.720 101.605 85.860 101.760 ;
        RECT 87.945 101.715 88.235 101.760 ;
        RECT 66.330 101.560 66.620 101.605 ;
        RECT 68.190 101.560 68.480 101.605 ;
        RECT 70.970 101.560 71.260 101.605 ;
        RECT 66.330 101.420 71.260 101.560 ;
        RECT 66.330 101.375 66.620 101.420 ;
        RECT 68.190 101.375 68.480 101.420 ;
        RECT 70.970 101.375 71.260 101.420 ;
        RECT 85.645 101.375 85.935 101.605 ;
        RECT 86.570 101.560 86.860 101.605 ;
        RECT 88.430 101.560 88.720 101.605 ;
        RECT 91.210 101.560 91.500 101.605 ;
        RECT 86.570 101.420 91.500 101.560 ;
        RECT 86.570 101.375 86.860 101.420 ;
        RECT 88.430 101.375 88.720 101.420 ;
        RECT 91.210 101.375 91.500 101.420 ;
        RECT 69.530 101.220 69.850 101.280 ;
        RECT 71.830 101.220 72.150 101.280 ;
        RECT 65.940 101.080 72.150 101.220 ;
        RECT 69.530 101.020 69.850 101.080 ;
        RECT 71.830 101.020 72.150 101.080 ;
        RECT 73.670 101.220 73.990 101.280 ;
        RECT 74.835 101.220 75.125 101.265 ;
        RECT 73.670 101.080 75.125 101.220 ;
        RECT 73.670 101.020 73.990 101.080 ;
        RECT 74.835 101.035 75.125 101.080 ;
        RECT 80.570 101.020 80.890 101.280 ;
        RECT 81.965 101.220 82.255 101.265 ;
        RECT 87.470 101.220 87.790 101.280 ;
        RECT 81.965 101.080 87.790 101.220 ;
        RECT 81.965 101.035 82.255 101.080 ;
        RECT 87.470 101.020 87.790 101.080 ;
        RECT 89.770 101.220 90.090 101.280 ;
        RECT 95.075 101.220 95.365 101.265 ;
        RECT 89.770 101.080 95.365 101.220 ;
        RECT 89.770 101.020 90.090 101.080 ;
        RECT 95.075 101.035 95.365 101.080 ;
        RECT 102.650 101.020 102.970 101.280 ;
        RECT 104.490 101.220 104.810 101.280 ;
        RECT 105.425 101.220 105.715 101.265 ;
        RECT 104.490 101.080 105.715 101.220 ;
        RECT 104.490 101.020 104.810 101.080 ;
        RECT 105.425 101.035 105.715 101.080 ;
        RECT 107.250 101.020 107.570 101.280 ;
        RECT 5.520 100.400 113.620 100.880 ;
        RECT 23.070 100.200 23.390 100.260 ;
        RECT 23.545 100.200 23.835 100.245 ;
        RECT 23.070 100.060 23.835 100.200 ;
        RECT 23.070 100.000 23.390 100.060 ;
        RECT 23.545 100.015 23.835 100.060 ;
        RECT 26.750 100.000 27.070 100.260 ;
        RECT 45.610 100.000 45.930 100.260 ;
        RECT 67.690 100.200 68.010 100.260 ;
        RECT 68.165 100.200 68.455 100.245 ;
        RECT 67.690 100.060 68.455 100.200 ;
        RECT 67.690 100.000 68.010 100.060 ;
        RECT 68.165 100.015 68.455 100.060 ;
        RECT 8.370 99.860 8.660 99.905 ;
        RECT 10.230 99.860 10.520 99.905 ;
        RECT 13.010 99.860 13.300 99.905 ;
        RECT 8.370 99.720 13.300 99.860 ;
        RECT 8.370 99.675 8.660 99.720 ;
        RECT 10.230 99.675 10.520 99.720 ;
        RECT 13.010 99.675 13.300 99.720 ;
        RECT 33.210 99.860 33.500 99.905 ;
        RECT 35.070 99.860 35.360 99.905 ;
        RECT 37.850 99.860 38.140 99.905 ;
        RECT 33.210 99.720 38.140 99.860 ;
        RECT 33.210 99.675 33.500 99.720 ;
        RECT 35.070 99.675 35.360 99.720 ;
        RECT 37.850 99.675 38.140 99.720 ;
        RECT 51.100 99.860 51.390 99.905 ;
        RECT 53.880 99.860 54.170 99.905 ;
        RECT 55.740 99.860 56.030 99.905 ;
        RECT 51.100 99.720 56.030 99.860 ;
        RECT 51.100 99.675 51.390 99.720 ;
        RECT 53.880 99.675 54.170 99.720 ;
        RECT 55.740 99.675 56.030 99.720 ;
        RECT 57.130 99.860 57.420 99.905 ;
        RECT 58.990 99.860 59.280 99.905 ;
        RECT 61.770 99.860 62.060 99.905 ;
        RECT 57.130 99.720 62.060 99.860 ;
        RECT 57.130 99.675 57.420 99.720 ;
        RECT 58.990 99.675 59.280 99.720 ;
        RECT 61.770 99.675 62.060 99.720 ;
        RECT 84.270 99.860 84.560 99.905 ;
        RECT 86.130 99.860 86.420 99.905 ;
        RECT 88.910 99.860 89.200 99.905 ;
        RECT 84.270 99.720 89.200 99.860 ;
        RECT 84.270 99.675 84.560 99.720 ;
        RECT 86.130 99.675 86.420 99.720 ;
        RECT 88.910 99.675 89.200 99.720 ;
        RECT 95.290 99.860 95.610 99.920 ;
        RECT 103.130 99.860 103.420 99.905 ;
        RECT 104.990 99.860 105.280 99.905 ;
        RECT 107.770 99.860 108.060 99.905 ;
        RECT 95.290 99.720 98.740 99.860 ;
        RECT 95.290 99.660 95.610 99.720 ;
        RECT 6.970 99.520 7.290 99.580 ;
        RECT 7.905 99.520 8.195 99.565 ;
        RECT 13.410 99.520 13.730 99.580 ;
        RECT 6.970 99.380 13.730 99.520 ;
        RECT 6.970 99.320 7.290 99.380 ;
        RECT 7.905 99.335 8.195 99.380 ;
        RECT 13.410 99.320 13.730 99.380 ;
        RECT 14.790 99.520 15.110 99.580 ;
        RECT 22.165 99.520 22.455 99.565 ;
        RECT 29.525 99.520 29.815 99.565 ;
        RECT 30.890 99.520 31.210 99.580 ;
        RECT 14.790 99.380 21.920 99.520 ;
        RECT 14.790 99.320 15.110 99.380 ;
        RECT 9.730 98.980 10.050 99.240 ;
        RECT 16.630 99.225 16.950 99.240 ;
        RECT 13.010 99.180 13.300 99.225 ;
        RECT 10.765 99.040 13.300 99.180 ;
        RECT 10.765 98.885 10.980 99.040 ;
        RECT 13.010 98.995 13.300 99.040 ;
        RECT 16.630 99.180 17.165 99.225 ;
        RECT 21.245 99.180 21.535 99.225 ;
        RECT 16.630 99.040 21.535 99.180 ;
        RECT 21.780 99.180 21.920 99.380 ;
        RECT 22.165 99.380 31.210 99.520 ;
        RECT 22.165 99.335 22.455 99.380 ;
        RECT 29.525 99.335 29.815 99.380 ;
        RECT 30.890 99.320 31.210 99.380 ;
        RECT 32.745 99.520 33.035 99.565 ;
        RECT 41.930 99.520 42.250 99.580 ;
        RECT 46.070 99.520 46.390 99.580 ;
        RECT 32.745 99.380 46.390 99.520 ;
        RECT 32.745 99.335 33.035 99.380 ;
        RECT 41.930 99.320 42.250 99.380 ;
        RECT 46.070 99.320 46.390 99.380 ;
        RECT 53.430 99.520 53.750 99.580 ;
        RECT 56.205 99.520 56.495 99.565 ;
        RECT 56.665 99.520 56.955 99.565 ;
        RECT 53.430 99.380 56.955 99.520 ;
        RECT 53.430 99.320 53.750 99.380 ;
        RECT 56.205 99.335 56.495 99.380 ;
        RECT 56.665 99.335 56.955 99.380 ;
        RECT 80.570 99.520 80.890 99.580 ;
        RECT 85.645 99.520 85.935 99.565 ;
        RECT 80.570 99.380 85.935 99.520 ;
        RECT 80.570 99.320 80.890 99.380 ;
        RECT 85.645 99.335 85.935 99.380 ;
        RECT 87.010 99.520 87.330 99.580 ;
        RECT 98.600 99.565 98.740 99.720 ;
        RECT 103.130 99.720 108.060 99.860 ;
        RECT 103.130 99.675 103.420 99.720 ;
        RECT 104.990 99.675 105.280 99.720 ;
        RECT 107.770 99.675 108.060 99.720 ;
        RECT 87.010 99.380 96.900 99.520 ;
        RECT 87.010 99.320 87.330 99.380 ;
        RECT 23.070 99.180 23.390 99.240 ;
        RECT 24.005 99.180 24.295 99.225 ;
        RECT 21.780 99.040 24.295 99.180 ;
        RECT 16.630 98.995 17.165 99.040 ;
        RECT 21.245 98.995 21.535 99.040 ;
        RECT 16.630 98.980 16.950 98.995 ;
        RECT 23.070 98.980 23.390 99.040 ;
        RECT 24.005 98.995 24.295 99.040 ;
        RECT 26.305 99.180 26.595 99.225 ;
        RECT 27.210 99.180 27.530 99.240 ;
        RECT 26.305 99.040 27.530 99.180 ;
        RECT 26.305 98.995 26.595 99.040 ;
        RECT 27.210 98.980 27.530 99.040 ;
        RECT 28.605 99.180 28.895 99.225 ;
        RECT 29.970 99.180 30.290 99.240 ;
        RECT 28.605 99.040 30.290 99.180 ;
        RECT 28.605 98.995 28.895 99.040 ;
        RECT 29.970 98.980 30.290 99.040 ;
        RECT 31.350 98.980 31.670 99.240 ;
        RECT 34.585 99.180 34.875 99.225 ;
        RECT 37.850 99.180 38.140 99.225 ;
        RECT 32.360 99.040 34.875 99.180 ;
        RECT 8.830 98.840 9.120 98.885 ;
        RECT 10.690 98.840 10.980 98.885 ;
        RECT 8.830 98.700 10.980 98.840 ;
        RECT 8.830 98.655 9.120 98.700 ;
        RECT 10.690 98.655 10.980 98.700 ;
        RECT 11.610 98.840 11.900 98.885 ;
        RECT 12.490 98.840 12.810 98.900 ;
        RECT 14.870 98.840 15.160 98.885 ;
        RECT 11.610 98.700 15.160 98.840 ;
        RECT 11.610 98.655 11.900 98.700 ;
        RECT 12.490 98.640 12.810 98.700 ;
        RECT 14.870 98.655 15.160 98.700 ;
        RECT 20.785 98.840 21.075 98.885 ;
        RECT 22.610 98.840 22.930 98.900 ;
        RECT 29.065 98.840 29.355 98.885 ;
        RECT 20.785 98.700 29.355 98.840 ;
        RECT 20.785 98.655 21.075 98.700 ;
        RECT 22.610 98.640 22.930 98.700 ;
        RECT 29.065 98.655 29.355 98.700 ;
        RECT 18.470 98.500 18.790 98.560 ;
        RECT 18.945 98.500 19.235 98.545 ;
        RECT 18.470 98.360 19.235 98.500 ;
        RECT 18.470 98.300 18.790 98.360 ;
        RECT 18.945 98.315 19.235 98.360 ;
        RECT 23.990 98.500 24.310 98.560 ;
        RECT 32.360 98.545 32.500 99.040 ;
        RECT 34.585 98.995 34.875 99.040 ;
        RECT 35.605 99.040 38.140 99.180 ;
        RECT 35.605 98.885 35.820 99.040 ;
        RECT 37.850 98.995 38.140 99.040 ;
        RECT 42.390 98.980 42.710 99.240 ;
        RECT 46.530 98.980 46.850 99.240 ;
        RECT 47.450 98.980 47.770 99.240 ;
        RECT 51.100 99.180 51.390 99.225 ;
        RECT 51.100 99.040 53.635 99.180 ;
        RECT 51.100 98.995 51.390 99.040 ;
        RECT 33.670 98.840 33.960 98.885 ;
        RECT 35.530 98.840 35.820 98.885 ;
        RECT 33.670 98.700 35.820 98.840 ;
        RECT 33.670 98.655 33.960 98.700 ;
        RECT 35.530 98.655 35.820 98.700 ;
        RECT 36.450 98.840 36.740 98.885 ;
        RECT 39.170 98.840 39.490 98.900 ;
        RECT 41.470 98.885 41.790 98.900 ;
        RECT 39.710 98.840 40.000 98.885 ;
        RECT 36.450 98.700 40.000 98.840 ;
        RECT 36.450 98.655 36.740 98.700 ;
        RECT 39.170 98.640 39.490 98.700 ;
        RECT 39.710 98.655 40.000 98.700 ;
        RECT 41.470 98.840 42.005 98.885 ;
        RECT 47.540 98.840 47.680 98.980 ;
        RECT 52.510 98.885 52.830 98.900 ;
        RECT 41.470 98.700 47.680 98.840 ;
        RECT 49.240 98.840 49.530 98.885 ;
        RECT 52.500 98.840 52.830 98.885 ;
        RECT 49.240 98.700 52.830 98.840 ;
        RECT 41.470 98.655 42.005 98.700 ;
        RECT 49.240 98.655 49.530 98.700 ;
        RECT 52.500 98.655 52.830 98.700 ;
        RECT 53.420 98.885 53.635 99.040 ;
        RECT 54.350 98.980 54.670 99.240 ;
        RECT 58.490 98.980 58.810 99.240 ;
        RECT 61.770 99.180 62.060 99.225 ;
        RECT 59.525 99.040 62.060 99.180 ;
        RECT 59.525 98.885 59.740 99.040 ;
        RECT 61.770 98.995 62.060 99.040 ;
        RECT 69.070 98.980 69.390 99.240 ;
        RECT 73.210 98.980 73.530 99.240 ;
        RECT 76.890 99.180 77.210 99.240 ;
        RECT 83.805 99.180 84.095 99.225 ;
        RECT 88.910 99.180 89.200 99.225 ;
        RECT 76.890 99.040 84.095 99.180 ;
        RECT 76.890 98.980 77.210 99.040 ;
        RECT 83.805 98.995 84.095 99.040 ;
        RECT 86.665 99.040 89.200 99.180 ;
        RECT 53.420 98.840 53.710 98.885 ;
        RECT 55.280 98.840 55.570 98.885 ;
        RECT 53.420 98.700 55.570 98.840 ;
        RECT 53.420 98.655 53.710 98.700 ;
        RECT 55.280 98.655 55.570 98.700 ;
        RECT 57.590 98.840 57.880 98.885 ;
        RECT 59.450 98.840 59.740 98.885 ;
        RECT 57.590 98.700 59.740 98.840 ;
        RECT 57.590 98.655 57.880 98.700 ;
        RECT 59.450 98.655 59.740 98.700 ;
        RECT 60.330 98.885 60.650 98.900 ;
        RECT 86.665 98.885 86.880 99.040 ;
        RECT 88.910 98.995 89.200 99.040 ;
        RECT 94.845 99.180 95.135 99.225 ;
        RECT 94.845 99.040 96.440 99.180 ;
        RECT 94.845 98.995 95.135 99.040 ;
        RECT 60.330 98.840 60.660 98.885 ;
        RECT 63.630 98.840 63.920 98.885 ;
        RECT 60.330 98.700 63.920 98.840 ;
        RECT 60.330 98.655 60.660 98.700 ;
        RECT 63.630 98.655 63.920 98.700 ;
        RECT 84.730 98.840 85.020 98.885 ;
        RECT 86.590 98.840 86.880 98.885 ;
        RECT 84.730 98.700 86.880 98.840 ;
        RECT 84.730 98.655 85.020 98.700 ;
        RECT 86.590 98.655 86.880 98.700 ;
        RECT 87.470 98.885 87.790 98.900 ;
        RECT 87.470 98.840 87.800 98.885 ;
        RECT 90.770 98.840 91.060 98.885 ;
        RECT 87.470 98.700 91.060 98.840 ;
        RECT 87.470 98.655 87.800 98.700 ;
        RECT 90.770 98.655 91.060 98.700 ;
        RECT 41.470 98.640 41.790 98.655 ;
        RECT 52.510 98.640 52.830 98.655 ;
        RECT 60.330 98.640 60.650 98.655 ;
        RECT 87.470 98.640 87.790 98.655 ;
        RECT 25.385 98.500 25.675 98.545 ;
        RECT 23.990 98.360 25.675 98.500 ;
        RECT 23.990 98.300 24.310 98.360 ;
        RECT 25.385 98.315 25.675 98.360 ;
        RECT 32.285 98.315 32.575 98.545 ;
        RECT 43.325 98.500 43.615 98.545 ;
        RECT 44.690 98.500 45.010 98.560 ;
        RECT 43.325 98.360 45.010 98.500 ;
        RECT 43.325 98.315 43.615 98.360 ;
        RECT 44.690 98.300 45.010 98.360 ;
        RECT 46.530 98.500 46.850 98.560 ;
        RECT 47.235 98.500 47.525 98.545 ;
        RECT 46.530 98.360 47.525 98.500 ;
        RECT 46.530 98.300 46.850 98.360 ;
        RECT 47.235 98.315 47.525 98.360 ;
        RECT 62.630 98.500 62.950 98.560 ;
        RECT 65.635 98.500 65.925 98.545 ;
        RECT 62.630 98.360 65.925 98.500 ;
        RECT 62.630 98.300 62.950 98.360 ;
        RECT 65.635 98.315 65.925 98.360 ;
        RECT 89.310 98.500 89.630 98.560 ;
        RECT 92.775 98.500 93.065 98.545 ;
        RECT 89.310 98.360 93.065 98.500 ;
        RECT 89.310 98.300 89.630 98.360 ;
        RECT 92.775 98.315 93.065 98.360 ;
        RECT 93.450 98.500 93.770 98.560 ;
        RECT 96.300 98.545 96.440 99.040 ;
        RECT 93.925 98.500 94.215 98.545 ;
        RECT 93.450 98.360 94.215 98.500 ;
        RECT 93.450 98.300 93.770 98.360 ;
        RECT 93.925 98.315 94.215 98.360 ;
        RECT 96.225 98.315 96.515 98.545 ;
        RECT 96.760 98.500 96.900 99.380 ;
        RECT 98.525 99.335 98.815 99.565 ;
        RECT 99.445 99.520 99.735 99.565 ;
        RECT 104.030 99.520 104.350 99.580 ;
        RECT 99.445 99.380 104.350 99.520 ;
        RECT 99.445 99.335 99.735 99.380 ;
        RECT 104.030 99.320 104.350 99.380 ;
        RECT 104.490 99.320 104.810 99.580 ;
        RECT 98.050 99.180 98.370 99.240 ;
        RECT 100.365 99.180 100.655 99.225 ;
        RECT 102.650 99.180 102.970 99.240 ;
        RECT 107.770 99.180 108.060 99.225 ;
        RECT 98.050 99.040 102.970 99.180 ;
        RECT 98.050 98.980 98.370 99.040 ;
        RECT 100.365 98.995 100.655 99.040 ;
        RECT 102.650 98.980 102.970 99.040 ;
        RECT 105.525 99.040 108.060 99.180 ;
        RECT 99.890 98.840 100.210 98.900 ;
        RECT 105.525 98.885 105.740 99.040 ;
        RECT 107.770 98.995 108.060 99.040 ;
        RECT 98.140 98.700 100.210 98.840 ;
        RECT 98.140 98.545 98.280 98.700 ;
        RECT 99.890 98.640 100.210 98.700 ;
        RECT 103.590 98.840 103.880 98.885 ;
        RECT 105.450 98.840 105.740 98.885 ;
        RECT 103.590 98.700 105.740 98.840 ;
        RECT 103.590 98.655 103.880 98.700 ;
        RECT 105.450 98.655 105.740 98.700 ;
        RECT 106.370 98.840 106.660 98.885 ;
        RECT 107.250 98.840 107.570 98.900 ;
        RECT 109.630 98.840 109.920 98.885 ;
        RECT 106.370 98.700 109.920 98.840 ;
        RECT 106.370 98.655 106.660 98.700 ;
        RECT 107.250 98.640 107.570 98.700 ;
        RECT 109.630 98.655 109.920 98.700 ;
        RECT 98.065 98.500 98.355 98.545 ;
        RECT 96.760 98.360 98.355 98.500 ;
        RECT 98.065 98.315 98.355 98.360 ;
        RECT 111.635 98.500 111.925 98.545 ;
        RECT 111.635 98.360 113.920 98.500 ;
        RECT 111.635 98.315 111.925 98.360 ;
        RECT 5.520 97.680 113.620 98.160 ;
        RECT 9.730 97.480 10.050 97.540 ;
        RECT 11.125 97.480 11.415 97.525 ;
        RECT 9.730 97.340 11.415 97.480 ;
        RECT 9.730 97.280 10.050 97.340 ;
        RECT 11.125 97.295 11.415 97.340 ;
        RECT 12.490 97.480 12.810 97.540 ;
        RECT 13.425 97.480 13.715 97.525 ;
        RECT 12.490 97.340 13.715 97.480 ;
        RECT 12.490 97.280 12.810 97.340 ;
        RECT 13.425 97.295 13.715 97.340 ;
        RECT 17.550 97.280 17.870 97.540 ;
        RECT 31.350 97.480 31.670 97.540 ;
        RECT 33.205 97.480 33.495 97.525 ;
        RECT 31.350 97.340 33.495 97.480 ;
        RECT 31.350 97.280 31.670 97.340 ;
        RECT 33.205 97.295 33.495 97.340 ;
        RECT 35.045 97.480 35.335 97.525 ;
        RECT 41.470 97.480 41.790 97.540 ;
        RECT 35.045 97.340 41.790 97.480 ;
        RECT 35.045 97.295 35.335 97.340 ;
        RECT 41.470 97.280 41.790 97.340 ;
        RECT 52.510 97.480 52.830 97.540 ;
        RECT 58.045 97.480 58.335 97.525 ;
        RECT 52.510 97.340 58.335 97.480 ;
        RECT 52.510 97.280 52.830 97.340 ;
        RECT 58.045 97.295 58.335 97.340 ;
        RECT 58.490 97.480 58.810 97.540 ;
        RECT 59.885 97.480 60.175 97.525 ;
        RECT 73.210 97.480 73.530 97.540 ;
        RECT 76.890 97.480 77.210 97.540 ;
        RECT 58.490 97.340 60.175 97.480 ;
        RECT 58.490 97.280 58.810 97.340 ;
        RECT 59.885 97.295 60.175 97.340 ;
        RECT 65.480 97.340 77.210 97.480 ;
        RECT 14.330 97.140 14.650 97.200 ;
        RECT 12.120 97.000 14.650 97.140 ;
        RECT 12.120 96.845 12.260 97.000 ;
        RECT 14.330 96.940 14.650 97.000 ;
        RECT 33.650 97.140 33.970 97.200 ;
        RECT 35.505 97.140 35.795 97.185 ;
        RECT 33.650 97.000 35.795 97.140 ;
        RECT 33.650 96.940 33.970 97.000 ;
        RECT 35.505 96.955 35.795 97.000 ;
        RECT 38.710 97.140 39.030 97.200 ;
        RECT 39.580 97.140 39.870 97.185 ;
        RECT 42.840 97.140 43.130 97.185 ;
        RECT 38.710 97.000 43.130 97.140 ;
        RECT 38.710 96.940 39.030 97.000 ;
        RECT 39.580 96.955 39.870 97.000 ;
        RECT 42.840 96.955 43.130 97.000 ;
        RECT 43.760 97.140 44.050 97.185 ;
        RECT 45.620 97.140 45.910 97.185 ;
        RECT 43.760 97.000 45.910 97.140 ;
        RECT 43.760 96.955 44.050 97.000 ;
        RECT 45.620 96.955 45.910 97.000 ;
        RECT 46.070 97.140 46.390 97.200 ;
        RECT 53.430 97.140 53.750 97.200 ;
        RECT 46.070 97.000 53.750 97.140 ;
        RECT 12.045 96.615 12.335 96.845 ;
        RECT 13.885 96.800 14.175 96.845 ;
        RECT 14.790 96.800 15.110 96.860 ;
        RECT 13.885 96.660 15.110 96.800 ;
        RECT 13.885 96.615 14.175 96.660 ;
        RECT 14.790 96.600 15.110 96.660 ;
        RECT 18.470 96.600 18.790 96.860 ;
        RECT 18.945 96.615 19.235 96.845 ;
        RECT 13.410 96.460 13.730 96.520 ;
        RECT 19.020 96.460 19.160 96.615 ;
        RECT 20.310 96.600 20.630 96.860 ;
        RECT 23.070 96.800 23.390 96.860 ;
        RECT 37.790 96.845 38.110 96.860 ;
        RECT 30.445 96.800 30.735 96.845 ;
        RECT 23.070 96.660 30.735 96.800 ;
        RECT 23.070 96.600 23.390 96.660 ;
        RECT 30.445 96.615 30.735 96.660 ;
        RECT 37.575 96.615 38.110 96.845 ;
        RECT 41.440 96.800 41.730 96.845 ;
        RECT 43.760 96.800 43.975 96.955 ;
        RECT 46.070 96.940 46.390 97.000 ;
        RECT 41.440 96.660 43.975 96.800 ;
        RECT 41.440 96.615 41.730 96.660 ;
        RECT 37.790 96.600 38.110 96.615 ;
        RECT 44.690 96.600 45.010 96.860 ;
        RECT 46.620 96.845 46.760 97.000 ;
        RECT 53.430 96.940 53.750 97.000 ;
        RECT 46.545 96.615 46.835 96.845 ;
        RECT 46.990 96.600 47.310 96.860 ;
        RECT 57.570 96.800 57.890 96.860 ;
        RECT 58.505 96.800 58.795 96.845 ;
        RECT 57.570 96.660 58.795 96.800 ;
        RECT 57.570 96.600 57.890 96.660 ;
        RECT 58.505 96.615 58.795 96.660 ;
        RECT 60.805 96.800 61.095 96.845 ;
        RECT 61.710 96.800 62.030 96.860 ;
        RECT 65.480 96.845 65.620 97.340 ;
        RECT 73.210 97.280 73.530 97.340 ;
        RECT 76.890 97.280 77.210 97.340 ;
        RECT 79.650 97.480 79.970 97.540 ;
        RECT 83.345 97.480 83.635 97.525 ;
        RECT 79.650 97.340 83.635 97.480 ;
        RECT 79.650 97.280 79.970 97.340 ;
        RECT 83.345 97.295 83.635 97.340 ;
        RECT 83.790 97.480 84.110 97.540 ;
        RECT 87.485 97.480 87.775 97.525 ;
        RECT 83.790 97.340 87.775 97.480 ;
        RECT 83.790 97.280 84.110 97.340 ;
        RECT 87.485 97.295 87.775 97.340 ;
        RECT 89.310 97.480 89.630 97.540 ;
        RECT 89.785 97.480 90.075 97.525 ;
        RECT 98.050 97.480 98.370 97.540 ;
        RECT 89.310 97.340 90.075 97.480 ;
        RECT 89.310 97.280 89.630 97.340 ;
        RECT 89.785 97.295 90.075 97.340 ;
        RECT 91.700 97.340 98.370 97.480 ;
        RECT 69.070 97.185 69.390 97.200 ;
        RECT 66.330 97.140 66.620 97.185 ;
        RECT 68.190 97.140 68.480 97.185 ;
        RECT 66.330 97.000 68.480 97.140 ;
        RECT 66.330 96.955 66.620 97.000 ;
        RECT 68.190 96.955 68.480 97.000 ;
        RECT 60.805 96.660 62.030 96.800 ;
        RECT 60.805 96.615 61.095 96.660 ;
        RECT 61.710 96.600 62.030 96.660 ;
        RECT 65.405 96.615 65.695 96.845 ;
        RECT 68.265 96.800 68.480 96.955 ;
        RECT 69.070 97.140 69.400 97.185 ;
        RECT 72.370 97.140 72.660 97.185 ;
        RECT 77.810 97.140 78.130 97.200 ;
        RECT 69.070 97.000 72.660 97.140 ;
        RECT 69.070 96.955 69.400 97.000 ;
        RECT 72.370 96.955 72.660 97.000 ;
        RECT 76.980 97.000 78.130 97.140 ;
        RECT 69.070 96.940 69.390 96.955 ;
        RECT 70.510 96.800 70.800 96.845 ;
        RECT 68.265 96.660 70.800 96.800 ;
        RECT 70.510 96.615 70.800 96.660 ;
        RECT 75.050 96.600 75.370 96.860 ;
        RECT 76.980 96.845 77.120 97.000 ;
        RECT 77.810 96.940 78.130 97.000 ;
        RECT 78.285 97.140 78.575 97.185 ;
        RECT 78.730 97.140 79.050 97.200 ;
        RECT 82.870 97.140 83.190 97.200 ;
        RECT 78.285 97.000 79.050 97.140 ;
        RECT 78.285 96.955 78.575 97.000 ;
        RECT 78.730 96.940 79.050 97.000 ;
        RECT 79.740 97.000 83.190 97.140 ;
        RECT 79.740 96.845 79.880 97.000 ;
        RECT 82.870 96.940 83.190 97.000 ;
        RECT 86.550 97.140 86.870 97.200 ;
        RECT 88.390 97.140 88.710 97.200 ;
        RECT 91.700 97.140 91.840 97.340 ;
        RECT 98.050 97.280 98.370 97.340 ;
        RECT 99.890 97.480 100.210 97.540 ;
        RECT 100.595 97.480 100.885 97.525 ;
        RECT 99.890 97.340 100.885 97.480 ;
        RECT 99.890 97.280 100.210 97.340 ;
        RECT 100.595 97.295 100.885 97.340 ;
        RECT 106.330 97.480 106.650 97.540 ;
        RECT 107.265 97.480 107.555 97.525 ;
        RECT 106.330 97.340 107.555 97.480 ;
        RECT 106.330 97.280 106.650 97.340 ;
        RECT 107.265 97.295 107.555 97.340 ;
        RECT 86.550 97.000 91.840 97.140 ;
        RECT 86.550 96.940 86.870 97.000 ;
        RECT 88.390 96.940 88.710 97.000 ;
        RECT 75.985 96.800 76.275 96.845 ;
        RECT 75.600 96.660 76.275 96.800 ;
        RECT 30.890 96.460 31.210 96.520 ;
        RECT 36.425 96.460 36.715 96.505 ;
        RECT 41.930 96.460 42.250 96.520 ;
        RECT 47.910 96.460 48.230 96.520 ;
        RECT 13.410 96.320 22.380 96.460 ;
        RECT 13.410 96.260 13.730 96.320 ;
        RECT 22.240 95.840 22.380 96.320 ;
        RECT 30.890 96.320 48.230 96.460 ;
        RECT 30.890 96.260 31.210 96.320 ;
        RECT 36.425 96.275 36.715 96.320 ;
        RECT 41.930 96.260 42.250 96.320 ;
        RECT 47.910 96.260 48.230 96.320 ;
        RECT 67.230 96.260 67.550 96.520 ;
        RECT 72.290 96.460 72.610 96.520 ;
        RECT 74.375 96.460 74.665 96.505 ;
        RECT 75.600 96.460 75.740 96.660 ;
        RECT 75.985 96.615 76.275 96.660 ;
        RECT 76.445 96.615 76.735 96.845 ;
        RECT 76.905 96.615 77.195 96.845 ;
        RECT 79.665 96.800 79.955 96.845 ;
        RECT 77.440 96.660 79.955 96.800 ;
        RECT 72.290 96.320 75.740 96.460 ;
        RECT 72.290 96.260 72.610 96.320 ;
        RECT 74.375 96.275 74.665 96.320 ;
        RECT 41.440 96.120 41.730 96.165 ;
        RECT 44.220 96.120 44.510 96.165 ;
        RECT 46.080 96.120 46.370 96.165 ;
        RECT 41.440 95.980 46.370 96.120 ;
        RECT 41.440 95.935 41.730 95.980 ;
        RECT 44.220 95.935 44.510 95.980 ;
        RECT 46.080 95.935 46.370 95.980 ;
        RECT 53.430 95.920 53.750 96.180 ;
        RECT 65.870 96.120 66.160 96.165 ;
        RECT 67.730 96.120 68.020 96.165 ;
        RECT 70.510 96.120 70.800 96.165 ;
        RECT 65.870 95.980 70.800 96.120 ;
        RECT 65.870 95.935 66.160 95.980 ;
        RECT 67.730 95.935 68.020 95.980 ;
        RECT 70.510 95.935 70.800 95.980 ;
        RECT 75.970 96.120 76.290 96.180 ;
        RECT 76.520 96.120 76.660 96.615 ;
        RECT 77.440 96.460 77.580 96.660 ;
        RECT 79.665 96.615 79.955 96.660 ;
        RECT 80.570 96.600 80.890 96.860 ;
        RECT 85.185 96.800 85.475 96.845 ;
        RECT 88.850 96.800 89.170 96.860 ;
        RECT 85.185 96.660 89.170 96.800 ;
        RECT 85.185 96.615 85.475 96.660 ;
        RECT 75.970 95.980 76.660 96.120 ;
        RECT 76.980 96.320 77.580 96.460 ;
        RECT 78.745 96.460 79.035 96.505 ;
        RECT 85.260 96.460 85.400 96.615 ;
        RECT 88.850 96.600 89.170 96.660 ;
        RECT 89.325 96.800 89.615 96.845 ;
        RECT 89.770 96.800 90.090 96.860 ;
        RECT 91.700 96.845 91.840 97.000 ;
        RECT 92.550 97.140 92.840 97.185 ;
        RECT 94.410 97.140 94.700 97.185 ;
        RECT 92.550 97.000 94.700 97.140 ;
        RECT 92.550 96.955 92.840 97.000 ;
        RECT 94.410 96.955 94.700 97.000 ;
        RECT 95.330 97.140 95.620 97.185 ;
        RECT 98.590 97.140 98.880 97.185 ;
        RECT 101.745 97.140 102.035 97.185 ;
        RECT 95.330 97.000 102.035 97.140 ;
        RECT 95.330 96.955 95.620 97.000 ;
        RECT 98.590 96.955 98.880 97.000 ;
        RECT 101.745 96.955 102.035 97.000 ;
        RECT 89.325 96.660 90.090 96.800 ;
        RECT 89.325 96.615 89.615 96.660 ;
        RECT 89.770 96.600 90.090 96.660 ;
        RECT 91.625 96.615 91.915 96.845 ;
        RECT 93.450 96.600 93.770 96.860 ;
        RECT 94.485 96.800 94.700 96.955 ;
        RECT 96.730 96.800 97.020 96.845 ;
        RECT 94.485 96.660 97.020 96.800 ;
        RECT 96.730 96.615 97.020 96.660 ;
        RECT 97.220 96.660 101.960 96.800 ;
        RECT 78.745 96.320 85.400 96.460 ;
        RECT 75.970 95.920 76.290 95.980 ;
        RECT 22.150 95.780 22.470 95.840 ;
        RECT 26.765 95.780 27.055 95.825 ;
        RECT 22.150 95.640 27.055 95.780 ;
        RECT 22.150 95.580 22.470 95.640 ;
        RECT 26.765 95.595 27.055 95.640 ;
        RECT 29.970 95.580 30.290 95.840 ;
        RECT 65.390 95.780 65.710 95.840 ;
        RECT 76.980 95.780 77.120 96.320 ;
        RECT 78.745 96.275 79.035 96.320 ;
        RECT 85.630 96.260 85.950 96.520 ;
        RECT 86.565 96.460 86.855 96.505 ;
        RECT 90.705 96.460 90.995 96.505 ;
        RECT 94.370 96.460 94.690 96.520 ;
        RECT 86.565 96.320 94.690 96.460 ;
        RECT 86.565 96.275 86.855 96.320 ;
        RECT 90.705 96.275 90.995 96.320 ;
        RECT 94.370 96.260 94.690 96.320 ;
        RECT 95.290 96.460 95.610 96.520 ;
        RECT 97.220 96.460 97.360 96.660 ;
        RECT 95.290 96.320 97.360 96.460 ;
        RECT 101.820 96.460 101.960 96.660 ;
        RECT 102.190 96.600 102.510 96.860 ;
        RECT 105.425 96.800 105.715 96.845 ;
        RECT 113.780 96.800 113.920 98.360 ;
        RECT 102.740 96.660 113.920 96.800 ;
        RECT 102.740 96.460 102.880 96.660 ;
        RECT 105.425 96.615 105.715 96.660 ;
        RECT 101.820 96.320 102.880 96.460 ;
        RECT 95.290 96.260 95.610 96.320 ;
        RECT 104.490 96.260 104.810 96.520 ;
        RECT 104.950 96.260 105.270 96.520 ;
        RECT 92.090 96.120 92.380 96.165 ;
        RECT 93.950 96.120 94.240 96.165 ;
        RECT 96.730 96.120 97.020 96.165 ;
        RECT 92.090 95.980 97.020 96.120 ;
        RECT 92.090 95.935 92.380 95.980 ;
        RECT 93.950 95.935 94.240 95.980 ;
        RECT 96.730 95.935 97.020 95.980 ;
        RECT 65.390 95.640 77.120 95.780 ;
        RECT 65.390 95.580 65.710 95.640 ;
        RECT 5.520 94.960 113.620 95.440 ;
        RECT 14.330 94.560 14.650 94.820 ;
        RECT 38.710 94.760 39.030 94.820 ;
        RECT 41.945 94.760 42.235 94.805 ;
        RECT 38.710 94.620 42.235 94.760 ;
        RECT 38.710 94.560 39.030 94.620 ;
        RECT 41.945 94.575 42.235 94.620 ;
        RECT 42.390 94.760 42.710 94.820 ;
        RECT 44.705 94.760 44.995 94.805 ;
        RECT 42.390 94.620 44.995 94.760 ;
        RECT 42.390 94.560 42.710 94.620 ;
        RECT 44.705 94.575 44.995 94.620 ;
        RECT 49.290 94.560 49.610 94.820 ;
        RECT 53.890 94.560 54.210 94.820 ;
        RECT 67.230 94.760 67.550 94.820 ;
        RECT 67.705 94.760 67.995 94.805 ;
        RECT 67.230 94.620 67.995 94.760 ;
        RECT 67.230 94.560 67.550 94.620 ;
        RECT 67.705 94.575 67.995 94.620 ;
        RECT 102.190 94.760 102.510 94.820 ;
        RECT 102.190 94.620 110.470 94.760 ;
        RECT 102.190 94.560 102.510 94.620 ;
        RECT 22.630 94.420 22.920 94.465 ;
        RECT 24.490 94.420 24.780 94.465 ;
        RECT 27.270 94.420 27.560 94.465 ;
        RECT 95.290 94.420 95.610 94.480 ;
        RECT 22.630 94.280 27.560 94.420 ;
        RECT 22.630 94.235 22.920 94.280 ;
        RECT 24.490 94.235 24.780 94.280 ;
        RECT 27.270 94.235 27.560 94.280 ;
        RECT 46.160 94.280 47.680 94.420 ;
        RECT 17.565 94.080 17.855 94.125 ;
        RECT 23.070 94.080 23.390 94.140 ;
        RECT 17.565 93.940 23.390 94.080 ;
        RECT 17.565 93.895 17.855 93.940 ;
        RECT 23.070 93.880 23.390 93.940 ;
        RECT 23.990 93.880 24.310 94.140 ;
        RECT 12.045 93.555 12.335 93.785 ;
        RECT 13.885 93.740 14.175 93.785 ;
        RECT 14.790 93.740 15.110 93.800 ;
        RECT 13.885 93.600 15.110 93.740 ;
        RECT 13.885 93.555 14.175 93.600 ;
        RECT 12.120 93.400 12.260 93.555 ;
        RECT 14.790 93.540 15.110 93.600 ;
        RECT 16.185 93.740 16.475 93.785 ;
        RECT 16.630 93.740 16.950 93.800 ;
        RECT 16.185 93.600 16.950 93.740 ;
        RECT 16.185 93.555 16.475 93.600 ;
        RECT 16.630 93.540 16.950 93.600 ;
        RECT 22.150 93.540 22.470 93.800 ;
        RECT 27.270 93.740 27.560 93.785 ;
        RECT 25.025 93.600 27.560 93.740 ;
        RECT 18.930 93.400 19.250 93.460 ;
        RECT 25.025 93.445 25.240 93.600 ;
        RECT 27.270 93.555 27.560 93.600 ;
        RECT 42.405 93.740 42.695 93.785 ;
        RECT 42.850 93.740 43.170 93.800 ;
        RECT 46.160 93.740 46.300 94.280 ;
        RECT 46.530 94.080 46.850 94.140 ;
        RECT 47.005 94.080 47.295 94.125 ;
        RECT 46.530 93.940 47.295 94.080 ;
        RECT 46.530 93.880 46.850 93.940 ;
        RECT 47.005 93.895 47.295 93.940 ;
        RECT 42.405 93.600 46.300 93.740 ;
        RECT 42.405 93.555 42.695 93.600 ;
        RECT 42.850 93.540 43.170 93.600 ;
        RECT 12.120 93.260 19.250 93.400 ;
        RECT 18.930 93.200 19.250 93.260 ;
        RECT 23.090 93.400 23.380 93.445 ;
        RECT 24.950 93.400 25.240 93.445 ;
        RECT 23.090 93.260 25.240 93.400 ;
        RECT 23.090 93.215 23.380 93.260 ;
        RECT 24.950 93.215 25.240 93.260 ;
        RECT 25.870 93.400 26.160 93.445 ;
        RECT 29.130 93.400 29.420 93.445 ;
        RECT 29.970 93.400 30.290 93.460 ;
        RECT 25.870 93.260 30.290 93.400 ;
        RECT 47.080 93.400 47.220 93.895 ;
        RECT 47.540 93.740 47.680 94.280 ;
        RECT 86.180 94.280 95.610 94.420 ;
        RECT 47.910 94.080 48.230 94.140 ;
        RECT 51.130 94.080 51.450 94.140 ;
        RECT 47.910 93.940 51.450 94.080 ;
        RECT 47.910 93.880 48.230 93.940 ;
        RECT 51.130 93.880 51.450 93.940 ;
        RECT 51.590 93.880 51.910 94.140 ;
        RECT 57.570 94.080 57.890 94.140 ;
        RECT 53.520 93.940 57.890 94.080 ;
        RECT 49.765 93.740 50.055 93.785 ;
        RECT 53.520 93.740 53.660 93.940 ;
        RECT 57.570 93.880 57.890 93.940 ;
        RECT 83.805 94.080 84.095 94.125 ;
        RECT 85.630 94.080 85.950 94.140 ;
        RECT 86.180 94.125 86.320 94.280 ;
        RECT 95.290 94.220 95.610 94.280 ;
        RECT 100.365 94.420 100.655 94.465 ;
        RECT 101.290 94.420 101.580 94.465 ;
        RECT 103.150 94.420 103.440 94.465 ;
        RECT 105.930 94.420 106.220 94.465 ;
        RECT 100.365 94.280 101.040 94.420 ;
        RECT 100.365 94.235 100.655 94.280 ;
        RECT 83.805 93.940 85.950 94.080 ;
        RECT 83.805 93.895 84.095 93.940 ;
        RECT 85.630 93.880 85.950 93.940 ;
        RECT 86.105 93.895 86.395 94.125 ;
        RECT 88.405 94.080 88.695 94.125 ;
        RECT 89.770 94.080 90.090 94.140 ;
        RECT 88.405 93.940 90.090 94.080 ;
        RECT 88.405 93.895 88.695 93.940 ;
        RECT 89.770 93.880 90.090 93.940 ;
        RECT 98.050 94.080 98.370 94.140 ;
        RECT 100.900 94.080 101.040 94.280 ;
        RECT 101.290 94.280 106.220 94.420 ;
        RECT 101.290 94.235 101.580 94.280 ;
        RECT 103.150 94.235 103.440 94.280 ;
        RECT 105.930 94.235 106.220 94.280 ;
        RECT 104.950 94.080 105.270 94.140 ;
        RECT 109.795 94.080 110.085 94.125 ;
        RECT 98.050 93.940 100.120 94.080 ;
        RECT 100.900 93.940 102.880 94.080 ;
        RECT 98.050 93.880 98.370 93.940 ;
        RECT 47.540 93.600 53.660 93.740 ;
        RECT 53.890 93.740 54.210 93.800 ;
        RECT 55.285 93.740 55.575 93.785 ;
        RECT 53.890 93.600 55.575 93.740 ;
        RECT 49.765 93.555 50.055 93.600 ;
        RECT 53.890 93.540 54.210 93.600 ;
        RECT 55.285 93.555 55.575 93.600 ;
        RECT 55.745 93.555 56.035 93.785 ;
        RECT 68.625 93.740 68.915 93.785 ;
        RECT 70.450 93.740 70.770 93.800 ;
        RECT 68.625 93.600 70.770 93.740 ;
        RECT 68.625 93.555 68.915 93.600 ;
        RECT 52.065 93.400 52.355 93.445 ;
        RECT 55.820 93.400 55.960 93.555 ;
        RECT 70.450 93.540 70.770 93.600 ;
        RECT 72.750 93.540 73.070 93.800 ;
        RECT 82.870 93.740 83.190 93.800 ;
        RECT 85.185 93.740 85.475 93.785 ;
        RECT 87.010 93.740 87.330 93.800 ;
        RECT 87.485 93.740 87.775 93.785 ;
        RECT 82.870 93.600 87.775 93.740 ;
        RECT 82.870 93.540 83.190 93.600 ;
        RECT 85.185 93.555 85.475 93.600 ;
        RECT 87.010 93.540 87.330 93.600 ;
        RECT 87.485 93.555 87.775 93.600 ;
        RECT 91.150 93.540 91.470 93.800 ;
        RECT 99.445 93.555 99.735 93.785 ;
        RECT 99.980 93.740 100.120 93.940 ;
        RECT 102.740 93.785 102.880 93.940 ;
        RECT 104.950 93.940 110.085 94.080 ;
        RECT 110.330 94.080 110.470 94.620 ;
        RECT 110.330 93.940 110.700 94.080 ;
        RECT 104.950 93.880 105.270 93.940 ;
        RECT 109.795 93.895 110.085 93.940 ;
        RECT 110.560 93.800 110.700 93.940 ;
        RECT 100.825 93.740 101.115 93.785 ;
        RECT 99.980 93.600 101.115 93.740 ;
        RECT 100.825 93.555 101.115 93.600 ;
        RECT 102.665 93.555 102.955 93.785 ;
        RECT 105.930 93.740 106.220 93.785 ;
        RECT 103.685 93.600 106.220 93.740 ;
        RECT 47.080 93.260 55.960 93.400 ;
        RECT 99.520 93.400 99.660 93.555 ;
        RECT 103.685 93.445 103.900 93.600 ;
        RECT 105.930 93.555 106.220 93.600 ;
        RECT 110.470 93.540 110.790 93.800 ;
        RECT 101.750 93.400 102.040 93.445 ;
        RECT 103.610 93.400 103.900 93.445 ;
        RECT 99.520 93.260 101.500 93.400 ;
        RECT 25.870 93.215 26.160 93.260 ;
        RECT 29.130 93.215 29.420 93.260 ;
        RECT 29.970 93.200 30.290 93.260 ;
        RECT 52.065 93.215 52.355 93.260 ;
        RECT 9.730 93.060 10.050 93.120 ;
        RECT 11.125 93.060 11.415 93.105 ;
        RECT 9.730 92.920 11.415 93.060 ;
        RECT 9.730 92.860 10.050 92.920 ;
        RECT 11.125 92.875 11.415 92.920 ;
        RECT 12.490 93.060 12.810 93.120 ;
        RECT 13.425 93.060 13.715 93.105 ;
        RECT 12.490 92.920 13.715 93.060 ;
        RECT 12.490 92.860 12.810 92.920 ;
        RECT 13.425 92.875 13.715 92.920 ;
        RECT 16.645 93.060 16.935 93.105 ;
        RECT 20.770 93.060 21.090 93.120 ;
        RECT 16.645 92.920 21.090 93.060 ;
        RECT 16.645 92.875 16.935 92.920 ;
        RECT 20.770 92.860 21.090 92.920 ;
        RECT 30.430 93.060 30.750 93.120 ;
        RECT 31.135 93.060 31.425 93.105 ;
        RECT 30.430 92.920 31.425 93.060 ;
        RECT 30.430 92.860 30.750 92.920 ;
        RECT 31.135 92.875 31.425 92.920 ;
        RECT 41.010 93.060 41.330 93.120 ;
        RECT 46.545 93.060 46.835 93.105 ;
        RECT 41.010 92.920 46.835 93.060 ;
        RECT 41.010 92.860 41.330 92.920 ;
        RECT 46.545 92.875 46.835 92.920 ;
        RECT 52.510 93.060 52.830 93.120 ;
        RECT 54.365 93.060 54.655 93.105 ;
        RECT 52.510 92.920 54.655 93.060 ;
        RECT 52.510 92.860 52.830 92.920 ;
        RECT 54.365 92.875 54.655 92.920 ;
        RECT 76.890 93.060 77.210 93.120 ;
        RECT 79.205 93.060 79.495 93.105 ;
        RECT 76.890 92.920 79.495 93.060 ;
        RECT 76.890 92.860 77.210 92.920 ;
        RECT 79.205 92.875 79.495 92.920 ;
        RECT 81.030 93.060 81.350 93.120 ;
        RECT 81.965 93.060 82.255 93.105 ;
        RECT 81.030 92.920 82.255 93.060 ;
        RECT 81.030 92.860 81.350 92.920 ;
        RECT 81.965 92.875 82.255 92.920 ;
        RECT 82.870 93.060 83.190 93.120 ;
        RECT 84.265 93.060 84.555 93.105 ;
        RECT 82.870 92.920 84.555 93.060 ;
        RECT 82.870 92.860 83.190 92.920 ;
        RECT 84.265 92.875 84.555 92.920 ;
        RECT 86.550 92.860 86.870 93.120 ;
        RECT 90.230 92.860 90.550 93.120 ;
        RECT 101.360 93.060 101.500 93.260 ;
        RECT 101.750 93.260 103.900 93.400 ;
        RECT 101.750 93.215 102.040 93.260 ;
        RECT 103.610 93.215 103.900 93.260 ;
        RECT 104.530 93.400 104.820 93.445 ;
        RECT 107.790 93.400 108.080 93.445 ;
        RECT 110.945 93.400 111.235 93.445 ;
        RECT 104.530 93.260 111.235 93.400 ;
        RECT 104.530 93.215 104.820 93.260 ;
        RECT 107.790 93.215 108.080 93.260 ;
        RECT 110.945 93.215 111.235 93.260 ;
        RECT 106.330 93.060 106.650 93.120 ;
        RECT 101.360 92.920 106.650 93.060 ;
        RECT 106.330 92.860 106.650 92.920 ;
        RECT 5.520 92.240 113.620 92.720 ;
        RECT 27.210 91.840 27.530 92.100 ;
        RECT 29.065 92.040 29.355 92.085 ;
        RECT 30.430 92.040 30.750 92.100 ;
        RECT 29.065 91.900 30.750 92.040 ;
        RECT 29.065 91.855 29.355 91.900 ;
        RECT 8.830 91.700 9.120 91.745 ;
        RECT 10.690 91.700 10.980 91.745 ;
        RECT 8.830 91.560 10.980 91.700 ;
        RECT 8.830 91.515 9.120 91.560 ;
        RECT 10.690 91.515 10.980 91.560 ;
        RECT 11.610 91.700 11.900 91.745 ;
        RECT 12.490 91.700 12.810 91.760 ;
        RECT 14.870 91.700 15.160 91.745 ;
        RECT 11.610 91.560 15.160 91.700 ;
        RECT 11.610 91.515 11.900 91.560 ;
        RECT 9.730 91.160 10.050 91.420 ;
        RECT 10.765 91.360 10.980 91.515 ;
        RECT 12.490 91.500 12.810 91.560 ;
        RECT 14.870 91.515 15.160 91.560 ;
        RECT 19.865 91.700 20.155 91.745 ;
        RECT 19.865 91.560 27.440 91.700 ;
        RECT 19.865 91.515 20.155 91.560 ;
        RECT 27.300 91.420 27.440 91.560 ;
        RECT 13.010 91.360 13.300 91.405 ;
        RECT 10.765 91.220 13.300 91.360 ;
        RECT 13.010 91.175 13.300 91.220 ;
        RECT 19.390 91.160 19.710 91.420 ;
        RECT 22.610 91.360 22.930 91.420 ;
        RECT 24.465 91.360 24.755 91.405 ;
        RECT 22.610 91.220 24.755 91.360 ;
        RECT 22.610 91.160 22.930 91.220 ;
        RECT 24.465 91.175 24.755 91.220 ;
        RECT 25.385 91.175 25.675 91.405 ;
        RECT 27.210 91.360 27.530 91.420 ;
        RECT 29.140 91.360 29.280 91.855 ;
        RECT 30.430 91.840 30.750 91.900 ;
        RECT 51.130 92.040 51.450 92.100 ;
        RECT 58.045 92.040 58.335 92.085 ;
        RECT 51.130 91.900 58.335 92.040 ;
        RECT 51.130 91.840 51.450 91.900 ;
        RECT 58.045 91.855 58.335 91.900 ;
        RECT 69.070 92.040 69.390 92.100 ;
        RECT 69.545 92.040 69.835 92.085 ;
        RECT 69.070 91.900 69.835 92.040 ;
        RECT 69.070 91.840 69.390 91.900 ;
        RECT 69.545 91.855 69.835 91.900 ;
        RECT 70.450 91.840 70.770 92.100 ;
        RECT 72.290 92.040 72.610 92.100 ;
        RECT 72.765 92.040 73.055 92.085 ;
        RECT 72.290 91.900 73.055 92.040 ;
        RECT 72.290 91.840 72.610 91.900 ;
        RECT 72.765 91.855 73.055 91.900 ;
        RECT 79.190 92.040 79.510 92.100 ;
        RECT 81.505 92.040 81.795 92.085 ;
        RECT 104.950 92.040 105.270 92.100 ;
        RECT 79.190 91.900 81.795 92.040 ;
        RECT 79.190 91.840 79.510 91.900 ;
        RECT 81.505 91.855 81.795 91.900 ;
        RECT 88.020 91.900 105.270 92.040 ;
        RECT 29.525 91.700 29.815 91.745 ;
        RECT 37.790 91.700 38.110 91.760 ;
        RECT 41.010 91.700 41.330 91.760 ;
        RECT 59.425 91.700 59.715 91.745 ;
        RECT 60.345 91.700 60.635 91.745 ;
        RECT 83.805 91.700 84.095 91.745 ;
        RECT 29.525 91.560 48.600 91.700 ;
        RECT 29.525 91.515 29.815 91.560 ;
        RECT 37.790 91.500 38.110 91.560 ;
        RECT 41.010 91.500 41.330 91.560 ;
        RECT 32.745 91.360 33.035 91.405 ;
        RECT 33.190 91.360 33.510 91.420 ;
        RECT 27.210 91.220 29.280 91.360 ;
        RECT 29.600 91.220 33.510 91.360 ;
        RECT 7.905 91.020 8.195 91.065 ;
        RECT 8.810 91.020 9.130 91.080 ;
        RECT 7.905 90.880 9.130 91.020 ;
        RECT 7.905 90.835 8.195 90.880 ;
        RECT 8.810 90.820 9.130 90.880 ;
        RECT 20.325 91.020 20.615 91.065 ;
        RECT 23.070 91.020 23.390 91.080 ;
        RECT 25.460 91.020 25.600 91.175 ;
        RECT 27.210 91.160 27.530 91.220 ;
        RECT 29.600 91.020 29.740 91.220 ;
        RECT 32.745 91.175 33.035 91.220 ;
        RECT 33.190 91.160 33.510 91.220 ;
        RECT 33.650 91.160 33.970 91.420 ;
        RECT 48.460 91.405 48.600 91.560 ;
        RECT 59.425 91.560 84.095 91.700 ;
        RECT 59.425 91.515 59.715 91.560 ;
        RECT 60.345 91.515 60.635 91.560 ;
        RECT 83.805 91.515 84.095 91.560 ;
        RECT 48.385 91.175 48.675 91.405 ;
        RECT 49.305 91.360 49.595 91.405 ;
        RECT 51.605 91.360 51.895 91.405 ;
        RECT 49.305 91.220 51.895 91.360 ;
        RECT 49.305 91.175 49.595 91.220 ;
        RECT 51.605 91.175 51.895 91.220 ;
        RECT 52.050 91.360 52.370 91.420 ;
        RECT 52.985 91.360 53.275 91.405 ;
        RECT 52.050 91.220 53.275 91.360 ;
        RECT 20.325 90.880 25.140 91.020 ;
        RECT 25.460 90.880 29.740 91.020 ;
        RECT 30.445 91.020 30.735 91.065 ;
        RECT 41.930 91.020 42.250 91.080 ;
        RECT 30.445 90.880 42.250 91.020 ;
        RECT 20.325 90.835 20.615 90.880 ;
        RECT 23.070 90.820 23.390 90.880 ;
        RECT 8.370 90.680 8.660 90.725 ;
        RECT 10.230 90.680 10.520 90.725 ;
        RECT 13.010 90.680 13.300 90.725 ;
        RECT 8.370 90.540 13.300 90.680 ;
        RECT 8.370 90.495 8.660 90.540 ;
        RECT 10.230 90.495 10.520 90.540 ;
        RECT 13.010 90.495 13.300 90.540 ;
        RECT 16.875 90.680 17.165 90.725 ;
        RECT 20.770 90.680 21.090 90.740 ;
        RECT 16.875 90.540 21.090 90.680 ;
        RECT 25.000 90.680 25.140 90.880 ;
        RECT 30.445 90.835 30.735 90.880 ;
        RECT 30.520 90.680 30.660 90.835 ;
        RECT 41.930 90.820 42.250 90.880 ;
        RECT 47.450 91.020 47.770 91.080 ;
        RECT 50.685 91.020 50.975 91.065 ;
        RECT 47.450 90.880 50.975 91.020 ;
        RECT 51.680 91.020 51.820 91.175 ;
        RECT 52.050 91.160 52.370 91.220 ;
        RECT 52.985 91.175 53.275 91.220 ;
        RECT 53.890 91.160 54.210 91.420 ;
        RECT 60.790 91.360 61.110 91.420 ;
        RECT 61.265 91.360 61.555 91.405 ;
        RECT 60.790 91.220 61.555 91.360 ;
        RECT 60.790 91.160 61.110 91.220 ;
        RECT 61.265 91.175 61.555 91.220 ;
        RECT 62.170 91.160 62.490 91.420 ;
        RECT 63.565 91.360 63.855 91.405 ;
        RECT 64.470 91.360 64.790 91.420 ;
        RECT 63.565 91.220 64.790 91.360 ;
        RECT 63.565 91.175 63.855 91.220 ;
        RECT 64.470 91.160 64.790 91.220 ;
        RECT 69.070 91.160 69.390 91.420 ;
        RECT 72.290 91.160 72.610 91.420 ;
        RECT 74.590 91.360 74.910 91.420 ;
        RECT 75.525 91.360 75.815 91.405 ;
        RECT 74.590 91.220 75.815 91.360 ;
        RECT 74.590 91.160 74.910 91.220 ;
        RECT 75.525 91.175 75.815 91.220 ;
        RECT 76.445 91.175 76.735 91.405 ;
        RECT 76.905 91.175 77.195 91.405 ;
        RECT 77.365 91.175 77.655 91.405 ;
        RECT 77.810 91.360 78.130 91.420 ;
        RECT 79.205 91.360 79.495 91.405 ;
        RECT 77.810 91.220 79.495 91.360 ;
        RECT 53.980 91.020 54.120 91.160 ;
        RECT 65.390 91.020 65.710 91.080 ;
        RECT 51.680 90.880 65.710 91.020 ;
        RECT 47.450 90.820 47.770 90.880 ;
        RECT 50.685 90.835 50.975 90.880 ;
        RECT 65.390 90.820 65.710 90.880 ;
        RECT 71.830 91.020 72.150 91.080 ;
        RECT 73.210 91.020 73.530 91.080 ;
        RECT 71.830 90.880 73.530 91.020 ;
        RECT 71.830 90.820 72.150 90.880 ;
        RECT 73.210 90.820 73.530 90.880 ;
        RECT 73.670 91.020 73.990 91.080 ;
        RECT 76.520 91.020 76.660 91.175 ;
        RECT 73.670 90.880 76.660 91.020 ;
        RECT 73.670 90.820 73.990 90.880 ;
        RECT 25.000 90.540 30.660 90.680 ;
        RECT 75.970 90.680 76.290 90.740 ;
        RECT 76.980 90.680 77.120 91.175 ;
        RECT 77.440 91.020 77.580 91.175 ;
        RECT 77.810 91.160 78.130 91.220 ;
        RECT 79.205 91.175 79.495 91.220 ;
        RECT 80.585 91.360 80.875 91.405 ;
        RECT 81.950 91.360 82.270 91.420 ;
        RECT 80.585 91.220 82.270 91.360 ;
        RECT 80.585 91.175 80.875 91.220 ;
        RECT 81.950 91.160 82.270 91.220 ;
        RECT 85.645 91.360 85.935 91.405 ;
        RECT 85.645 91.220 86.780 91.360 ;
        RECT 85.645 91.175 85.935 91.220 ;
        RECT 78.270 91.020 78.590 91.080 ;
        RECT 77.440 90.880 78.590 91.020 ;
        RECT 78.270 90.820 78.590 90.880 ;
        RECT 80.110 90.820 80.430 91.080 ;
        RECT 83.790 91.020 84.110 91.080 ;
        RECT 86.105 91.020 86.395 91.065 ;
        RECT 83.790 90.880 86.395 91.020 ;
        RECT 86.640 91.020 86.780 91.220 ;
        RECT 87.010 91.160 87.330 91.420 ;
        RECT 88.020 91.405 88.160 91.900 ;
        RECT 104.950 91.840 105.270 91.900 ;
        RECT 95.290 91.745 95.610 91.760 ;
        RECT 89.330 91.700 89.620 91.745 ;
        RECT 91.190 91.700 91.480 91.745 ;
        RECT 89.330 91.560 91.480 91.700 ;
        RECT 89.330 91.515 89.620 91.560 ;
        RECT 91.190 91.515 91.480 91.560 ;
        RECT 92.110 91.700 92.400 91.745 ;
        RECT 95.290 91.700 95.660 91.745 ;
        RECT 92.110 91.560 95.660 91.700 ;
        RECT 92.110 91.515 92.400 91.560 ;
        RECT 95.290 91.515 95.660 91.560 ;
        RECT 99.910 91.700 100.200 91.745 ;
        RECT 101.770 91.700 102.060 91.745 ;
        RECT 99.910 91.560 102.060 91.700 ;
        RECT 99.910 91.515 100.200 91.560 ;
        RECT 101.770 91.515 102.060 91.560 ;
        RECT 102.690 91.700 102.980 91.745 ;
        RECT 105.950 91.700 106.240 91.745 ;
        RECT 110.945 91.700 111.235 91.745 ;
        RECT 102.690 91.560 111.235 91.700 ;
        RECT 102.690 91.515 102.980 91.560 ;
        RECT 105.950 91.515 106.240 91.560 ;
        RECT 110.945 91.515 111.235 91.560 ;
        RECT 87.945 91.175 88.235 91.405 ;
        RECT 88.390 91.160 88.710 91.420 ;
        RECT 90.230 91.160 90.550 91.420 ;
        RECT 91.265 91.360 91.480 91.515 ;
        RECT 95.290 91.500 95.610 91.515 ;
        RECT 93.510 91.360 93.800 91.405 ;
        RECT 91.265 91.220 93.800 91.360 ;
        RECT 93.510 91.175 93.800 91.220 ;
        RECT 98.050 91.360 98.370 91.420 ;
        RECT 98.985 91.360 99.275 91.405 ;
        RECT 98.050 91.220 99.275 91.360 ;
        RECT 101.845 91.360 102.060 91.515 ;
        RECT 104.090 91.360 104.380 91.405 ;
        RECT 101.845 91.220 104.380 91.360 ;
        RECT 98.050 91.160 98.370 91.220 ;
        RECT 98.985 91.175 99.275 91.220 ;
        RECT 104.090 91.175 104.380 91.220 ;
        RECT 110.010 91.160 110.330 91.420 ;
        RECT 110.470 91.160 110.790 91.420 ;
        RECT 94.370 91.020 94.690 91.080 ;
        RECT 86.640 90.880 94.690 91.020 ;
        RECT 83.790 90.820 84.110 90.880 ;
        RECT 86.105 90.835 86.395 90.880 ;
        RECT 94.370 90.820 94.690 90.880 ;
        RECT 100.825 91.020 101.115 91.065 ;
        RECT 100.825 90.880 109.320 91.020 ;
        RECT 100.825 90.835 101.115 90.880 ;
        RECT 75.970 90.540 77.120 90.680 ;
        RECT 78.745 90.680 79.035 90.725 ;
        RECT 85.170 90.680 85.490 90.740 ;
        RECT 109.180 90.725 109.320 90.880 ;
        RECT 78.745 90.540 85.490 90.680 ;
        RECT 16.875 90.495 17.165 90.540 ;
        RECT 20.770 90.480 21.090 90.540 ;
        RECT 75.970 90.480 76.290 90.540 ;
        RECT 78.745 90.495 79.035 90.540 ;
        RECT 85.170 90.480 85.490 90.540 ;
        RECT 88.870 90.680 89.160 90.725 ;
        RECT 90.730 90.680 91.020 90.725 ;
        RECT 93.510 90.680 93.800 90.725 ;
        RECT 88.870 90.540 93.800 90.680 ;
        RECT 88.870 90.495 89.160 90.540 ;
        RECT 90.730 90.495 91.020 90.540 ;
        RECT 93.510 90.495 93.800 90.540 ;
        RECT 99.450 90.680 99.740 90.725 ;
        RECT 101.310 90.680 101.600 90.725 ;
        RECT 104.090 90.680 104.380 90.725 ;
        RECT 99.450 90.540 104.380 90.680 ;
        RECT 99.450 90.495 99.740 90.540 ;
        RECT 101.310 90.495 101.600 90.540 ;
        RECT 104.090 90.495 104.380 90.540 ;
        RECT 109.105 90.495 109.395 90.725 ;
        RECT 17.550 90.140 17.870 90.400 ;
        RECT 26.305 90.340 26.595 90.385 ;
        RECT 26.750 90.340 27.070 90.400 ;
        RECT 26.305 90.200 27.070 90.340 ;
        RECT 26.305 90.155 26.595 90.200 ;
        RECT 26.750 90.140 27.070 90.200 ;
        RECT 31.810 90.140 32.130 90.400 ;
        RECT 50.225 90.340 50.515 90.385 ;
        RECT 50.670 90.340 50.990 90.400 ;
        RECT 50.225 90.200 50.990 90.340 ;
        RECT 50.225 90.155 50.515 90.200 ;
        RECT 50.670 90.140 50.990 90.200 ;
        RECT 51.590 90.340 51.910 90.400 ;
        RECT 52.525 90.340 52.815 90.385 ;
        RECT 51.590 90.200 52.815 90.340 ;
        RECT 51.590 90.140 51.910 90.200 ;
        RECT 52.525 90.155 52.815 90.200 ;
        RECT 53.890 90.340 54.210 90.400 ;
        RECT 54.825 90.340 55.115 90.385 ;
        RECT 53.890 90.200 55.115 90.340 ;
        RECT 53.890 90.140 54.210 90.200 ;
        RECT 54.825 90.155 55.115 90.200 ;
        RECT 63.090 90.140 63.410 90.400 ;
        RECT 80.585 90.340 80.875 90.385 ;
        RECT 81.030 90.340 81.350 90.400 ;
        RECT 80.585 90.200 81.350 90.340 ;
        RECT 80.585 90.155 80.875 90.200 ;
        RECT 81.030 90.140 81.350 90.200 ;
        RECT 96.670 90.340 96.990 90.400 ;
        RECT 97.375 90.340 97.665 90.385 ;
        RECT 96.670 90.200 97.665 90.340 ;
        RECT 96.670 90.140 96.990 90.200 ;
        RECT 97.375 90.155 97.665 90.200 ;
        RECT 107.955 90.340 108.245 90.385 ;
        RECT 108.630 90.340 108.950 90.400 ;
        RECT 107.955 90.200 108.950 90.340 ;
        RECT 107.955 90.155 108.245 90.200 ;
        RECT 108.630 90.140 108.950 90.200 ;
        RECT 5.520 89.520 113.620 90.000 ;
        RECT 18.930 89.120 19.250 89.380 ;
        RECT 48.830 89.320 49.150 89.380 ;
        RECT 49.305 89.320 49.595 89.365 ;
        RECT 48.830 89.180 49.595 89.320 ;
        RECT 48.830 89.120 49.150 89.180 ;
        RECT 49.305 89.135 49.595 89.180 ;
        RECT 51.590 89.120 51.910 89.380 ;
        RECT 65.390 89.120 65.710 89.380 ;
        RECT 77.365 89.320 77.655 89.365 ;
        RECT 77.810 89.320 78.130 89.380 ;
        RECT 77.365 89.180 78.130 89.320 ;
        RECT 77.365 89.135 77.655 89.180 ;
        RECT 77.810 89.120 78.130 89.180 ;
        RECT 79.665 89.135 79.955 89.365 ;
        RECT 80.570 89.320 80.890 89.380 ;
        RECT 81.045 89.320 81.335 89.365 ;
        RECT 80.570 89.180 81.335 89.320 ;
        RECT 9.290 88.980 9.580 89.025 ;
        RECT 11.150 88.980 11.440 89.025 ;
        RECT 13.930 88.980 14.220 89.025 ;
        RECT 9.290 88.840 14.220 88.980 ;
        RECT 9.290 88.795 9.580 88.840 ;
        RECT 11.150 88.795 11.440 88.840 ;
        RECT 13.930 88.795 14.220 88.840 ;
        RECT 17.795 88.980 18.085 89.025 ;
        RECT 19.390 88.980 19.710 89.040 ;
        RECT 51.130 88.980 51.450 89.040 ;
        RECT 17.795 88.840 21.460 88.980 ;
        RECT 17.795 88.795 18.085 88.840 ;
        RECT 19.390 88.780 19.710 88.840 ;
        RECT 8.810 88.640 9.130 88.700 ;
        RECT 13.410 88.640 13.730 88.700 ;
        RECT 21.320 88.685 21.460 88.840 ;
        RECT 50.760 88.840 51.450 88.980 ;
        RECT 8.810 88.500 13.730 88.640 ;
        RECT 8.810 88.440 9.130 88.500 ;
        RECT 13.410 88.440 13.730 88.500 ;
        RECT 21.245 88.455 21.535 88.685 ;
        RECT 22.165 88.640 22.455 88.685 ;
        RECT 23.070 88.640 23.390 88.700 ;
        RECT 33.190 88.640 33.510 88.700 ;
        RECT 49.750 88.640 50.070 88.700 ;
        RECT 50.760 88.685 50.900 88.840 ;
        RECT 51.130 88.780 51.450 88.840 ;
        RECT 55.290 88.980 55.580 89.025 ;
        RECT 57.150 88.980 57.440 89.025 ;
        RECT 59.930 88.980 60.220 89.025 ;
        RECT 55.290 88.840 60.220 88.980 ;
        RECT 79.740 88.980 79.880 89.135 ;
        RECT 80.570 89.120 80.890 89.180 ;
        RECT 81.045 89.135 81.335 89.180 ;
        RECT 83.330 89.120 83.650 89.380 ;
        RECT 86.550 89.120 86.870 89.380 ;
        RECT 87.485 89.320 87.775 89.365 ;
        RECT 87.930 89.320 88.250 89.380 ;
        RECT 87.485 89.180 88.250 89.320 ;
        RECT 87.485 89.135 87.775 89.180 ;
        RECT 87.930 89.120 88.250 89.180 ;
        RECT 90.705 89.320 90.995 89.365 ;
        RECT 91.150 89.320 91.470 89.380 ;
        RECT 90.705 89.180 91.470 89.320 ;
        RECT 90.705 89.135 90.995 89.180 ;
        RECT 91.150 89.120 91.470 89.180 ;
        RECT 95.290 89.320 95.610 89.380 ;
        RECT 96.685 89.320 96.975 89.365 ;
        RECT 95.290 89.180 96.975 89.320 ;
        RECT 95.290 89.120 95.610 89.180 ;
        RECT 96.685 89.135 96.975 89.180 ;
        RECT 105.885 89.320 106.175 89.365 ;
        RECT 110.010 89.320 110.330 89.380 ;
        RECT 105.885 89.180 110.330 89.320 ;
        RECT 105.885 89.135 106.175 89.180 ;
        RECT 110.010 89.120 110.330 89.180 ;
        RECT 82.870 88.980 83.190 89.040 ;
        RECT 79.740 88.840 83.190 88.980 ;
        RECT 55.290 88.795 55.580 88.840 ;
        RECT 57.150 88.795 57.440 88.840 ;
        RECT 59.930 88.795 60.220 88.840 ;
        RECT 82.870 88.780 83.190 88.840 ;
        RECT 89.770 88.980 90.090 89.040 ;
        RECT 89.770 88.840 93.220 88.980 ;
        RECT 89.770 88.780 90.090 88.840 ;
        RECT 22.165 88.500 23.390 88.640 ;
        RECT 22.165 88.455 22.455 88.500 ;
        RECT 23.070 88.440 23.390 88.500 ;
        RECT 24.080 88.500 27.900 88.640 ;
        RECT 24.080 88.360 24.220 88.500 ;
        RECT 10.650 88.100 10.970 88.360 ;
        RECT 13.930 88.300 14.220 88.345 ;
        RECT 11.685 88.160 14.220 88.300 ;
        RECT 11.685 88.005 11.900 88.160 ;
        RECT 13.930 88.115 14.220 88.160 ;
        RECT 20.770 88.100 21.090 88.360 ;
        RECT 23.990 88.100 24.310 88.360 ;
        RECT 24.465 88.115 24.755 88.345 ;
        RECT 9.750 87.960 10.040 88.005 ;
        RECT 11.610 87.960 11.900 88.005 ;
        RECT 9.750 87.820 11.900 87.960 ;
        RECT 9.750 87.775 10.040 87.820 ;
        RECT 11.610 87.775 11.900 87.820 ;
        RECT 12.530 87.960 12.820 88.005 ;
        RECT 14.330 87.960 14.650 88.020 ;
        RECT 15.790 87.960 16.080 88.005 ;
        RECT 12.530 87.820 16.080 87.960 ;
        RECT 12.530 87.775 12.820 87.820 ;
        RECT 14.330 87.760 14.650 87.820 ;
        RECT 15.790 87.775 16.080 87.820 ;
        RECT 16.630 87.960 16.950 88.020 ;
        RECT 24.540 87.960 24.680 88.115 ;
        RECT 27.210 88.100 27.530 88.360 ;
        RECT 27.760 88.345 27.900 88.500 ;
        RECT 33.190 88.500 50.070 88.640 ;
        RECT 33.190 88.440 33.510 88.500 ;
        RECT 49.750 88.440 50.070 88.500 ;
        RECT 50.685 88.455 50.975 88.685 ;
        RECT 78.270 88.440 78.590 88.700 ;
        RECT 78.730 88.440 79.050 88.700 ;
        RECT 81.490 88.440 81.810 88.700 ;
        RECT 86.105 88.640 86.395 88.685 ;
        RECT 88.390 88.640 88.710 88.700 ;
        RECT 93.080 88.685 93.220 88.840 ;
        RECT 106.330 88.780 106.650 89.040 ;
        RECT 86.105 88.500 88.710 88.640 ;
        RECT 86.105 88.455 86.395 88.500 ;
        RECT 88.390 88.440 88.710 88.500 ;
        RECT 93.005 88.455 93.295 88.685 ;
        RECT 93.925 88.640 94.215 88.685 ;
        RECT 94.370 88.640 94.690 88.700 ;
        RECT 103.125 88.640 103.415 88.685 ;
        RECT 104.490 88.640 104.810 88.700 ;
        RECT 109.105 88.640 109.395 88.685 ;
        RECT 93.925 88.500 109.395 88.640 ;
        RECT 93.925 88.455 94.215 88.500 ;
        RECT 94.370 88.440 94.690 88.500 ;
        RECT 103.125 88.455 103.415 88.500 ;
        RECT 104.490 88.440 104.810 88.500 ;
        RECT 109.105 88.455 109.395 88.500 ;
        RECT 27.685 88.300 27.975 88.345 ;
        RECT 33.280 88.300 33.420 88.440 ;
        RECT 27.685 88.160 33.420 88.300 ;
        RECT 40.565 88.300 40.855 88.345 ;
        RECT 46.530 88.300 46.850 88.360 ;
        RECT 40.565 88.160 46.850 88.300 ;
        RECT 27.685 88.115 27.975 88.160 ;
        RECT 40.565 88.115 40.855 88.160 ;
        RECT 46.530 88.100 46.850 88.160 ;
        RECT 49.290 88.300 49.610 88.360 ;
        RECT 50.225 88.300 50.515 88.345 ;
        RECT 49.290 88.160 50.515 88.300 ;
        RECT 49.290 88.100 49.610 88.160 ;
        RECT 50.225 88.115 50.515 88.160 ;
        RECT 51.130 88.300 51.450 88.360 ;
        RECT 53.430 88.300 53.750 88.360 ;
        RECT 54.825 88.300 55.115 88.345 ;
        RECT 51.130 88.160 55.115 88.300 ;
        RECT 51.130 88.100 51.450 88.160 ;
        RECT 53.430 88.100 53.750 88.160 ;
        RECT 54.825 88.115 55.115 88.160 ;
        RECT 56.650 88.100 56.970 88.360 ;
        RECT 59.930 88.300 60.220 88.345 ;
        RECT 57.685 88.160 60.220 88.300 ;
        RECT 16.630 87.820 24.680 87.960 ;
        RECT 46.990 87.960 47.310 88.020 ;
        RECT 57.685 88.005 57.900 88.160 ;
        RECT 59.930 88.115 60.220 88.160 ;
        RECT 60.790 88.300 61.110 88.360 ;
        RECT 64.945 88.300 65.235 88.345 ;
        RECT 60.790 88.160 65.235 88.300 ;
        RECT 60.790 88.100 61.110 88.160 ;
        RECT 64.945 88.115 65.235 88.160 ;
        RECT 68.165 88.300 68.455 88.345 ;
        RECT 73.670 88.300 73.990 88.360 ;
        RECT 68.165 88.160 73.990 88.300 ;
        RECT 68.165 88.115 68.455 88.160 ;
        RECT 73.670 88.100 73.990 88.160 ;
        RECT 74.145 88.300 74.435 88.345 ;
        RECT 74.590 88.300 74.910 88.360 ;
        RECT 74.145 88.160 74.910 88.300 ;
        RECT 74.145 88.115 74.435 88.160 ;
        RECT 74.590 88.100 74.910 88.160 ;
        RECT 75.065 88.115 75.355 88.345 ;
        RECT 51.605 87.960 51.895 88.005 ;
        RECT 46.990 87.820 51.895 87.960 ;
        RECT 16.630 87.760 16.950 87.820 ;
        RECT 46.990 87.760 47.310 87.820 ;
        RECT 51.605 87.775 51.895 87.820 ;
        RECT 55.750 87.960 56.040 88.005 ;
        RECT 57.610 87.960 57.900 88.005 ;
        RECT 55.750 87.820 57.900 87.960 ;
        RECT 55.750 87.775 56.040 87.820 ;
        RECT 57.610 87.775 57.900 87.820 ;
        RECT 58.530 87.960 58.820 88.005 ;
        RECT 61.790 87.960 62.080 88.005 ;
        RECT 63.090 87.960 63.410 88.020 ;
        RECT 58.530 87.820 63.410 87.960 ;
        RECT 58.530 87.775 58.820 87.820 ;
        RECT 61.790 87.775 62.080 87.820 ;
        RECT 63.090 87.760 63.410 87.820 ;
        RECT 72.290 87.960 72.610 88.020 ;
        RECT 75.140 87.960 75.280 88.115 ;
        RECT 75.510 88.100 75.830 88.360 ;
        RECT 75.985 88.300 76.275 88.345 ;
        RECT 78.360 88.300 78.500 88.440 ;
        RECT 75.985 88.160 78.500 88.300 ;
        RECT 79.665 88.300 79.955 88.345 ;
        RECT 80.110 88.300 80.430 88.360 ;
        RECT 79.665 88.160 80.430 88.300 ;
        RECT 75.985 88.115 76.275 88.160 ;
        RECT 79.665 88.115 79.955 88.160 ;
        RECT 80.110 88.100 80.430 88.160 ;
        RECT 82.425 88.300 82.715 88.345 ;
        RECT 83.330 88.300 83.650 88.360 ;
        RECT 82.425 88.160 83.650 88.300 ;
        RECT 82.425 88.115 82.715 88.160 ;
        RECT 83.330 88.100 83.650 88.160 ;
        RECT 85.170 88.100 85.490 88.360 ;
        RECT 86.550 88.100 86.870 88.360 ;
        RECT 87.010 88.300 87.330 88.360 ;
        RECT 88.865 88.300 89.155 88.345 ;
        RECT 87.010 88.160 89.155 88.300 ;
        RECT 87.010 88.100 87.330 88.160 ;
        RECT 88.865 88.115 89.155 88.160 ;
        RECT 89.785 88.115 90.075 88.345 ;
        RECT 92.545 88.300 92.835 88.345 ;
        RECT 96.670 88.300 96.990 88.360 ;
        RECT 92.545 88.160 96.990 88.300 ;
        RECT 92.545 88.115 92.835 88.160 ;
        RECT 72.290 87.820 75.280 87.960 ;
        RECT 77.810 87.960 78.130 88.020 ;
        RECT 78.285 87.960 78.575 88.005 ;
        RECT 77.810 87.820 78.575 87.960 ;
        RECT 72.290 87.760 72.610 87.820 ;
        RECT 77.810 87.760 78.130 87.820 ;
        RECT 78.285 87.775 78.575 87.820 ;
        RECT 79.190 87.960 79.510 88.020 ;
        RECT 81.045 87.960 81.335 88.005 ;
        RECT 79.190 87.820 81.335 87.960 ;
        RECT 89.860 87.960 90.000 88.115 ;
        RECT 96.670 88.100 96.990 88.160 ;
        RECT 97.130 88.300 97.450 88.360 ;
        RECT 102.190 88.300 102.510 88.360 ;
        RECT 97.130 88.160 102.510 88.300 ;
        RECT 97.130 88.100 97.450 88.160 ;
        RECT 102.190 88.100 102.510 88.160 ;
        RECT 104.950 88.300 105.270 88.360 ;
        RECT 108.185 88.300 108.475 88.345 ;
        RECT 104.950 88.160 108.475 88.300 ;
        RECT 104.950 88.100 105.270 88.160 ;
        RECT 108.185 88.115 108.475 88.160 ;
        RECT 104.045 87.960 104.335 88.005 ;
        RECT 108.630 87.960 108.950 88.020 ;
        RECT 89.860 87.820 108.950 87.960 ;
        RECT 79.190 87.760 79.510 87.820 ;
        RECT 81.045 87.775 81.335 87.820 ;
        RECT 104.045 87.775 104.335 87.820 ;
        RECT 108.630 87.760 108.950 87.820 ;
        RECT 22.610 87.620 22.930 87.680 ;
        RECT 23.085 87.620 23.375 87.665 ;
        RECT 22.610 87.480 23.375 87.620 ;
        RECT 22.610 87.420 22.930 87.480 ;
        RECT 23.085 87.435 23.375 87.480 ;
        RECT 28.590 87.420 28.910 87.680 ;
        RECT 38.710 87.620 39.030 87.680 ;
        RECT 63.550 87.665 63.870 87.680 ;
        RECT 39.645 87.620 39.935 87.665 ;
        RECT 38.710 87.480 39.935 87.620 ;
        RECT 38.710 87.420 39.030 87.480 ;
        RECT 39.645 87.435 39.935 87.480 ;
        RECT 63.550 87.435 64.085 87.665 ;
        RECT 65.850 87.620 66.170 87.680 ;
        RECT 67.245 87.620 67.535 87.665 ;
        RECT 65.850 87.480 67.535 87.620 ;
        RECT 63.550 87.420 63.870 87.435 ;
        RECT 65.850 87.420 66.170 87.480 ;
        RECT 67.245 87.435 67.535 87.480 ;
        RECT 77.350 87.620 77.670 87.680 ;
        RECT 80.585 87.620 80.875 87.665 ;
        RECT 77.350 87.480 80.875 87.620 ;
        RECT 77.350 87.420 77.670 87.480 ;
        RECT 80.585 87.435 80.875 87.480 ;
        RECT 82.870 87.620 83.190 87.680 ;
        RECT 87.945 87.620 88.235 87.665 ;
        RECT 82.870 87.480 88.235 87.620 ;
        RECT 82.870 87.420 83.190 87.480 ;
        RECT 87.945 87.435 88.235 87.480 ;
        RECT 103.570 87.420 103.890 87.680 ;
        RECT 5.520 86.800 113.620 87.280 ;
        RECT 15.265 86.600 15.555 86.645 ;
        RECT 13.730 86.460 15.555 86.600 ;
        RECT 10.650 86.260 10.970 86.320 ;
        RECT 13.730 86.260 13.870 86.460 ;
        RECT 15.265 86.415 15.555 86.460 ;
        RECT 21.230 86.600 21.550 86.660 ;
        RECT 23.990 86.600 24.310 86.660 ;
        RECT 21.230 86.460 24.310 86.600 ;
        RECT 21.230 86.400 21.550 86.460 ;
        RECT 23.990 86.400 24.310 86.460 ;
        RECT 46.530 86.400 46.850 86.660 ;
        RECT 56.650 86.600 56.970 86.660 ;
        RECT 57.585 86.600 57.875 86.645 ;
        RECT 56.650 86.460 57.875 86.600 ;
        RECT 56.650 86.400 56.970 86.460 ;
        RECT 57.585 86.415 57.875 86.460 ;
        RECT 58.965 86.415 59.255 86.645 ;
        RECT 61.265 86.600 61.555 86.645 ;
        RECT 62.630 86.600 62.950 86.660 ;
        RECT 63.550 86.600 63.870 86.660 ;
        RECT 61.265 86.460 63.870 86.600 ;
        RECT 61.265 86.415 61.555 86.460 ;
        RECT 10.650 86.120 13.870 86.260 ;
        RECT 10.650 86.060 10.970 86.120 ;
        RECT 14.330 86.060 14.650 86.320 ;
        RECT 19.390 86.260 19.710 86.320 ;
        RECT 37.810 86.260 38.100 86.305 ;
        RECT 39.670 86.260 39.960 86.305 ;
        RECT 19.390 86.120 22.840 86.260 ;
        RECT 19.390 86.060 19.710 86.120 ;
        RECT 14.790 85.720 15.110 85.980 ;
        RECT 16.185 85.920 16.475 85.965 ;
        RECT 17.550 85.920 17.870 85.980 ;
        RECT 16.185 85.780 17.870 85.920 ;
        RECT 16.185 85.735 16.475 85.780 ;
        RECT 17.550 85.720 17.870 85.780 ;
        RECT 21.230 85.920 21.550 85.980 ;
        RECT 22.700 85.965 22.840 86.120 ;
        RECT 37.810 86.120 39.960 86.260 ;
        RECT 37.810 86.075 38.100 86.120 ;
        RECT 39.670 86.075 39.960 86.120 ;
        RECT 40.590 86.260 40.880 86.305 ;
        RECT 42.390 86.260 42.710 86.320 ;
        RECT 43.850 86.260 44.140 86.305 ;
        RECT 40.590 86.120 44.140 86.260 ;
        RECT 40.590 86.075 40.880 86.120 ;
        RECT 21.705 85.920 21.995 85.965 ;
        RECT 21.230 85.780 21.995 85.920 ;
        RECT 21.230 85.720 21.550 85.780 ;
        RECT 21.705 85.735 21.995 85.780 ;
        RECT 22.625 85.735 22.915 85.965 ;
        RECT 23.990 85.720 24.310 85.980 ;
        RECT 32.270 85.720 32.590 85.980 ;
        RECT 35.505 85.920 35.795 85.965 ;
        RECT 37.330 85.920 37.650 85.980 ;
        RECT 35.505 85.780 37.650 85.920 ;
        RECT 35.505 85.735 35.795 85.780 ;
        RECT 20.770 85.580 21.090 85.640 ;
        RECT 23.085 85.580 23.375 85.625 ;
        RECT 20.770 85.440 23.375 85.580 ;
        RECT 20.770 85.380 21.090 85.440 ;
        RECT 23.085 85.395 23.375 85.440 ;
        RECT 29.970 85.580 30.290 85.640 ;
        RECT 35.580 85.580 35.720 85.735 ;
        RECT 37.330 85.720 37.650 85.780 ;
        RECT 38.710 85.720 39.030 85.980 ;
        RECT 39.745 85.920 39.960 86.075 ;
        RECT 42.390 86.060 42.710 86.120 ;
        RECT 43.850 86.075 44.140 86.120 ;
        RECT 53.905 86.260 54.195 86.305 ;
        RECT 54.365 86.260 54.655 86.305 ;
        RECT 53.905 86.120 54.655 86.260 ;
        RECT 53.905 86.075 54.195 86.120 ;
        RECT 54.365 86.075 54.655 86.120 ;
        RECT 41.990 85.920 42.280 85.965 ;
        RECT 39.745 85.780 42.280 85.920 ;
        RECT 41.990 85.735 42.280 85.780 ;
        RECT 47.910 85.920 48.230 85.980 ;
        RECT 48.385 85.920 48.675 85.965 ;
        RECT 47.910 85.780 48.675 85.920 ;
        RECT 47.910 85.720 48.230 85.780 ;
        RECT 48.385 85.735 48.675 85.780 ;
        RECT 48.845 85.920 49.135 85.965 ;
        RECT 50.210 85.920 50.530 85.980 ;
        RECT 50.685 85.920 50.975 85.965 ;
        RECT 48.845 85.780 49.980 85.920 ;
        RECT 48.845 85.735 49.135 85.780 ;
        RECT 29.970 85.440 35.720 85.580 ;
        RECT 29.970 85.380 30.290 85.440 ;
        RECT 36.870 85.380 37.190 85.640 ;
        RECT 47.450 85.580 47.770 85.640 ;
        RECT 49.305 85.580 49.595 85.625 ;
        RECT 47.450 85.440 49.595 85.580 ;
        RECT 47.450 85.380 47.770 85.440 ;
        RECT 49.305 85.395 49.595 85.440 ;
        RECT 49.840 85.580 49.980 85.780 ;
        RECT 50.210 85.780 50.975 85.920 ;
        RECT 50.210 85.720 50.530 85.780 ;
        RECT 50.685 85.735 50.975 85.780 ;
        RECT 51.605 85.735 51.895 85.965 ;
        RECT 51.680 85.580 51.820 85.735 ;
        RECT 52.050 85.720 52.370 85.980 ;
        RECT 52.525 85.920 52.815 85.965 ;
        RECT 52.970 85.920 53.290 85.980 ;
        RECT 52.525 85.780 53.290 85.920 ;
        RECT 52.525 85.735 52.815 85.780 ;
        RECT 52.970 85.720 53.290 85.780 ;
        RECT 53.430 85.920 53.750 85.980 ;
        RECT 55.745 85.920 56.035 85.965 ;
        RECT 53.430 85.780 56.035 85.920 ;
        RECT 53.430 85.720 53.750 85.780 ;
        RECT 55.745 85.735 56.035 85.780 ;
        RECT 58.505 85.920 58.795 85.965 ;
        RECT 59.040 85.920 59.180 86.415 ;
        RECT 62.630 86.400 62.950 86.460 ;
        RECT 63.550 86.400 63.870 86.460 ;
        RECT 73.670 86.400 73.990 86.660 ;
        RECT 75.510 86.600 75.830 86.660 ;
        RECT 75.510 86.460 77.580 86.600 ;
        RECT 75.510 86.400 75.830 86.460 ;
        RECT 60.805 86.260 61.095 86.305 ;
        RECT 63.090 86.260 63.410 86.320 ;
        RECT 60.805 86.120 63.410 86.260 ;
        RECT 60.805 86.075 61.095 86.120 ;
        RECT 63.090 86.060 63.410 86.120 ;
        RECT 64.010 86.060 64.330 86.320 ;
        RECT 64.950 86.260 65.240 86.305 ;
        RECT 66.810 86.260 67.100 86.305 ;
        RECT 64.950 86.120 67.100 86.260 ;
        RECT 64.950 86.075 65.240 86.120 ;
        RECT 66.810 86.075 67.100 86.120 ;
        RECT 67.730 86.260 68.020 86.305 ;
        RECT 70.990 86.260 71.280 86.305 ;
        RECT 71.830 86.260 72.150 86.320 ;
        RECT 67.730 86.120 72.150 86.260 ;
        RECT 67.730 86.075 68.020 86.120 ;
        RECT 70.990 86.075 71.280 86.120 ;
        RECT 64.100 85.920 64.240 86.060 ;
        RECT 58.505 85.780 59.180 85.920 ;
        RECT 62.260 85.780 65.620 85.920 ;
        RECT 58.505 85.735 58.795 85.780 ;
        RECT 49.840 85.440 51.820 85.580 ;
        RECT 37.350 85.240 37.640 85.285 ;
        RECT 39.210 85.240 39.500 85.285 ;
        RECT 41.990 85.240 42.280 85.285 ;
        RECT 37.350 85.100 42.280 85.240 ;
        RECT 37.350 85.055 37.640 85.100 ;
        RECT 39.210 85.055 39.500 85.100 ;
        RECT 41.990 85.055 42.280 85.100 ;
        RECT 20.785 84.900 21.075 84.945 ;
        RECT 21.230 84.900 21.550 84.960 ;
        RECT 20.785 84.760 21.550 84.900 ;
        RECT 20.785 84.715 21.075 84.760 ;
        RECT 21.230 84.700 21.550 84.760 ;
        RECT 24.925 84.900 25.215 84.945 ;
        RECT 28.130 84.900 28.450 84.960 ;
        RECT 24.925 84.760 28.450 84.900 ;
        RECT 24.925 84.715 25.215 84.760 ;
        RECT 28.130 84.700 28.450 84.760 ;
        RECT 32.730 84.900 33.050 84.960 ;
        RECT 33.205 84.900 33.495 84.945 ;
        RECT 32.730 84.760 33.495 84.900 ;
        RECT 32.730 84.700 33.050 84.760 ;
        RECT 33.205 84.715 33.495 84.760 ;
        RECT 35.490 84.900 35.810 84.960 ;
        RECT 35.965 84.900 36.255 84.945 ;
        RECT 35.490 84.760 36.255 84.900 ;
        RECT 35.490 84.700 35.810 84.760 ;
        RECT 35.965 84.715 36.255 84.760 ;
        RECT 44.690 84.900 45.010 84.960 ;
        RECT 45.855 84.900 46.145 84.945 ;
        RECT 49.840 84.900 49.980 85.440 ;
        RECT 55.270 85.380 55.590 85.640 ;
        RECT 62.260 85.625 62.400 85.780 ;
        RECT 62.185 85.395 62.475 85.625 ;
        RECT 63.550 85.580 63.870 85.640 ;
        RECT 64.025 85.580 64.315 85.625 ;
        RECT 63.550 85.440 64.315 85.580 ;
        RECT 65.480 85.580 65.620 85.780 ;
        RECT 65.850 85.720 66.170 85.980 ;
        RECT 66.885 85.920 67.100 86.075 ;
        RECT 71.830 86.060 72.150 86.120 ;
        RECT 72.290 86.260 72.610 86.320 ;
        RECT 72.995 86.260 73.285 86.305 ;
        RECT 75.985 86.260 76.275 86.305 ;
        RECT 72.290 86.120 76.275 86.260 ;
        RECT 77.440 86.260 77.580 86.460 ;
        RECT 77.810 86.400 78.130 86.660 ;
        RECT 78.270 86.600 78.590 86.660 ;
        RECT 79.190 86.600 79.510 86.660 ;
        RECT 78.270 86.460 79.510 86.600 ;
        RECT 78.270 86.400 78.590 86.460 ;
        RECT 79.190 86.400 79.510 86.460 ;
        RECT 80.570 86.260 80.890 86.320 ;
        RECT 77.440 86.120 80.890 86.260 ;
        RECT 72.290 86.060 72.610 86.120 ;
        RECT 72.995 86.075 73.285 86.120 ;
        RECT 75.985 86.075 76.275 86.120 ;
        RECT 69.130 85.920 69.420 85.965 ;
        RECT 66.885 85.780 69.420 85.920 ;
        RECT 69.130 85.735 69.420 85.780 ;
        RECT 75.525 85.920 75.815 85.965 ;
        RECT 77.350 85.920 77.670 85.980 ;
        RECT 75.525 85.780 78.960 85.920 ;
        RECT 75.525 85.735 75.815 85.780 ;
        RECT 77.350 85.720 77.670 85.780 ;
        RECT 73.210 85.580 73.530 85.640 ;
        RECT 76.445 85.580 76.735 85.625 ;
        RECT 77.810 85.580 78.130 85.640 ;
        RECT 65.480 85.440 78.130 85.580 ;
        RECT 78.820 85.580 78.960 85.780 ;
        RECT 79.190 85.720 79.510 85.980 ;
        RECT 79.740 85.965 79.880 86.120 ;
        RECT 80.570 86.060 80.890 86.120 ;
        RECT 79.665 85.735 79.955 85.965 ;
        RECT 80.125 85.735 80.415 85.965 ;
        RECT 81.045 85.920 81.335 85.965 ;
        RECT 82.410 85.920 82.730 85.980 ;
        RECT 81.045 85.780 82.730 85.920 ;
        RECT 81.045 85.735 81.335 85.780 ;
        RECT 80.200 85.580 80.340 85.735 ;
        RECT 82.410 85.720 82.730 85.780 ;
        RECT 78.820 85.440 80.340 85.580 ;
        RECT 63.550 85.380 63.870 85.440 ;
        RECT 64.025 85.395 64.315 85.440 ;
        RECT 73.210 85.380 73.530 85.440 ;
        RECT 76.445 85.395 76.735 85.440 ;
        RECT 77.810 85.380 78.130 85.440 ;
        RECT 56.665 85.240 56.955 85.285 ;
        RECT 57.110 85.240 57.430 85.300 ;
        RECT 56.665 85.100 57.430 85.240 ;
        RECT 56.665 85.055 56.955 85.100 ;
        RECT 57.110 85.040 57.430 85.100 ;
        RECT 64.490 85.240 64.780 85.285 ;
        RECT 66.350 85.240 66.640 85.285 ;
        RECT 69.130 85.240 69.420 85.285 ;
        RECT 64.490 85.100 69.420 85.240 ;
        RECT 64.490 85.055 64.780 85.100 ;
        RECT 66.350 85.055 66.640 85.100 ;
        RECT 69.130 85.055 69.420 85.100 ;
        RECT 44.690 84.760 49.980 84.900 ;
        RECT 53.890 84.900 54.210 84.960 ;
        RECT 54.365 84.900 54.655 84.945 ;
        RECT 53.890 84.760 54.655 84.900 ;
        RECT 44.690 84.700 45.010 84.760 ;
        RECT 45.855 84.715 46.145 84.760 ;
        RECT 53.890 84.700 54.210 84.760 ;
        RECT 54.365 84.715 54.655 84.760 ;
        RECT 72.750 84.900 73.070 84.960 ;
        RECT 90.230 84.900 90.550 84.960 ;
        RECT 93.910 84.900 94.230 84.960 ;
        RECT 72.750 84.760 94.230 84.900 ;
        RECT 72.750 84.700 73.070 84.760 ;
        RECT 90.230 84.700 90.550 84.760 ;
        RECT 93.910 84.700 94.230 84.760 ;
        RECT 5.520 84.080 113.620 84.560 ;
        RECT 14.790 83.880 15.110 83.940 ;
        RECT 29.970 83.880 30.290 83.940 ;
        RECT 14.790 83.740 30.290 83.880 ;
        RECT 14.790 83.680 15.110 83.740 ;
        RECT 29.970 83.680 30.290 83.740 ;
        RECT 34.570 83.880 34.890 83.940 ;
        RECT 39.875 83.880 40.165 83.925 ;
        RECT 34.570 83.740 41.470 83.880 ;
        RECT 34.570 83.680 34.890 83.740 ;
        RECT 39.875 83.695 40.165 83.740 ;
        RECT 21.710 83.540 22.000 83.585 ;
        RECT 23.570 83.540 23.860 83.585 ;
        RECT 26.350 83.540 26.640 83.585 ;
        RECT 21.710 83.400 26.640 83.540 ;
        RECT 21.710 83.355 22.000 83.400 ;
        RECT 23.570 83.355 23.860 83.400 ;
        RECT 26.350 83.355 26.640 83.400 ;
        RECT 31.370 83.540 31.660 83.585 ;
        RECT 33.230 83.540 33.520 83.585 ;
        RECT 36.010 83.540 36.300 83.585 ;
        RECT 31.370 83.400 36.300 83.540 ;
        RECT 41.330 83.540 41.470 83.740 ;
        RECT 46.990 83.680 47.310 83.940 ;
        RECT 55.270 83.880 55.590 83.940 ;
        RECT 57.570 83.880 57.890 83.940 ;
        RECT 55.270 83.740 57.890 83.880 ;
        RECT 55.270 83.680 55.590 83.740 ;
        RECT 57.570 83.680 57.890 83.740 ;
        RECT 70.925 83.880 71.215 83.925 ;
        RECT 71.830 83.880 72.150 83.940 ;
        RECT 70.925 83.740 72.150 83.880 ;
        RECT 70.925 83.695 71.215 83.740 ;
        RECT 71.830 83.680 72.150 83.740 ;
        RECT 77.350 83.880 77.670 83.940 ;
        RECT 82.655 83.880 82.945 83.925 ;
        RECT 103.570 83.880 103.890 83.940 ;
        RECT 105.870 83.880 106.190 83.940 ;
        RECT 111.175 83.880 111.465 83.925 ;
        RECT 77.350 83.740 82.945 83.880 ;
        RECT 77.350 83.680 77.670 83.740 ;
        RECT 82.655 83.695 82.945 83.740 ;
        RECT 93.080 83.740 111.465 83.880 ;
        RECT 47.910 83.540 48.230 83.600 ;
        RECT 49.750 83.540 50.070 83.600 ;
        RECT 59.885 83.540 60.175 83.585 ;
        RECT 72.750 83.540 73.070 83.600 ;
        RECT 41.330 83.400 48.370 83.540 ;
        RECT 31.370 83.355 31.660 83.400 ;
        RECT 33.230 83.355 33.520 83.400 ;
        RECT 36.010 83.355 36.300 83.400 ;
        RECT 47.910 83.340 48.370 83.400 ;
        RECT 49.750 83.400 73.070 83.540 ;
        RECT 49.750 83.340 50.070 83.400 ;
        RECT 59.885 83.355 60.175 83.400 ;
        RECT 72.750 83.340 73.070 83.400 ;
        RECT 74.150 83.540 74.440 83.585 ;
        RECT 76.010 83.540 76.300 83.585 ;
        RECT 78.790 83.540 79.080 83.585 ;
        RECT 74.150 83.400 79.080 83.540 ;
        RECT 74.150 83.355 74.440 83.400 ;
        RECT 76.010 83.355 76.300 83.400 ;
        RECT 78.790 83.355 79.080 83.400 ;
        RECT 21.245 83.200 21.535 83.245 ;
        RECT 22.150 83.200 22.470 83.260 ;
        RECT 30.905 83.200 31.195 83.245 ;
        RECT 21.245 83.060 31.195 83.200 ;
        RECT 21.245 83.015 21.535 83.060 ;
        RECT 22.150 83.000 22.470 83.060 ;
        RECT 30.905 83.015 31.195 83.060 ;
        RECT 32.730 83.000 33.050 83.260 ;
        RECT 36.870 83.200 37.190 83.260 ;
        RECT 46.990 83.200 47.310 83.260 ;
        RECT 36.870 83.060 47.310 83.200 ;
        RECT 48.230 83.200 48.370 83.340 ;
        RECT 63.550 83.200 63.870 83.260 ;
        RECT 73.685 83.200 73.975 83.245 ;
        RECT 76.890 83.200 77.210 83.260 ;
        RECT 93.080 83.245 93.220 83.740 ;
        RECT 103.570 83.680 103.890 83.740 ;
        RECT 105.870 83.680 106.190 83.740 ;
        RECT 111.175 83.695 111.465 83.740 ;
        RECT 97.130 83.540 97.450 83.600 ;
        RECT 102.670 83.540 102.960 83.585 ;
        RECT 104.530 83.540 104.820 83.585 ;
        RECT 107.310 83.540 107.600 83.585 ;
        RECT 97.130 83.340 97.590 83.540 ;
        RECT 102.670 83.400 107.600 83.540 ;
        RECT 102.670 83.355 102.960 83.400 ;
        RECT 104.530 83.355 104.820 83.400 ;
        RECT 107.310 83.355 107.600 83.400 ;
        RECT 48.230 83.060 49.520 83.200 ;
        RECT 36.870 83.000 37.190 83.060 ;
        RECT 46.990 83.000 47.310 83.060 ;
        RECT 23.070 82.660 23.390 82.920 ;
        RECT 26.350 82.860 26.640 82.905 ;
        RECT 36.010 82.860 36.300 82.905 ;
        RECT 24.105 82.720 26.640 82.860 ;
        RECT 24.105 82.565 24.320 82.720 ;
        RECT 26.350 82.675 26.640 82.720 ;
        RECT 33.765 82.720 36.300 82.860 ;
        RECT 22.170 82.520 22.460 82.565 ;
        RECT 24.030 82.520 24.320 82.565 ;
        RECT 22.170 82.380 24.320 82.520 ;
        RECT 22.170 82.335 22.460 82.380 ;
        RECT 24.030 82.335 24.320 82.380 ;
        RECT 24.950 82.520 25.240 82.565 ;
        RECT 28.210 82.520 28.500 82.565 ;
        RECT 29.050 82.520 29.370 82.580 ;
        RECT 33.765 82.565 33.980 82.720 ;
        RECT 36.010 82.675 36.300 82.720 ;
        RECT 37.330 82.860 37.650 82.920 ;
        RECT 41.025 82.860 41.315 82.905 ;
        RECT 37.330 82.720 41.315 82.860 ;
        RECT 37.330 82.660 37.650 82.720 ;
        RECT 41.025 82.675 41.315 82.720 ;
        RECT 41.485 82.860 41.775 82.905 ;
        RECT 42.390 82.860 42.710 82.920 ;
        RECT 49.380 82.905 49.520 83.060 ;
        RECT 63.550 83.060 77.210 83.200 ;
        RECT 63.550 83.000 63.870 83.060 ;
        RECT 73.685 83.015 73.975 83.060 ;
        RECT 76.890 83.000 77.210 83.060 ;
        RECT 93.005 83.015 93.295 83.245 ;
        RECT 94.830 83.000 95.150 83.260 ;
        RECT 41.485 82.720 42.710 82.860 ;
        RECT 41.485 82.675 41.775 82.720 ;
        RECT 24.950 82.380 29.370 82.520 ;
        RECT 24.950 82.335 25.240 82.380 ;
        RECT 28.210 82.335 28.500 82.380 ;
        RECT 29.050 82.320 29.370 82.380 ;
        RECT 31.830 82.520 32.120 82.565 ;
        RECT 33.690 82.520 33.980 82.565 ;
        RECT 31.830 82.380 33.980 82.520 ;
        RECT 31.830 82.335 32.120 82.380 ;
        RECT 33.690 82.335 33.980 82.380 ;
        RECT 34.610 82.520 34.900 82.565 ;
        RECT 35.490 82.520 35.810 82.580 ;
        RECT 37.870 82.520 38.160 82.565 ;
        RECT 34.610 82.380 38.160 82.520 ;
        RECT 41.100 82.520 41.240 82.675 ;
        RECT 42.390 82.660 42.710 82.720 ;
        RECT 48.385 82.675 48.675 82.905 ;
        RECT 48.845 82.675 49.135 82.905 ;
        RECT 49.305 82.675 49.595 82.905 ;
        RECT 41.930 82.520 42.250 82.580 ;
        RECT 41.100 82.380 42.250 82.520 ;
        RECT 34.610 82.335 34.900 82.380 ;
        RECT 35.490 82.320 35.810 82.380 ;
        RECT 37.870 82.335 38.160 82.380 ;
        RECT 41.930 82.320 42.250 82.380 ;
        RECT 27.670 82.180 27.990 82.240 ;
        RECT 30.215 82.180 30.505 82.225 ;
        RECT 34.110 82.180 34.430 82.240 ;
        RECT 27.670 82.040 34.430 82.180 ;
        RECT 48.460 82.180 48.600 82.675 ;
        RECT 48.920 82.520 49.060 82.675 ;
        RECT 50.210 82.660 50.530 82.920 ;
        RECT 67.230 82.860 67.550 82.920 ;
        RECT 69.070 82.860 69.390 82.920 ;
        RECT 71.370 82.860 71.690 82.920 ;
        RECT 67.230 82.720 71.690 82.860 ;
        RECT 67.230 82.660 67.550 82.720 ;
        RECT 69.070 82.660 69.390 82.720 ;
        RECT 71.370 82.660 71.690 82.720 ;
        RECT 72.290 82.660 72.610 82.920 ;
        RECT 75.525 82.860 75.815 82.905 ;
        RECT 78.790 82.860 79.080 82.905 ;
        RECT 73.300 82.720 75.815 82.860 ;
        RECT 52.050 82.520 52.370 82.580 ;
        RECT 48.920 82.380 52.370 82.520 ;
        RECT 52.050 82.320 52.370 82.380 ;
        RECT 59.870 82.520 60.190 82.580 ;
        RECT 60.790 82.520 61.110 82.580 ;
        RECT 59.870 82.380 61.110 82.520 ;
        RECT 59.870 82.320 60.190 82.380 ;
        RECT 60.790 82.320 61.110 82.380 ;
        RECT 52.970 82.180 53.290 82.240 ;
        RECT 73.300 82.225 73.440 82.720 ;
        RECT 75.525 82.675 75.815 82.720 ;
        RECT 76.545 82.720 79.080 82.860 ;
        RECT 76.545 82.565 76.760 82.720 ;
        RECT 78.790 82.675 79.080 82.720 ;
        RECT 93.910 82.660 94.230 82.920 ;
        RECT 97.450 82.905 97.590 83.340 ;
        RECT 98.050 83.200 98.370 83.260 ;
        RECT 102.205 83.200 102.495 83.245 ;
        RECT 98.050 83.060 102.495 83.200 ;
        RECT 98.050 83.000 98.370 83.060 ;
        RECT 102.205 83.015 102.495 83.060 ;
        RECT 104.045 83.200 104.335 83.245 ;
        RECT 106.330 83.200 106.650 83.260 ;
        RECT 104.045 83.060 106.650 83.200 ;
        RECT 104.045 83.015 104.335 83.060 ;
        RECT 106.330 83.000 106.650 83.060 ;
        RECT 97.185 82.720 97.590 82.905 ;
        RECT 107.310 82.860 107.600 82.905 ;
        RECT 105.065 82.720 107.600 82.860 ;
        RECT 97.185 82.675 97.475 82.720 ;
        RECT 74.610 82.520 74.900 82.565 ;
        RECT 76.470 82.520 76.760 82.565 ;
        RECT 74.610 82.380 76.760 82.520 ;
        RECT 74.610 82.335 74.900 82.380 ;
        RECT 76.470 82.335 76.760 82.380 ;
        RECT 77.390 82.520 77.680 82.565 ;
        RECT 79.650 82.520 79.970 82.580 ;
        RECT 105.065 82.565 105.280 82.720 ;
        RECT 107.310 82.675 107.600 82.720 ;
        RECT 80.650 82.520 80.940 82.565 ;
        RECT 77.390 82.380 80.940 82.520 ;
        RECT 77.390 82.335 77.680 82.380 ;
        RECT 79.650 82.320 79.970 82.380 ;
        RECT 80.650 82.335 80.940 82.380 ;
        RECT 103.130 82.520 103.420 82.565 ;
        RECT 104.990 82.520 105.280 82.565 ;
        RECT 103.130 82.380 105.280 82.520 ;
        RECT 103.130 82.335 103.420 82.380 ;
        RECT 104.990 82.335 105.280 82.380 ;
        RECT 105.910 82.520 106.200 82.565 ;
        RECT 109.170 82.520 109.460 82.565 ;
        RECT 110.930 82.520 111.250 82.580 ;
        RECT 105.910 82.380 111.250 82.520 ;
        RECT 105.910 82.335 106.200 82.380 ;
        RECT 109.170 82.335 109.460 82.380 ;
        RECT 110.930 82.320 111.250 82.380 ;
        RECT 48.460 82.040 53.290 82.180 ;
        RECT 27.670 81.980 27.990 82.040 ;
        RECT 30.215 81.995 30.505 82.040 ;
        RECT 34.110 81.980 34.430 82.040 ;
        RECT 52.970 81.980 53.290 82.040 ;
        RECT 73.225 81.995 73.515 82.225 ;
        RECT 96.670 81.980 96.990 82.240 ;
        RECT 5.520 81.360 113.620 81.840 ;
        RECT 23.070 80.960 23.390 81.220 ;
        RECT 24.465 80.975 24.755 81.205 ;
        RECT 26.765 81.160 27.055 81.205 ;
        RECT 27.670 81.160 27.990 81.220 ;
        RECT 26.765 81.020 27.990 81.160 ;
        RECT 26.765 80.975 27.055 81.020 ;
        RECT 16.630 80.820 16.950 80.880 ;
        RECT 11.200 80.680 16.950 80.820 ;
        RECT 11.200 80.525 11.340 80.680 ;
        RECT 16.630 80.620 16.950 80.680 ;
        RECT 11.125 80.295 11.415 80.525 ;
        RECT 12.505 80.480 12.795 80.525 ;
        RECT 16.185 80.480 16.475 80.525 ;
        RECT 18.930 80.480 19.250 80.540 ;
        RECT 12.505 80.340 13.870 80.480 ;
        RECT 12.505 80.295 12.795 80.340 ;
        RECT 13.730 79.800 13.870 80.340 ;
        RECT 16.185 80.340 19.250 80.480 ;
        RECT 16.185 80.295 16.475 80.340 ;
        RECT 18.930 80.280 19.250 80.340 ;
        RECT 24.005 80.480 24.295 80.525 ;
        RECT 24.540 80.480 24.680 80.975 ;
        RECT 27.670 80.960 27.990 81.020 ;
        RECT 29.050 80.960 29.370 81.220 ;
        RECT 32.270 80.960 32.590 81.220 ;
        RECT 34.570 80.960 34.890 81.220 ;
        RECT 44.690 80.960 45.010 81.220 ;
        RECT 72.290 81.160 72.610 81.220 ;
        RECT 75.065 81.160 75.355 81.205 ;
        RECT 72.290 81.020 75.355 81.160 ;
        RECT 72.290 80.960 72.610 81.020 ;
        RECT 75.065 80.975 75.355 81.020 ;
        RECT 77.350 80.960 77.670 81.220 ;
        RECT 79.650 80.960 79.970 81.220 ;
        RECT 92.990 81.160 93.310 81.220 ;
        RECT 97.590 81.160 97.910 81.220 ;
        RECT 92.990 81.020 97.910 81.160 ;
        RECT 92.990 80.960 93.310 81.020 ;
        RECT 97.590 80.960 97.910 81.020 ;
        RECT 104.505 80.975 104.795 81.205 ;
        RECT 71.370 80.820 71.690 80.880 ;
        RECT 92.090 80.820 92.380 80.865 ;
        RECT 93.950 80.820 94.240 80.865 ;
        RECT 35.580 80.680 46.300 80.820 ;
        RECT 24.005 80.340 24.680 80.480 ;
        RECT 24.005 80.295 24.295 80.340 ;
        RECT 26.305 80.295 26.595 80.525 ;
        RECT 29.525 80.480 29.815 80.525 ;
        RECT 29.970 80.480 30.290 80.540 ;
        RECT 29.525 80.340 30.290 80.480 ;
        RECT 29.525 80.295 29.815 80.340 ;
        RECT 16.645 79.955 16.935 80.185 ;
        RECT 17.565 80.140 17.855 80.185 ;
        RECT 19.850 80.140 20.170 80.200 ;
        RECT 17.565 80.000 20.170 80.140 ;
        RECT 17.565 79.955 17.855 80.000 ;
        RECT 14.345 79.800 14.635 79.845 ;
        RECT 13.730 79.660 14.635 79.800 ;
        RECT 16.720 79.800 16.860 79.955 ;
        RECT 19.850 79.940 20.170 80.000 ;
        RECT 23.070 80.140 23.390 80.200 ;
        RECT 26.380 80.140 26.520 80.295 ;
        RECT 29.970 80.280 30.290 80.340 ;
        RECT 34.110 80.280 34.430 80.540 ;
        RECT 35.580 80.185 35.720 80.680 ;
        RECT 41.945 80.480 42.235 80.525 ;
        RECT 41.945 80.340 43.080 80.480 ;
        RECT 41.945 80.295 42.235 80.340 ;
        RECT 23.070 80.000 26.520 80.140 ;
        RECT 27.685 80.140 27.975 80.185 ;
        RECT 35.505 80.140 35.795 80.185 ;
        RECT 27.685 80.000 35.795 80.140 ;
        RECT 23.070 79.940 23.390 80.000 ;
        RECT 27.685 79.955 27.975 80.000 ;
        RECT 35.505 79.955 35.795 80.000 ;
        RECT 23.160 79.800 23.300 79.940 ;
        RECT 16.720 79.660 23.300 79.800 ;
        RECT 14.345 79.615 14.635 79.660 ;
        RECT 7.890 79.460 8.210 79.520 ;
        RECT 10.205 79.460 10.495 79.505 ;
        RECT 7.890 79.320 10.495 79.460 ;
        RECT 7.890 79.260 8.210 79.320 ;
        RECT 10.205 79.275 10.495 79.320 ;
        RECT 11.570 79.260 11.890 79.520 ;
        RECT 19.850 79.460 20.170 79.520 ;
        RECT 27.760 79.460 27.900 79.955 ;
        RECT 42.940 79.845 43.080 80.340 ;
        RECT 45.150 79.940 45.470 80.200 ;
        RECT 46.160 80.185 46.300 80.680 ;
        RECT 71.370 80.680 80.340 80.820 ;
        RECT 71.370 80.620 71.690 80.680 ;
        RECT 76.905 80.480 77.195 80.525 ;
        RECT 77.350 80.480 77.670 80.540 ;
        RECT 80.200 80.525 80.340 80.680 ;
        RECT 92.090 80.680 94.240 80.820 ;
        RECT 92.090 80.635 92.380 80.680 ;
        RECT 93.950 80.635 94.240 80.680 ;
        RECT 94.870 80.820 95.160 80.865 ;
        RECT 96.670 80.820 96.990 80.880 ;
        RECT 98.130 80.820 98.420 80.865 ;
        RECT 94.870 80.680 98.420 80.820 ;
        RECT 94.870 80.635 95.160 80.680 ;
        RECT 76.905 80.340 77.670 80.480 ;
        RECT 76.905 80.295 77.195 80.340 ;
        RECT 77.350 80.280 77.670 80.340 ;
        RECT 80.125 80.480 80.415 80.525 ;
        RECT 84.250 80.480 84.570 80.540 ;
        RECT 80.125 80.340 84.570 80.480 ;
        RECT 80.125 80.295 80.415 80.340 ;
        RECT 84.250 80.280 84.570 80.340 ;
        RECT 89.770 80.280 90.090 80.540 ;
        RECT 91.165 80.480 91.455 80.525 ;
        RECT 94.025 80.480 94.240 80.635 ;
        RECT 96.670 80.620 96.990 80.680 ;
        RECT 98.130 80.635 98.420 80.680 ;
        RECT 96.270 80.480 96.560 80.525 ;
        RECT 91.165 80.340 93.680 80.480 ;
        RECT 94.025 80.340 96.560 80.480 ;
        RECT 91.165 80.295 91.455 80.340 ;
        RECT 46.085 80.140 46.375 80.185 ;
        RECT 47.450 80.140 47.770 80.200 ;
        RECT 46.085 80.000 47.770 80.140 ;
        RECT 46.085 79.955 46.375 80.000 ;
        RECT 47.450 79.940 47.770 80.000 ;
        RECT 77.810 79.940 78.130 80.200 ;
        RECT 93.005 80.140 93.295 80.185 ;
        RECT 90.780 80.000 93.295 80.140 ;
        RECT 93.540 80.140 93.680 80.340 ;
        RECT 96.270 80.295 96.560 80.340 ;
        RECT 102.665 80.480 102.955 80.525 ;
        RECT 103.570 80.480 103.890 80.540 ;
        RECT 102.665 80.340 103.890 80.480 ;
        RECT 104.580 80.480 104.720 80.975 ;
        RECT 106.330 80.960 106.650 81.220 ;
        RECT 110.930 80.960 111.250 81.220 ;
        RECT 105.885 80.480 106.175 80.525 ;
        RECT 104.580 80.340 106.175 80.480 ;
        RECT 102.665 80.295 102.955 80.340 ;
        RECT 103.570 80.280 103.890 80.340 ;
        RECT 105.885 80.295 106.175 80.340 ;
        RECT 107.250 80.280 107.570 80.540 ;
        RECT 110.025 80.480 110.315 80.525 ;
        RECT 110.470 80.480 110.790 80.540 ;
        RECT 110.025 80.340 110.790 80.480 ;
        RECT 110.025 80.295 110.315 80.340 ;
        RECT 110.470 80.280 110.790 80.340 ;
        RECT 98.050 80.140 98.370 80.200 ;
        RECT 93.540 80.000 98.370 80.140 ;
        RECT 90.780 79.845 90.920 80.000 ;
        RECT 93.005 79.955 93.295 80.000 ;
        RECT 98.050 79.940 98.370 80.000 ;
        RECT 101.730 79.940 102.050 80.200 ;
        RECT 102.205 79.955 102.495 80.185 ;
        RECT 42.865 79.615 43.155 79.845 ;
        RECT 90.705 79.615 90.995 79.845 ;
        RECT 91.630 79.800 91.920 79.845 ;
        RECT 93.490 79.800 93.780 79.845 ;
        RECT 96.270 79.800 96.560 79.845 ;
        RECT 91.630 79.660 96.560 79.800 ;
        RECT 91.630 79.615 91.920 79.660 ;
        RECT 93.490 79.615 93.780 79.660 ;
        RECT 96.270 79.615 96.560 79.660 ;
        RECT 19.850 79.320 27.900 79.460 ;
        RECT 39.170 79.460 39.490 79.520 ;
        RECT 41.025 79.460 41.315 79.505 ;
        RECT 39.170 79.320 41.315 79.460 ;
        RECT 19.850 79.260 20.170 79.320 ;
        RECT 39.170 79.260 39.490 79.320 ;
        RECT 41.025 79.275 41.315 79.320 ;
        RECT 97.590 79.460 97.910 79.520 ;
        RECT 100.135 79.460 100.425 79.505 ;
        RECT 102.280 79.460 102.420 79.955 ;
        RECT 97.590 79.320 102.420 79.460 ;
        RECT 102.650 79.460 102.970 79.520 ;
        RECT 104.965 79.460 105.255 79.505 ;
        RECT 102.650 79.320 105.255 79.460 ;
        RECT 97.590 79.260 97.910 79.320 ;
        RECT 100.135 79.275 100.425 79.320 ;
        RECT 102.650 79.260 102.970 79.320 ;
        RECT 104.965 79.275 105.255 79.320 ;
        RECT 107.710 79.460 108.030 79.520 ;
        RECT 109.565 79.460 109.855 79.505 ;
        RECT 107.710 79.320 109.855 79.460 ;
        RECT 107.710 79.260 108.030 79.320 ;
        RECT 109.565 79.275 109.855 79.320 ;
        RECT 5.520 78.640 113.620 79.120 ;
        RECT 22.610 78.240 22.930 78.500 ;
        RECT 23.530 78.440 23.850 78.500 ;
        RECT 24.465 78.440 24.755 78.485 ;
        RECT 23.530 78.300 24.755 78.440 ;
        RECT 23.530 78.240 23.850 78.300 ;
        RECT 24.465 78.255 24.755 78.300 ;
        RECT 26.305 78.440 26.595 78.485 ;
        RECT 26.750 78.440 27.070 78.500 ;
        RECT 26.305 78.300 27.070 78.440 ;
        RECT 26.305 78.255 26.595 78.300 ;
        RECT 26.750 78.240 27.070 78.300 ;
        RECT 76.430 78.440 76.750 78.500 ;
        RECT 78.745 78.440 79.035 78.485 ;
        RECT 76.430 78.300 79.035 78.440 ;
        RECT 76.430 78.240 76.750 78.300 ;
        RECT 78.745 78.255 79.035 78.300 ;
        RECT 81.045 78.440 81.335 78.485 ;
        RECT 83.790 78.440 84.110 78.500 ;
        RECT 81.045 78.300 84.110 78.440 ;
        RECT 81.045 78.255 81.335 78.300 ;
        RECT 83.790 78.240 84.110 78.300 ;
        RECT 89.770 78.440 90.090 78.500 ;
        RECT 96.225 78.440 96.515 78.485 ;
        RECT 101.730 78.440 102.050 78.500 ;
        RECT 104.490 78.440 104.810 78.500 ;
        RECT 89.770 78.300 96.515 78.440 ;
        RECT 89.770 78.240 90.090 78.300 ;
        RECT 96.225 78.255 96.515 78.300 ;
        RECT 99.980 78.300 104.810 78.440 ;
        RECT 9.290 78.100 9.580 78.145 ;
        RECT 11.150 78.100 11.440 78.145 ;
        RECT 13.930 78.100 14.220 78.145 ;
        RECT 9.290 77.960 14.220 78.100 ;
        RECT 9.290 77.915 9.580 77.960 ;
        RECT 11.150 77.915 11.440 77.960 ;
        RECT 13.930 77.915 14.220 77.960 ;
        RECT 21.690 78.100 22.010 78.160 ;
        RECT 27.225 78.100 27.515 78.145 ;
        RECT 21.690 77.960 27.515 78.100 ;
        RECT 21.690 77.900 22.010 77.960 ;
        RECT 27.225 77.915 27.515 77.960 ;
        RECT 51.610 78.100 51.900 78.145 ;
        RECT 53.470 78.100 53.760 78.145 ;
        RECT 56.250 78.100 56.540 78.145 ;
        RECT 51.610 77.960 56.540 78.100 ;
        RECT 51.610 77.915 51.900 77.960 ;
        RECT 53.470 77.915 53.760 77.960 ;
        RECT 56.250 77.915 56.540 77.960 ;
        RECT 58.030 78.100 58.350 78.160 ;
        RECT 61.710 78.100 62.030 78.160 ;
        RECT 58.030 77.960 62.030 78.100 ;
        RECT 58.030 77.900 58.350 77.960 ;
        RECT 61.710 77.900 62.030 77.960 ;
        RECT 68.165 78.100 68.455 78.145 ;
        RECT 93.910 78.100 94.230 78.160 ;
        RECT 68.165 77.960 94.230 78.100 ;
        RECT 68.165 77.915 68.455 77.960 ;
        RECT 93.910 77.900 94.230 77.960 ;
        RECT 8.810 77.560 9.130 77.820 ;
        RECT 10.665 77.760 10.955 77.805 ;
        RECT 11.570 77.760 11.890 77.820 ;
        RECT 10.665 77.620 11.890 77.760 ;
        RECT 10.665 77.575 10.955 77.620 ;
        RECT 11.570 77.560 11.890 77.620 ;
        RECT 13.410 77.760 13.730 77.820 ;
        RECT 13.410 77.620 20.080 77.760 ;
        RECT 13.410 77.560 13.730 77.620 ;
        RECT 19.940 77.465 20.080 77.620 ;
        RECT 22.610 77.560 22.930 77.820 ;
        RECT 23.990 77.760 24.310 77.820 ;
        RECT 25.385 77.760 25.675 77.805 ;
        RECT 23.990 77.620 25.675 77.760 ;
        RECT 23.990 77.560 24.310 77.620 ;
        RECT 25.385 77.575 25.675 77.620 ;
        RECT 46.990 77.760 47.310 77.820 ;
        RECT 51.130 77.760 51.450 77.820 ;
        RECT 46.990 77.620 51.450 77.760 ;
        RECT 46.990 77.560 47.310 77.620 ;
        RECT 51.130 77.560 51.450 77.620 ;
        RECT 59.410 77.760 59.730 77.820 ;
        RECT 60.115 77.760 60.405 77.805 ;
        RECT 63.105 77.760 63.395 77.805 ;
        RECT 59.410 77.620 63.395 77.760 ;
        RECT 59.410 77.560 59.730 77.620 ;
        RECT 60.115 77.575 60.405 77.620 ;
        RECT 63.105 77.575 63.395 77.620 ;
        RECT 64.010 77.560 64.330 77.820 ;
        RECT 79.190 77.760 79.510 77.820 ;
        RECT 80.125 77.760 80.415 77.805 ;
        RECT 93.465 77.760 93.755 77.805 ;
        RECT 97.130 77.760 97.450 77.820 ;
        RECT 98.525 77.760 98.815 77.805 ;
        RECT 79.190 77.620 80.415 77.760 ;
        RECT 79.190 77.560 79.510 77.620 ;
        RECT 80.125 77.575 80.415 77.620 ;
        RECT 90.320 77.620 92.760 77.760 ;
        RECT 90.320 77.480 90.460 77.620 ;
        RECT 13.930 77.420 14.220 77.465 ;
        RECT 11.685 77.280 14.220 77.420 ;
        RECT 11.685 77.125 11.900 77.280 ;
        RECT 13.930 77.235 14.220 77.280 ;
        RECT 19.865 77.235 20.155 77.465 ;
        RECT 23.530 77.220 23.850 77.480 ;
        RECT 26.305 77.420 26.595 77.465 ;
        RECT 27.670 77.420 27.990 77.480 ;
        RECT 26.305 77.280 27.990 77.420 ;
        RECT 26.305 77.235 26.595 77.280 ;
        RECT 27.670 77.220 27.990 77.280 ;
        RECT 41.485 77.420 41.775 77.465 ;
        RECT 41.930 77.420 42.250 77.480 ;
        RECT 44.690 77.420 45.010 77.480 ;
        RECT 41.485 77.280 45.010 77.420 ;
        RECT 41.485 77.235 41.775 77.280 ;
        RECT 41.930 77.220 42.250 77.280 ;
        RECT 44.690 77.220 45.010 77.280 ;
        RECT 52.970 77.220 53.290 77.480 ;
        RECT 56.250 77.420 56.540 77.465 ;
        RECT 54.005 77.280 56.540 77.420 ;
        RECT 9.750 77.080 10.040 77.125 ;
        RECT 11.610 77.080 11.900 77.125 ;
        RECT 9.750 76.940 11.900 77.080 ;
        RECT 9.750 76.895 10.040 76.940 ;
        RECT 11.610 76.895 11.900 76.940 ;
        RECT 12.530 77.080 12.820 77.125 ;
        RECT 15.790 77.080 16.080 77.125 ;
        RECT 19.405 77.080 19.695 77.125 ;
        RECT 12.530 76.940 19.695 77.080 ;
        RECT 12.530 76.895 12.820 76.940 ;
        RECT 15.790 76.895 16.080 76.940 ;
        RECT 19.405 76.895 19.695 76.940 ;
        RECT 22.150 76.880 22.470 77.140 ;
        RECT 24.925 77.080 25.215 77.125 ;
        RECT 26.750 77.080 27.070 77.140 ;
        RECT 54.005 77.125 54.220 77.280 ;
        RECT 56.250 77.235 56.540 77.280 ;
        RECT 62.630 77.220 62.950 77.480 ;
        RECT 64.930 77.220 65.250 77.480 ;
        RECT 65.865 77.235 66.155 77.465 ;
        RECT 24.925 76.940 27.070 77.080 ;
        RECT 24.925 76.895 25.215 76.940 ;
        RECT 26.750 76.880 27.070 76.940 ;
        RECT 52.070 77.080 52.360 77.125 ;
        RECT 53.930 77.080 54.220 77.125 ;
        RECT 52.070 76.940 54.220 77.080 ;
        RECT 52.070 76.895 52.360 76.940 ;
        RECT 53.930 76.895 54.220 76.940 ;
        RECT 54.850 77.080 55.140 77.125 ;
        RECT 56.650 77.080 56.970 77.140 ;
        RECT 58.110 77.080 58.400 77.125 ;
        RECT 54.850 76.940 58.400 77.080 ;
        RECT 62.720 77.080 62.860 77.220 ;
        RECT 65.940 77.080 66.080 77.235 ;
        RECT 66.310 77.220 66.630 77.480 ;
        RECT 66.785 77.420 67.075 77.465 ;
        RECT 67.690 77.420 68.010 77.480 ;
        RECT 69.545 77.420 69.835 77.465 ;
        RECT 66.785 77.280 68.010 77.420 ;
        RECT 66.785 77.235 67.075 77.280 ;
        RECT 67.690 77.220 68.010 77.280 ;
        RECT 68.240 77.280 69.835 77.420 ;
        RECT 62.720 76.940 66.080 77.080 ;
        RECT 54.850 76.895 55.140 76.940 ;
        RECT 56.650 76.880 56.970 76.940 ;
        RECT 58.110 76.895 58.400 76.940 ;
        RECT 17.795 76.740 18.085 76.785 ;
        RECT 23.070 76.740 23.390 76.800 ;
        RECT 17.795 76.600 23.390 76.740 ;
        RECT 17.795 76.555 18.085 76.600 ;
        RECT 23.070 76.540 23.390 76.600 ;
        RECT 41.470 76.740 41.790 76.800 ;
        RECT 41.945 76.740 42.235 76.785 ;
        RECT 41.470 76.600 42.235 76.740 ;
        RECT 41.470 76.540 41.790 76.600 ;
        RECT 41.945 76.555 42.235 76.600 ;
        RECT 60.790 76.540 61.110 76.800 ;
        RECT 61.710 76.740 62.030 76.800 ;
        RECT 64.470 76.740 64.790 76.800 ;
        RECT 68.240 76.740 68.380 77.280 ;
        RECT 69.545 77.235 69.835 77.280 ;
        RECT 76.905 77.420 77.195 77.465 ;
        RECT 78.730 77.420 79.050 77.480 ;
        RECT 76.905 77.280 79.050 77.420 ;
        RECT 76.905 77.235 77.195 77.280 ;
        RECT 78.730 77.220 79.050 77.280 ;
        RECT 79.650 77.220 79.970 77.480 ;
        RECT 90.230 77.220 90.550 77.480 ;
        RECT 92.620 77.465 92.760 77.620 ;
        RECT 93.465 77.620 98.815 77.760 ;
        RECT 93.465 77.575 93.755 77.620 ;
        RECT 97.130 77.560 97.450 77.620 ;
        RECT 98.525 77.575 98.815 77.620 ;
        RECT 99.445 77.760 99.735 77.805 ;
        RECT 99.980 77.760 100.120 78.300 ;
        RECT 101.730 78.240 102.050 78.300 ;
        RECT 104.490 78.240 104.810 78.300 ;
        RECT 101.290 78.100 101.580 78.145 ;
        RECT 103.150 78.100 103.440 78.145 ;
        RECT 105.930 78.100 106.220 78.145 ;
        RECT 101.290 77.960 106.220 78.100 ;
        RECT 101.290 77.915 101.580 77.960 ;
        RECT 103.150 77.915 103.440 77.960 ;
        RECT 105.930 77.915 106.220 77.960 ;
        RECT 99.445 77.620 100.120 77.760 ;
        RECT 99.445 77.575 99.735 77.620 ;
        RECT 102.650 77.560 102.970 77.820 ;
        RECT 103.570 77.760 103.890 77.820 ;
        RECT 109.795 77.760 110.085 77.805 ;
        RECT 103.200 77.620 110.085 77.760 ;
        RECT 91.165 77.235 91.455 77.465 ;
        RECT 92.545 77.235 92.835 77.465 ;
        RECT 98.050 77.420 98.370 77.480 ;
        RECT 100.825 77.420 101.115 77.465 ;
        RECT 103.200 77.420 103.340 77.620 ;
        RECT 103.570 77.560 103.890 77.620 ;
        RECT 109.795 77.575 110.085 77.620 ;
        RECT 105.930 77.420 106.220 77.465 ;
        RECT 98.050 77.280 101.115 77.420 ;
        RECT 81.030 76.880 81.350 77.140 ;
        RECT 91.240 77.080 91.380 77.235 ;
        RECT 98.050 77.220 98.370 77.280 ;
        RECT 100.825 77.235 101.115 77.280 ;
        RECT 101.360 77.280 103.340 77.420 ;
        RECT 103.685 77.280 106.220 77.420 ;
        RECT 101.360 77.080 101.500 77.280 ;
        RECT 103.685 77.125 103.900 77.280 ;
        RECT 105.930 77.235 106.220 77.280 ;
        RECT 107.710 77.125 108.030 77.140 ;
        RECT 91.240 76.940 101.500 77.080 ;
        RECT 101.750 77.080 102.040 77.125 ;
        RECT 103.610 77.080 103.900 77.125 ;
        RECT 101.750 76.940 103.900 77.080 ;
        RECT 101.750 76.895 102.040 76.940 ;
        RECT 103.610 76.895 103.900 76.940 ;
        RECT 104.530 77.080 104.820 77.125 ;
        RECT 107.710 77.080 108.080 77.125 ;
        RECT 104.530 76.940 108.080 77.080 ;
        RECT 104.530 76.895 104.820 76.940 ;
        RECT 107.710 76.895 108.080 76.940 ;
        RECT 107.710 76.880 108.030 76.895 ;
        RECT 61.710 76.600 68.380 76.740 ;
        RECT 61.710 76.540 62.030 76.600 ;
        RECT 64.470 76.540 64.790 76.600 ;
        RECT 69.070 76.540 69.390 76.800 ;
        RECT 77.810 76.540 78.130 76.800 ;
        RECT 87.930 76.740 88.250 76.800 ;
        RECT 89.325 76.740 89.615 76.785 ;
        RECT 87.930 76.600 89.615 76.740 ;
        RECT 87.930 76.540 88.250 76.600 ;
        RECT 89.325 76.555 89.615 76.600 ;
        RECT 91.610 76.540 91.930 76.800 ;
        RECT 97.590 76.740 97.910 76.800 ;
        RECT 98.065 76.740 98.355 76.785 ;
        RECT 97.590 76.600 98.355 76.740 ;
        RECT 97.590 76.540 97.910 76.600 ;
        RECT 98.065 76.555 98.355 76.600 ;
        RECT 5.520 75.920 113.620 76.400 ;
        RECT 16.630 75.520 16.950 75.780 ;
        RECT 18.930 75.520 19.250 75.780 ;
        RECT 25.845 75.720 26.135 75.765 ;
        RECT 26.750 75.720 27.070 75.780 ;
        RECT 25.845 75.580 27.070 75.720 ;
        RECT 25.845 75.535 26.135 75.580 ;
        RECT 26.750 75.520 27.070 75.580 ;
        RECT 45.610 75.720 45.930 75.780 ;
        RECT 49.750 75.720 50.070 75.780 ;
        RECT 52.050 75.720 52.370 75.780 ;
        RECT 45.610 75.580 49.520 75.720 ;
        RECT 45.610 75.520 45.930 75.580 ;
        RECT 7.910 75.380 8.200 75.425 ;
        RECT 9.770 75.380 10.060 75.425 ;
        RECT 7.910 75.240 10.060 75.380 ;
        RECT 7.910 75.195 8.200 75.240 ;
        RECT 9.770 75.195 10.060 75.240 ;
        RECT 10.690 75.380 10.980 75.425 ;
        RECT 12.490 75.380 12.810 75.440 ;
        RECT 13.950 75.380 14.240 75.425 ;
        RECT 10.690 75.240 14.240 75.380 ;
        RECT 10.690 75.195 10.980 75.240 ;
        RECT 6.985 75.040 7.275 75.085 ;
        RECT 8.350 75.040 8.670 75.100 ;
        RECT 6.985 74.900 8.670 75.040 ;
        RECT 9.845 75.040 10.060 75.195 ;
        RECT 12.490 75.180 12.810 75.240 ;
        RECT 13.950 75.195 14.240 75.240 ;
        RECT 15.955 75.380 16.245 75.425 ;
        RECT 19.020 75.380 19.160 75.520 ;
        RECT 24.910 75.380 25.230 75.440 ;
        RECT 41.470 75.425 41.790 75.440 ;
        RECT 15.955 75.240 19.160 75.380 ;
        RECT 15.955 75.195 16.245 75.240 ;
        RECT 12.090 75.040 12.380 75.085 ;
        RECT 9.845 74.900 12.380 75.040 ;
        RECT 6.985 74.855 7.275 74.900 ;
        RECT 8.350 74.840 8.670 74.900 ;
        RECT 12.090 74.855 12.380 74.900 ;
        RECT 15.250 75.040 15.570 75.100 ;
        RECT 18.485 75.040 18.775 75.085 ;
        RECT 15.250 74.900 18.775 75.040 ;
        RECT 15.250 74.840 15.570 74.900 ;
        RECT 18.485 74.855 18.775 74.900 ;
        RECT 7.890 74.700 8.210 74.760 ;
        RECT 8.825 74.700 9.115 74.745 ;
        RECT 7.890 74.560 9.115 74.700 ;
        RECT 7.890 74.500 8.210 74.560 ;
        RECT 8.825 74.515 9.115 74.560 ;
        RECT 7.450 74.360 7.740 74.405 ;
        RECT 9.310 74.360 9.600 74.405 ;
        RECT 12.090 74.360 12.380 74.405 ;
        RECT 7.450 74.220 12.380 74.360 ;
        RECT 7.450 74.175 7.740 74.220 ;
        RECT 9.310 74.175 9.600 74.220 ;
        RECT 12.090 74.175 12.380 74.220 ;
        RECT 18.560 74.020 18.700 74.855 ;
        RECT 19.020 74.360 19.160 75.240 ;
        RECT 24.080 75.240 25.230 75.380 ;
        RECT 22.625 74.855 22.915 75.085 ;
        RECT 23.070 75.040 23.390 75.100 ;
        RECT 24.080 75.085 24.220 75.240 ;
        RECT 24.910 75.180 25.230 75.240 ;
        RECT 38.730 75.380 39.020 75.425 ;
        RECT 40.590 75.380 40.880 75.425 ;
        RECT 38.730 75.240 40.880 75.380 ;
        RECT 38.730 75.195 39.020 75.240 ;
        RECT 40.590 75.195 40.880 75.240 ;
        RECT 23.545 75.040 23.835 75.085 ;
        RECT 23.070 74.900 23.835 75.040 ;
        RECT 19.850 74.500 20.170 74.760 ;
        RECT 22.700 74.700 22.840 74.855 ;
        RECT 23.070 74.840 23.390 74.900 ;
        RECT 23.545 74.855 23.835 74.900 ;
        RECT 24.005 74.855 24.295 75.085 ;
        RECT 24.465 75.040 24.755 75.085 ;
        RECT 26.290 75.040 26.610 75.100 ;
        RECT 33.205 75.040 33.495 75.085 ;
        RECT 24.465 74.900 33.495 75.040 ;
        RECT 24.465 74.855 24.755 74.900 ;
        RECT 26.290 74.840 26.610 74.900 ;
        RECT 33.205 74.855 33.495 74.900 ;
        RECT 33.280 74.700 33.420 74.855 ;
        RECT 33.650 74.840 33.970 75.100 ;
        RECT 34.110 74.840 34.430 75.100 ;
        RECT 35.030 74.840 35.350 75.100 ;
        RECT 39.170 75.040 39.490 75.100 ;
        RECT 39.645 75.040 39.935 75.085 ;
        RECT 39.170 74.900 39.935 75.040 ;
        RECT 40.665 75.040 40.880 75.195 ;
        RECT 41.470 75.380 41.800 75.425 ;
        RECT 44.770 75.380 45.060 75.425 ;
        RECT 41.470 75.240 45.060 75.380 ;
        RECT 49.380 75.380 49.520 75.580 ;
        RECT 49.750 75.580 52.370 75.720 ;
        RECT 49.750 75.520 50.070 75.580 ;
        RECT 52.050 75.520 52.370 75.580 ;
        RECT 52.970 75.720 53.290 75.780 ;
        RECT 54.365 75.720 54.655 75.765 ;
        RECT 52.970 75.580 54.655 75.720 ;
        RECT 52.970 75.520 53.290 75.580 ;
        RECT 54.365 75.535 54.655 75.580 ;
        RECT 56.205 75.720 56.495 75.765 ;
        RECT 56.650 75.720 56.970 75.780 ;
        RECT 63.550 75.720 63.870 75.780 ;
        RECT 56.205 75.580 56.970 75.720 ;
        RECT 56.205 75.535 56.495 75.580 ;
        RECT 56.650 75.520 56.970 75.580 ;
        RECT 60.420 75.580 63.870 75.720 ;
        RECT 51.145 75.380 51.435 75.425 ;
        RECT 51.605 75.380 51.895 75.425 ;
        RECT 49.380 75.240 50.900 75.380 ;
        RECT 41.470 75.195 41.800 75.240 ;
        RECT 44.770 75.195 45.060 75.240 ;
        RECT 41.470 75.180 41.790 75.195 ;
        RECT 42.910 75.040 43.200 75.085 ;
        RECT 40.665 74.900 43.200 75.040 ;
        RECT 39.170 74.840 39.490 74.900 ;
        RECT 39.645 74.855 39.935 74.900 ;
        RECT 42.910 74.855 43.200 74.900 ;
        RECT 47.910 74.840 48.230 75.100 ;
        RECT 48.845 74.855 49.135 75.085 ;
        RECT 49.305 74.855 49.595 75.085 ;
        RECT 49.765 74.855 50.055 75.085 ;
        RECT 50.760 75.040 50.900 75.240 ;
        RECT 51.145 75.240 51.895 75.380 ;
        RECT 51.145 75.195 51.435 75.240 ;
        RECT 51.605 75.195 51.895 75.240 ;
        RECT 50.760 74.900 52.740 75.040 ;
        RECT 34.570 74.700 34.890 74.760 ;
        RECT 36.870 74.700 37.190 74.760 ;
        RECT 37.805 74.700 38.095 74.745 ;
        RECT 22.700 74.560 24.680 74.700 ;
        RECT 33.280 74.560 33.880 74.700 ;
        RECT 24.540 74.420 24.680 74.560 ;
        RECT 23.070 74.360 23.390 74.420 ;
        RECT 19.020 74.220 23.390 74.360 ;
        RECT 23.070 74.160 23.390 74.220 ;
        RECT 24.450 74.160 24.770 74.420 ;
        RECT 25.370 74.020 25.690 74.080 ;
        RECT 18.560 73.880 25.690 74.020 ;
        RECT 25.370 73.820 25.690 73.880 ;
        RECT 31.350 74.020 31.670 74.080 ;
        RECT 31.825 74.020 32.115 74.065 ;
        RECT 31.350 73.880 32.115 74.020 ;
        RECT 33.740 74.020 33.880 74.560 ;
        RECT 34.570 74.560 38.095 74.700 ;
        RECT 34.570 74.500 34.890 74.560 ;
        RECT 36.870 74.500 37.190 74.560 ;
        RECT 37.805 74.515 38.095 74.560 ;
        RECT 45.150 74.700 45.470 74.760 ;
        RECT 46.775 74.700 47.065 74.745 ;
        RECT 48.920 74.700 49.060 74.855 ;
        RECT 45.150 74.560 49.060 74.700 ;
        RECT 45.150 74.500 45.470 74.560 ;
        RECT 46.775 74.515 47.065 74.560 ;
        RECT 38.270 74.360 38.560 74.405 ;
        RECT 40.130 74.360 40.420 74.405 ;
        RECT 42.910 74.360 43.200 74.405 ;
        RECT 38.270 74.220 43.200 74.360 ;
        RECT 49.380 74.360 49.520 74.855 ;
        RECT 49.840 74.700 49.980 74.855 ;
        RECT 51.130 74.700 51.450 74.760 ;
        RECT 49.840 74.560 51.450 74.700 ;
        RECT 51.130 74.500 51.450 74.560 ;
        RECT 51.590 74.500 51.910 74.760 ;
        RECT 52.050 74.500 52.370 74.760 ;
        RECT 52.600 74.700 52.740 74.900 ;
        RECT 52.970 74.840 53.290 75.100 ;
        RECT 55.285 74.855 55.575 75.085 ;
        RECT 55.745 75.040 56.035 75.085 ;
        RECT 58.030 75.040 58.350 75.100 ;
        RECT 60.420 75.085 60.560 75.580 ;
        RECT 63.550 75.520 63.870 75.580 ;
        RECT 78.730 75.520 79.050 75.780 ;
        RECT 79.205 75.720 79.495 75.765 ;
        RECT 81.030 75.720 81.350 75.780 ;
        RECT 79.205 75.580 81.350 75.720 ;
        RECT 79.205 75.535 79.495 75.580 ;
        RECT 81.030 75.520 81.350 75.580 ;
        RECT 88.865 75.720 89.155 75.765 ;
        RECT 92.990 75.720 93.310 75.780 ;
        RECT 88.865 75.580 93.310 75.720 ;
        RECT 88.865 75.535 89.155 75.580 ;
        RECT 92.990 75.520 93.310 75.580 ;
        RECT 93.465 75.720 93.755 75.765 ;
        RECT 95.750 75.720 96.070 75.780 ;
        RECT 96.225 75.720 96.515 75.765 ;
        RECT 93.465 75.580 95.520 75.720 ;
        RECT 93.465 75.535 93.755 75.580 ;
        RECT 61.270 75.380 61.560 75.425 ;
        RECT 63.130 75.380 63.420 75.425 ;
        RECT 61.270 75.240 63.420 75.380 ;
        RECT 61.270 75.195 61.560 75.240 ;
        RECT 63.130 75.195 63.420 75.240 ;
        RECT 64.050 75.380 64.340 75.425 ;
        RECT 67.310 75.380 67.600 75.425 ;
        RECT 69.070 75.380 69.390 75.440 ;
        RECT 64.050 75.240 69.390 75.380 ;
        RECT 64.050 75.195 64.340 75.240 ;
        RECT 67.310 75.195 67.600 75.240 ;
        RECT 55.745 74.900 58.350 75.040 ;
        RECT 55.745 74.855 56.035 74.900 ;
        RECT 55.360 74.700 55.500 74.855 ;
        RECT 58.030 74.840 58.350 74.900 ;
        RECT 60.345 74.855 60.635 75.085 ;
        RECT 60.790 74.840 61.110 75.100 ;
        RECT 63.205 75.040 63.420 75.195 ;
        RECT 69.070 75.180 69.390 75.240 ;
        RECT 76.445 75.380 76.735 75.425 ;
        RECT 77.350 75.380 77.670 75.440 ;
        RECT 76.445 75.240 81.720 75.380 ;
        RECT 76.445 75.195 76.735 75.240 ;
        RECT 77.350 75.180 77.670 75.240 ;
        RECT 81.580 75.100 81.720 75.240 ;
        RECT 82.040 75.240 88.160 75.380 ;
        RECT 65.450 75.040 65.740 75.085 ;
        RECT 63.205 74.900 65.740 75.040 ;
        RECT 65.450 74.855 65.740 74.900 ;
        RECT 71.370 75.040 71.690 75.100 ;
        RECT 71.845 75.040 72.135 75.085 ;
        RECT 71.370 74.900 72.135 75.040 ;
        RECT 71.370 74.840 71.690 74.900 ;
        RECT 71.845 74.855 72.135 74.900 ;
        RECT 72.305 75.040 72.595 75.085 ;
        RECT 73.670 75.040 73.990 75.100 ;
        RECT 76.905 75.040 77.195 75.085 ;
        RECT 72.305 74.900 77.195 75.040 ;
        RECT 72.305 74.855 72.595 74.900 ;
        RECT 73.670 74.840 73.990 74.900 ;
        RECT 76.905 74.855 77.195 74.900 ;
        RECT 78.270 75.040 78.590 75.100 ;
        RECT 80.585 75.040 80.875 75.085 ;
        RECT 78.270 74.900 80.875 75.040 ;
        RECT 78.270 74.840 78.590 74.900 ;
        RECT 80.585 74.855 80.875 74.900 ;
        RECT 81.030 74.840 81.350 75.100 ;
        RECT 81.490 74.840 81.810 75.100 ;
        RECT 60.880 74.700 61.020 74.840 ;
        RECT 52.600 74.560 54.120 74.700 ;
        RECT 55.360 74.560 61.020 74.700 ;
        RECT 61.250 74.700 61.570 74.760 ;
        RECT 62.185 74.700 62.475 74.745 ;
        RECT 61.250 74.560 62.475 74.700 ;
        RECT 49.750 74.360 50.070 74.420 ;
        RECT 49.380 74.220 50.070 74.360 ;
        RECT 51.680 74.360 51.820 74.500 ;
        RECT 53.980 74.405 54.120 74.560 ;
        RECT 61.250 74.500 61.570 74.560 ;
        RECT 62.185 74.515 62.475 74.560 ;
        RECT 64.010 74.700 64.330 74.760 ;
        RECT 72.765 74.700 73.055 74.745 ;
        RECT 75.525 74.700 75.815 74.745 ;
        RECT 64.010 74.560 75.815 74.700 ;
        RECT 64.010 74.500 64.330 74.560 ;
        RECT 72.765 74.515 73.055 74.560 ;
        RECT 75.525 74.515 75.815 74.560 ;
        RECT 75.970 74.700 76.290 74.760 ;
        RECT 82.040 74.700 82.180 75.240 ;
        RECT 82.410 74.840 82.730 75.100 ;
        RECT 83.790 75.040 84.110 75.100 ;
        RECT 84.265 75.040 84.555 75.085 ;
        RECT 86.090 75.040 86.410 75.100 ;
        RECT 83.790 74.900 86.410 75.040 ;
        RECT 83.790 74.840 84.110 74.900 ;
        RECT 84.265 74.855 84.555 74.900 ;
        RECT 86.090 74.840 86.410 74.900 ;
        RECT 86.565 75.040 86.855 75.085 ;
        RECT 87.470 75.040 87.790 75.100 ;
        RECT 88.020 75.085 88.160 75.240 ;
        RECT 93.910 75.180 94.230 75.440 ;
        RECT 95.380 75.380 95.520 75.580 ;
        RECT 95.750 75.580 96.515 75.720 ;
        RECT 95.750 75.520 96.070 75.580 ;
        RECT 96.225 75.535 96.515 75.580 ;
        RECT 98.970 75.520 99.290 75.780 ;
        RECT 103.570 75.720 103.890 75.780 ;
        RECT 105.425 75.720 105.715 75.765 ;
        RECT 103.570 75.580 105.715 75.720 ;
        RECT 103.570 75.520 103.890 75.580 ;
        RECT 105.425 75.535 105.715 75.580 ;
        RECT 105.870 75.520 106.190 75.780 ;
        RECT 107.250 75.720 107.570 75.780 ;
        RECT 107.725 75.720 108.015 75.765 ;
        RECT 107.250 75.580 108.015 75.720 ;
        RECT 107.250 75.520 107.570 75.580 ;
        RECT 107.725 75.535 108.015 75.580 ;
        RECT 98.510 75.380 98.830 75.440 ;
        RECT 95.380 75.240 98.830 75.380 ;
        RECT 98.510 75.180 98.830 75.240 ;
        RECT 86.565 74.900 87.790 75.040 ;
        RECT 86.565 74.855 86.855 74.900 ;
        RECT 87.470 74.840 87.790 74.900 ;
        RECT 87.945 74.855 88.235 75.085 ;
        RECT 91.165 74.855 91.455 75.085 ;
        RECT 92.545 75.040 92.835 75.085 ;
        RECT 93.450 75.040 93.770 75.100 ;
        RECT 92.545 74.900 93.770 75.040 ;
        RECT 92.545 74.855 92.835 74.900 ;
        RECT 75.970 74.560 82.180 74.700 ;
        RECT 75.970 74.500 76.290 74.560 ;
        RECT 87.010 74.500 87.330 74.760 ;
        RECT 51.680 74.220 52.280 74.360 ;
        RECT 38.270 74.175 38.560 74.220 ;
        RECT 40.130 74.175 40.420 74.220 ;
        RECT 42.910 74.175 43.200 74.220 ;
        RECT 49.750 74.160 50.070 74.220 ;
        RECT 51.590 74.020 51.910 74.080 ;
        RECT 52.140 74.065 52.280 74.220 ;
        RECT 53.905 74.175 54.195 74.405 ;
        RECT 60.810 74.360 61.100 74.405 ;
        RECT 62.670 74.360 62.960 74.405 ;
        RECT 65.450 74.360 65.740 74.405 ;
        RECT 60.810 74.220 65.740 74.360 ;
        RECT 60.810 74.175 61.100 74.220 ;
        RECT 62.670 74.175 62.960 74.220 ;
        RECT 65.450 74.175 65.740 74.220 ;
        RECT 66.770 74.360 67.090 74.420 ;
        RECT 69.315 74.360 69.605 74.405 ;
        RECT 71.370 74.360 71.690 74.420 ;
        RECT 66.770 74.220 71.690 74.360 ;
        RECT 66.770 74.160 67.090 74.220 ;
        RECT 69.315 74.175 69.605 74.220 ;
        RECT 71.370 74.160 71.690 74.220 ;
        RECT 72.290 74.360 72.610 74.420 ;
        RECT 91.240 74.360 91.380 74.855 ;
        RECT 93.450 74.840 93.770 74.900 ;
        RECT 95.290 74.840 95.610 75.100 ;
        RECT 96.670 74.840 96.990 75.100 ;
        RECT 98.050 74.840 98.370 75.100 ;
        RECT 92.070 74.500 92.390 74.760 ;
        RECT 94.385 74.700 94.675 74.745 ;
        RECT 94.000 74.560 94.675 74.700 ;
        RECT 94.000 74.420 94.140 74.560 ;
        RECT 94.385 74.515 94.675 74.560 ;
        RECT 97.130 74.500 97.450 74.760 ;
        RECT 104.490 74.500 104.810 74.760 ;
        RECT 72.290 74.220 91.380 74.360 ;
        RECT 72.290 74.160 72.610 74.220 ;
        RECT 93.910 74.160 94.230 74.420 ;
        RECT 33.740 73.880 51.910 74.020 ;
        RECT 31.350 73.820 31.670 73.880 ;
        RECT 31.825 73.835 32.115 73.880 ;
        RECT 51.590 73.820 51.910 73.880 ;
        RECT 52.065 73.835 52.355 74.065 ;
        RECT 70.005 74.020 70.295 74.065 ;
        RECT 71.830 74.020 72.150 74.080 ;
        RECT 70.005 73.880 72.150 74.020 ;
        RECT 70.005 73.835 70.295 73.880 ;
        RECT 71.830 73.820 72.150 73.880 ;
        RECT 74.130 74.020 74.450 74.080 ;
        RECT 80.570 74.020 80.890 74.080 ;
        RECT 74.130 73.880 80.890 74.020 ;
        RECT 74.130 73.820 74.450 73.880 ;
        RECT 80.570 73.820 80.890 73.880 ;
        RECT 83.790 73.820 84.110 74.080 ;
        RECT 87.930 73.820 88.250 74.080 ;
        RECT 91.610 73.820 91.930 74.080 ;
        RECT 94.370 73.820 94.690 74.080 ;
        RECT 94.830 74.020 95.150 74.080 ;
        RECT 96.685 74.020 96.975 74.065 ;
        RECT 94.830 73.880 96.975 74.020 ;
        RECT 94.830 73.820 95.150 73.880 ;
        RECT 96.685 73.835 96.975 73.880 ;
        RECT 5.520 73.200 113.620 73.680 ;
        RECT 12.490 72.800 12.810 73.060 ;
        RECT 20.785 73.000 21.075 73.045 ;
        RECT 22.150 73.000 22.470 73.060 ;
        RECT 20.785 72.860 22.470 73.000 ;
        RECT 20.785 72.815 21.075 72.860 ;
        RECT 22.150 72.800 22.470 72.860 ;
        RECT 28.130 72.800 28.450 73.060 ;
        RECT 29.510 73.000 29.830 73.060 ;
        RECT 30.445 73.000 30.735 73.045 ;
        RECT 29.510 72.860 30.735 73.000 ;
        RECT 29.510 72.800 29.830 72.860 ;
        RECT 30.445 72.815 30.735 72.860 ;
        RECT 31.810 72.800 32.130 73.060 ;
        RECT 33.190 73.000 33.510 73.060 ;
        RECT 34.125 73.000 34.415 73.045 ;
        RECT 64.010 73.000 64.330 73.060 ;
        RECT 33.190 72.860 34.415 73.000 ;
        RECT 33.190 72.800 33.510 72.860 ;
        RECT 34.125 72.815 34.415 72.860 ;
        RECT 34.660 72.860 57.340 73.000 ;
        RECT 21.690 72.660 22.010 72.720 ;
        RECT 24.910 72.660 25.230 72.720 ;
        RECT 33.650 72.660 33.970 72.720 ;
        RECT 34.660 72.660 34.800 72.860 ;
        RECT 21.690 72.520 34.800 72.660 ;
        RECT 35.050 72.660 35.340 72.705 ;
        RECT 36.910 72.660 37.200 72.705 ;
        RECT 39.690 72.660 39.980 72.705 ;
        RECT 35.050 72.520 39.980 72.660 ;
        RECT 21.690 72.460 22.010 72.520 ;
        RECT 24.910 72.460 25.230 72.520 ;
        RECT 12.965 71.980 13.255 72.025 ;
        RECT 13.410 71.980 13.730 72.040 ;
        RECT 21.935 71.980 22.225 72.025 ;
        RECT 12.965 71.840 13.730 71.980 ;
        RECT 12.965 71.795 13.255 71.840 ;
        RECT 13.410 71.780 13.730 71.840 ;
        RECT 21.320 71.840 22.225 71.980 ;
        RECT 21.320 71.300 21.460 71.840 ;
        RECT 21.935 71.795 22.225 71.840 ;
        RECT 22.625 71.795 22.915 72.025 ;
        RECT 23.070 72.010 23.390 72.040 ;
        RECT 23.070 71.965 23.400 72.010 ;
        RECT 24.005 71.980 24.295 72.025 ;
        RECT 24.450 71.980 24.770 72.040 ;
        RECT 23.070 71.825 23.570 71.965 ;
        RECT 24.005 71.840 24.770 71.980 ;
        RECT 22.700 71.640 22.840 71.795 ;
        RECT 23.070 71.780 23.400 71.825 ;
        RECT 24.005 71.795 24.295 71.840 ;
        RECT 24.450 71.780 24.770 71.840 ;
        RECT 25.370 71.780 25.690 72.040 ;
        RECT 25.920 72.025 26.060 72.520 ;
        RECT 33.650 72.460 33.970 72.520 ;
        RECT 35.050 72.475 35.340 72.520 ;
        RECT 36.910 72.475 37.200 72.520 ;
        RECT 39.690 72.475 39.980 72.520 ;
        RECT 50.210 72.460 50.530 72.720 ;
        RECT 28.130 72.320 28.450 72.380 ;
        RECT 26.380 72.180 28.450 72.320 ;
        RECT 26.380 72.040 26.520 72.180 ;
        RECT 28.130 72.120 28.450 72.180 ;
        RECT 32.270 72.120 32.590 72.380 ;
        RECT 34.570 72.120 34.890 72.380 ;
        RECT 36.425 72.320 36.715 72.365 ;
        RECT 43.310 72.320 43.630 72.380 ;
        RECT 36.425 72.180 43.630 72.320 ;
        RECT 36.425 72.135 36.715 72.180 ;
        RECT 43.310 72.120 43.630 72.180 ;
        RECT 47.910 72.120 48.230 72.380 ;
        RECT 48.370 72.320 48.690 72.380 ;
        RECT 50.300 72.320 50.440 72.460 ;
        RECT 53.890 72.320 54.210 72.380 ;
        RECT 48.370 72.180 54.210 72.320 ;
        RECT 57.200 72.320 57.340 72.860 ;
        RECT 59.960 72.860 64.330 73.000 ;
        RECT 59.960 72.720 60.100 72.860 ;
        RECT 64.010 72.800 64.330 72.860 ;
        RECT 65.405 73.000 65.695 73.045 ;
        RECT 72.290 73.000 72.610 73.060 ;
        RECT 65.405 72.860 72.610 73.000 ;
        RECT 65.405 72.815 65.695 72.860 ;
        RECT 72.290 72.800 72.610 72.860 ;
        RECT 72.750 73.000 73.070 73.060 ;
        RECT 74.590 73.000 74.910 73.060 ;
        RECT 81.030 73.000 81.350 73.060 ;
        RECT 72.750 72.860 81.350 73.000 ;
        RECT 72.750 72.800 73.070 72.860 ;
        RECT 74.590 72.800 74.910 72.860 ;
        RECT 81.030 72.800 81.350 72.860 ;
        RECT 81.490 73.000 81.810 73.060 ;
        RECT 85.875 73.000 86.165 73.045 ;
        RECT 81.490 72.860 86.165 73.000 ;
        RECT 81.490 72.800 81.810 72.860 ;
        RECT 85.875 72.815 86.165 72.860 ;
        RECT 94.370 72.800 94.690 73.060 ;
        RECT 57.585 72.660 57.875 72.705 ;
        RECT 59.870 72.660 60.190 72.720 ;
        RECT 57.585 72.520 60.190 72.660 ;
        RECT 57.585 72.475 57.875 72.520 ;
        RECT 59.870 72.460 60.190 72.520 ;
        RECT 61.725 72.660 62.015 72.705 ;
        RECT 63.550 72.660 63.870 72.720 ;
        RECT 75.970 72.660 76.290 72.720 ;
        RECT 61.725 72.520 76.290 72.660 ;
        RECT 61.725 72.475 62.015 72.520 ;
        RECT 63.550 72.460 63.870 72.520 ;
        RECT 75.970 72.460 76.290 72.520 ;
        RECT 77.370 72.660 77.660 72.705 ;
        RECT 79.230 72.660 79.520 72.705 ;
        RECT 82.010 72.660 82.300 72.705 ;
        RECT 96.670 72.660 96.990 72.720 ;
        RECT 77.370 72.520 82.300 72.660 ;
        RECT 77.370 72.475 77.660 72.520 ;
        RECT 79.230 72.475 79.520 72.520 ;
        RECT 82.010 72.475 82.300 72.520 ;
        RECT 82.960 72.520 96.990 72.660 ;
        RECT 58.030 72.320 58.350 72.380 ;
        RECT 66.310 72.320 66.630 72.380 ;
        RECT 69.085 72.320 69.375 72.365 ;
        RECT 57.200 72.180 67.460 72.320 ;
        RECT 48.370 72.120 48.690 72.180 ;
        RECT 25.845 71.795 26.135 72.025 ;
        RECT 25.920 71.640 26.060 71.795 ;
        RECT 26.290 71.780 26.610 72.040 ;
        RECT 29.050 71.780 29.370 72.040 ;
        RECT 29.525 71.795 29.815 72.025 ;
        RECT 31.350 71.980 31.670 72.040 ;
        RECT 31.825 71.980 32.115 72.025 ;
        RECT 31.350 71.840 32.115 71.980 ;
        RECT 22.700 71.500 26.060 71.640 ;
        RECT 22.150 71.300 22.470 71.360 ;
        RECT 26.380 71.300 26.520 71.780 ;
        RECT 27.685 71.640 27.975 71.685 ;
        RECT 28.145 71.640 28.435 71.685 ;
        RECT 27.685 71.500 28.435 71.640 ;
        RECT 27.685 71.455 27.975 71.500 ;
        RECT 28.145 71.455 28.435 71.500 ;
        RECT 21.320 71.160 26.520 71.300 ;
        RECT 27.210 71.300 27.530 71.360 ;
        RECT 29.600 71.300 29.740 71.795 ;
        RECT 31.350 71.780 31.670 71.840 ;
        RECT 31.825 71.795 32.115 71.840 ;
        RECT 33.205 71.980 33.495 72.025 ;
        RECT 33.650 71.980 33.970 72.040 ;
        RECT 39.690 71.980 39.980 72.025 ;
        RECT 33.205 71.840 33.970 71.980 ;
        RECT 33.205 71.795 33.495 71.840 ;
        RECT 33.650 71.780 33.970 71.840 ;
        RECT 37.445 71.840 39.980 71.980 ;
        RECT 37.445 71.685 37.660 71.840 ;
        RECT 39.690 71.795 39.980 71.840 ;
        RECT 45.150 71.980 45.470 72.040 ;
        RECT 48.920 72.025 49.060 72.180 ;
        RECT 53.890 72.120 54.210 72.180 ;
        RECT 58.030 72.120 58.350 72.180 ;
        RECT 46.545 71.980 46.835 72.025 ;
        RECT 45.150 71.840 46.835 71.980 ;
        RECT 45.150 71.780 45.470 71.840 ;
        RECT 46.545 71.795 46.835 71.840 ;
        RECT 48.845 71.795 49.135 72.025 ;
        RECT 49.765 71.795 50.055 72.025 ;
        RECT 41.470 71.685 41.790 71.700 ;
        RECT 35.510 71.640 35.800 71.685 ;
        RECT 37.370 71.640 37.660 71.685 ;
        RECT 35.510 71.500 37.660 71.640 ;
        RECT 35.510 71.455 35.800 71.500 ;
        RECT 37.370 71.455 37.660 71.500 ;
        RECT 38.290 71.640 38.580 71.685 ;
        RECT 41.470 71.640 41.840 71.685 ;
        RECT 38.290 71.500 41.840 71.640 ;
        RECT 38.290 71.455 38.580 71.500 ;
        RECT 41.470 71.455 41.840 71.500 ;
        RECT 42.850 71.640 43.170 71.700 ;
        RECT 43.555 71.640 43.845 71.685 ;
        RECT 47.005 71.640 47.295 71.685 ;
        RECT 49.840 71.640 49.980 71.795 ;
        RECT 50.210 71.780 50.530 72.040 ;
        RECT 50.685 71.980 50.975 72.025 ;
        RECT 51.130 71.980 51.450 72.040 ;
        RECT 50.685 71.840 56.880 71.980 ;
        RECT 50.685 71.795 50.975 71.840 ;
        RECT 51.130 71.780 51.450 71.840 ;
        RECT 42.850 71.500 49.980 71.640 ;
        RECT 51.590 71.640 51.910 71.700 ;
        RECT 56.205 71.640 56.495 71.685 ;
        RECT 51.590 71.500 56.495 71.640 ;
        RECT 41.470 71.440 41.790 71.455 ;
        RECT 42.850 71.440 43.170 71.500 ;
        RECT 43.555 71.455 43.845 71.500 ;
        RECT 47.005 71.455 47.295 71.500 ;
        RECT 51.590 71.440 51.910 71.500 ;
        RECT 56.205 71.455 56.495 71.500 ;
        RECT 27.210 71.160 29.740 71.300 ;
        RECT 44.230 71.300 44.550 71.360 ;
        RECT 44.705 71.300 44.995 71.345 ;
        RECT 44.230 71.160 44.995 71.300 ;
        RECT 22.150 71.100 22.470 71.160 ;
        RECT 27.210 71.100 27.530 71.160 ;
        RECT 44.230 71.100 44.550 71.160 ;
        RECT 44.705 71.115 44.995 71.160 ;
        RECT 50.210 71.300 50.530 71.360 ;
        RECT 52.065 71.300 52.355 71.345 ;
        RECT 50.210 71.160 52.355 71.300 ;
        RECT 56.740 71.300 56.880 71.840 ;
        RECT 58.490 71.780 58.810 72.040 ;
        RECT 59.410 71.780 59.730 72.040 ;
        RECT 59.960 72.025 60.100 72.180 ;
        RECT 59.885 71.795 60.175 72.025 ;
        RECT 60.330 71.780 60.650 72.040 ;
        RECT 62.185 71.990 62.475 72.025 ;
        RECT 62.630 71.990 62.950 72.040 ;
        RECT 62.185 71.850 62.950 71.990 ;
        RECT 62.185 71.795 62.475 71.850 ;
        RECT 62.630 71.780 62.950 71.850 ;
        RECT 63.090 71.780 63.410 72.040 ;
        RECT 63.640 72.025 63.780 72.180 ;
        RECT 66.310 72.120 66.630 72.180 ;
        RECT 63.565 71.795 63.855 72.025 ;
        RECT 64.010 71.780 64.330 72.040 ;
        RECT 64.930 71.980 65.250 72.040 ;
        RECT 65.865 71.980 66.155 72.025 ;
        RECT 64.930 71.840 66.155 71.980 ;
        RECT 64.930 71.780 65.250 71.840 ;
        RECT 65.865 71.795 66.155 71.840 ;
        RECT 66.770 71.780 67.090 72.040 ;
        RECT 67.320 72.025 67.460 72.180 ;
        RECT 69.085 72.180 76.660 72.320 ;
        RECT 69.085 72.135 69.375 72.180 ;
        RECT 67.245 71.795 67.535 72.025 ;
        RECT 67.690 71.780 68.010 72.040 ;
        RECT 71.385 71.980 71.675 72.025 ;
        RECT 71.830 71.980 72.150 72.040 ;
        RECT 71.385 71.840 72.150 71.980 ;
        RECT 71.385 71.795 71.675 71.840 ;
        RECT 71.830 71.780 72.150 71.840 ;
        RECT 72.290 71.980 72.610 72.040 ;
        RECT 72.765 71.980 73.055 72.025 ;
        RECT 72.290 71.840 73.055 71.980 ;
        RECT 72.290 71.780 72.610 71.840 ;
        RECT 72.765 71.795 73.055 71.840 ;
        RECT 73.670 71.780 73.990 72.040 ;
        RECT 74.130 71.780 74.450 72.040 ;
        RECT 74.605 71.990 74.895 72.025 ;
        RECT 74.605 71.850 75.740 71.990 ;
        RECT 74.605 71.795 74.895 71.850 ;
        RECT 64.100 71.640 64.240 71.780 ;
        RECT 67.780 71.640 67.920 71.780 ;
        RECT 64.100 71.500 67.920 71.640 ;
        RECT 75.600 71.640 75.740 71.850 ;
        RECT 76.520 71.980 76.660 72.180 ;
        RECT 76.890 72.120 77.210 72.380 ;
        RECT 77.810 72.320 78.130 72.380 ;
        RECT 78.745 72.320 79.035 72.365 ;
        RECT 82.960 72.320 83.100 72.520 ;
        RECT 96.670 72.460 96.990 72.520 ;
        RECT 77.810 72.180 79.035 72.320 ;
        RECT 77.810 72.120 78.130 72.180 ;
        RECT 78.745 72.135 79.035 72.180 ;
        RECT 79.280 72.180 83.100 72.320 ;
        RECT 92.545 72.320 92.835 72.365 ;
        RECT 97.590 72.320 97.910 72.380 ;
        RECT 92.545 72.180 97.910 72.320 ;
        RECT 79.280 71.980 79.420 72.180 ;
        RECT 92.545 72.135 92.835 72.180 ;
        RECT 97.590 72.120 97.910 72.180 ;
        RECT 82.010 71.980 82.300 72.025 ;
        RECT 76.520 71.840 79.420 71.980 ;
        RECT 79.765 71.840 82.300 71.980 ;
        RECT 77.350 71.640 77.670 71.700 ;
        RECT 79.765 71.685 79.980 71.840 ;
        RECT 82.010 71.795 82.300 71.840 ;
        RECT 90.230 71.980 90.550 72.040 ;
        RECT 93.465 71.980 93.755 72.025 ;
        RECT 90.230 71.840 93.755 71.980 ;
        RECT 90.230 71.780 90.550 71.840 ;
        RECT 93.465 71.795 93.755 71.840 ;
        RECT 83.790 71.685 84.110 71.700 ;
        RECT 75.600 71.500 77.670 71.640 ;
        RECT 77.350 71.440 77.670 71.500 ;
        RECT 77.830 71.640 78.120 71.685 ;
        RECT 79.690 71.640 79.980 71.685 ;
        RECT 77.830 71.500 79.980 71.640 ;
        RECT 77.830 71.455 78.120 71.500 ;
        RECT 79.690 71.455 79.980 71.500 ;
        RECT 80.610 71.640 80.900 71.685 ;
        RECT 83.790 71.640 84.160 71.685 ;
        RECT 80.610 71.500 84.160 71.640 ;
        RECT 80.610 71.455 80.900 71.500 ;
        RECT 83.790 71.455 84.160 71.500 ;
        RECT 83.790 71.440 84.110 71.455 ;
        RECT 64.470 71.300 64.790 71.360 ;
        RECT 56.740 71.160 64.790 71.300 ;
        RECT 50.210 71.100 50.530 71.160 ;
        RECT 52.065 71.115 52.355 71.160 ;
        RECT 64.470 71.100 64.790 71.160 ;
        RECT 70.450 71.100 70.770 71.360 ;
        RECT 75.985 71.300 76.275 71.345 ;
        RECT 79.190 71.300 79.510 71.360 ;
        RECT 75.985 71.160 79.510 71.300 ;
        RECT 75.985 71.115 76.275 71.160 ;
        RECT 79.190 71.100 79.510 71.160 ;
        RECT 86.090 71.300 86.410 71.360 ;
        RECT 94.370 71.300 94.690 71.360 ;
        RECT 86.090 71.160 94.690 71.300 ;
        RECT 86.090 71.100 86.410 71.160 ;
        RECT 94.370 71.100 94.690 71.160 ;
        RECT 5.520 70.480 113.620 70.960 ;
        RECT 14.805 70.280 15.095 70.325 ;
        RECT 16.630 70.280 16.950 70.340 ;
        RECT 14.805 70.140 23.300 70.280 ;
        RECT 14.805 70.095 15.095 70.140 ;
        RECT 16.630 70.080 16.950 70.140 ;
        RECT 17.550 69.940 17.870 70.000 ;
        RECT 19.850 69.940 20.170 70.000 ;
        RECT 16.260 69.800 20.170 69.940 ;
        RECT 15.250 69.060 15.570 69.320 ;
        RECT 16.260 69.305 16.400 69.800 ;
        RECT 17.550 69.740 17.870 69.800 ;
        RECT 19.850 69.740 20.170 69.800 ;
        RECT 20.325 69.940 20.615 69.985 ;
        RECT 20.785 69.940 21.075 69.985 ;
        RECT 20.325 69.800 21.075 69.940 ;
        RECT 20.325 69.755 20.615 69.800 ;
        RECT 20.785 69.755 21.075 69.800 ;
        RECT 21.690 69.940 22.010 70.000 ;
        RECT 21.690 69.800 22.840 69.940 ;
        RECT 21.690 69.740 22.010 69.800 ;
        RECT 18.945 69.600 19.235 69.645 ;
        RECT 18.945 69.460 21.000 69.600 ;
        RECT 18.945 69.415 19.235 69.460 ;
        RECT 20.860 69.320 21.000 69.460 ;
        RECT 22.150 69.400 22.470 69.660 ;
        RECT 22.700 69.645 22.840 69.800 ;
        RECT 23.160 69.645 23.300 70.140 ;
        RECT 26.750 70.080 27.070 70.340 ;
        RECT 30.890 70.280 31.210 70.340 ;
        RECT 34.125 70.280 34.415 70.325 ;
        RECT 30.890 70.140 34.415 70.280 ;
        RECT 30.890 70.080 31.210 70.140 ;
        RECT 34.125 70.095 34.415 70.140 ;
        RECT 39.185 70.095 39.475 70.325 ;
        RECT 41.025 70.280 41.315 70.325 ;
        RECT 42.850 70.280 43.170 70.340 ;
        RECT 41.025 70.140 43.170 70.280 ;
        RECT 41.025 70.095 41.315 70.140 ;
        RECT 26.840 69.940 26.980 70.080 ;
        RECT 25.460 69.800 26.980 69.940 ;
        RECT 28.605 69.940 28.895 69.985 ;
        RECT 31.825 69.940 32.115 69.985 ;
        RECT 28.605 69.800 32.115 69.940 ;
        RECT 25.460 69.645 25.600 69.800 ;
        RECT 28.605 69.755 28.895 69.800 ;
        RECT 31.825 69.755 32.115 69.800 ;
        RECT 22.625 69.415 22.915 69.645 ;
        RECT 23.085 69.415 23.375 69.645 ;
        RECT 24.005 69.600 24.295 69.645 ;
        RECT 25.385 69.600 25.675 69.645 ;
        RECT 24.005 69.460 25.675 69.600 ;
        RECT 24.005 69.415 24.295 69.460 ;
        RECT 25.385 69.415 25.675 69.460 ;
        RECT 16.185 69.075 16.475 69.305 ;
        RECT 18.010 69.060 18.330 69.320 ;
        RECT 19.850 69.060 20.170 69.320 ;
        RECT 20.770 69.060 21.090 69.320 ;
        RECT 22.700 69.260 22.840 69.415 ;
        RECT 26.290 69.400 26.610 69.660 ;
        RECT 26.765 69.415 27.055 69.645 ;
        RECT 27.225 69.600 27.515 69.645 ;
        RECT 28.130 69.600 28.450 69.660 ;
        RECT 27.225 69.460 28.450 69.600 ;
        RECT 27.225 69.415 27.515 69.460 ;
        RECT 26.840 69.260 26.980 69.415 ;
        RECT 28.130 69.400 28.450 69.460 ;
        RECT 33.190 69.400 33.510 69.660 ;
        RECT 37.805 69.600 38.095 69.645 ;
        RECT 39.260 69.600 39.400 70.095 ;
        RECT 42.850 70.080 43.170 70.140 ;
        RECT 43.310 70.080 43.630 70.340 ;
        RECT 51.590 70.080 51.910 70.340 ;
        RECT 52.510 70.080 52.830 70.340 ;
        RECT 53.890 70.280 54.210 70.340 ;
        RECT 59.425 70.280 59.715 70.325 ;
        RECT 53.890 70.140 59.715 70.280 ;
        RECT 53.890 70.080 54.210 70.140 ;
        RECT 59.425 70.095 59.715 70.140 ;
        RECT 41.470 69.940 41.790 70.000 ;
        RECT 45.165 69.940 45.455 69.985 ;
        RECT 41.470 69.800 45.455 69.940 ;
        RECT 41.470 69.740 41.790 69.800 ;
        RECT 45.165 69.755 45.455 69.800 ;
        RECT 50.210 69.740 50.530 70.000 ;
        RECT 51.680 69.940 51.820 70.080 ;
        RECT 54.810 69.940 55.130 70.000 ;
        RECT 51.680 69.800 55.130 69.940 ;
        RECT 59.500 69.940 59.640 70.095 ;
        RECT 61.250 70.080 61.570 70.340 ;
        RECT 62.170 70.280 62.490 70.340 ;
        RECT 63.550 70.280 63.870 70.340 ;
        RECT 72.290 70.280 72.610 70.340 ;
        RECT 62.170 70.140 63.870 70.280 ;
        RECT 62.170 70.080 62.490 70.140 ;
        RECT 63.550 70.080 63.870 70.140 ;
        RECT 64.100 70.140 72.610 70.280 ;
        RECT 64.100 69.940 64.240 70.140 ;
        RECT 72.290 70.080 72.610 70.140 ;
        RECT 73.670 70.280 73.990 70.340 ;
        RECT 76.445 70.280 76.735 70.325 ;
        RECT 73.670 70.140 76.735 70.280 ;
        RECT 73.670 70.080 73.990 70.140 ;
        RECT 76.445 70.095 76.735 70.140 ;
        RECT 76.905 70.095 77.195 70.325 ;
        RECT 59.500 69.800 64.240 69.940 ;
        RECT 69.085 69.940 69.375 69.985 ;
        RECT 70.450 69.940 70.770 70.000 ;
        RECT 69.085 69.800 70.770 69.940 ;
        RECT 54.810 69.740 55.130 69.800 ;
        RECT 69.085 69.755 69.375 69.800 ;
        RECT 70.450 69.740 70.770 69.800 ;
        RECT 71.365 69.940 72.015 69.985 ;
        RECT 72.750 69.940 73.070 70.000 ;
        RECT 74.965 69.940 75.255 69.985 ;
        RECT 71.365 69.800 75.255 69.940 ;
        RECT 71.365 69.755 72.015 69.800 ;
        RECT 72.750 69.740 73.070 69.800 ;
        RECT 74.665 69.755 75.255 69.800 ;
        RECT 37.805 69.460 39.400 69.600 ;
        RECT 37.805 69.415 38.095 69.460 ;
        RECT 44.230 69.400 44.550 69.660 ;
        RECT 44.690 69.400 45.010 69.660 ;
        RECT 51.590 69.400 51.910 69.660 ;
        RECT 59.870 69.600 60.190 69.660 ;
        RECT 60.345 69.600 60.635 69.645 ;
        RECT 59.870 69.460 60.635 69.600 ;
        RECT 59.870 69.400 60.190 69.460 ;
        RECT 60.345 69.415 60.635 69.460 ;
        RECT 62.170 69.400 62.490 69.660 ;
        RECT 62.630 69.400 62.950 69.660 ;
        RECT 63.105 69.415 63.395 69.645 ;
        RECT 64.025 69.600 64.315 69.645 ;
        RECT 66.770 69.600 67.090 69.660 ;
        RECT 64.025 69.460 67.090 69.600 ;
        RECT 64.025 69.415 64.315 69.460 ;
        RECT 22.700 69.120 26.980 69.260 ;
        RECT 29.510 69.260 29.830 69.320 ;
        RECT 32.285 69.260 32.575 69.305 ;
        RECT 29.510 69.120 32.575 69.260 ;
        RECT 29.510 69.060 29.830 69.120 ;
        RECT 32.285 69.075 32.575 69.120 ;
        RECT 41.485 69.075 41.775 69.305 ;
        RECT 42.405 69.260 42.695 69.305 ;
        RECT 47.910 69.260 48.230 69.320 ;
        RECT 42.405 69.120 50.900 69.260 ;
        RECT 42.405 69.075 42.695 69.120 ;
        RECT 11.570 68.580 11.890 68.640 ;
        RECT 18.100 68.625 18.240 69.060 ;
        RECT 26.290 68.920 26.610 68.980 ;
        RECT 41.560 68.920 41.700 69.075 ;
        RECT 47.910 69.060 48.230 69.120 ;
        RECT 42.850 68.920 43.170 68.980 ;
        RECT 26.290 68.780 43.170 68.920 ;
        RECT 50.760 68.920 50.900 69.120 ;
        RECT 51.130 69.060 51.450 69.320 ;
        RECT 53.445 69.260 53.735 69.305 ;
        RECT 51.680 69.120 53.735 69.260 ;
        RECT 51.680 68.920 51.820 69.120 ;
        RECT 53.445 69.075 53.735 69.120 ;
        RECT 50.760 68.780 51.820 68.920 ;
        RECT 60.330 68.920 60.650 68.980 ;
        RECT 63.180 68.920 63.320 69.415 ;
        RECT 66.770 69.400 67.090 69.460 ;
        RECT 68.170 69.600 68.460 69.645 ;
        RECT 70.005 69.600 70.295 69.645 ;
        RECT 73.585 69.600 73.875 69.645 ;
        RECT 68.170 69.460 73.875 69.600 ;
        RECT 68.170 69.415 68.460 69.460 ;
        RECT 70.005 69.415 70.295 69.460 ;
        RECT 73.585 69.415 73.875 69.460 ;
        RECT 74.665 69.440 74.955 69.755 ;
        RECT 67.690 69.060 68.010 69.320 ;
        RECT 69.070 69.260 69.390 69.320 ;
        RECT 76.980 69.260 77.120 70.095 ;
        RECT 93.450 70.080 93.770 70.340 ;
        RECT 79.190 69.740 79.510 70.000 ;
        RECT 86.090 69.940 86.410 70.000 ;
        RECT 86.090 69.800 92.300 69.940 ;
        RECT 86.090 69.740 86.410 69.800 ;
        RECT 77.810 69.400 78.130 69.660 ;
        RECT 90.245 69.600 90.535 69.645 ;
        RECT 90.690 69.600 91.010 69.660 ;
        RECT 78.360 69.460 91.010 69.600 ;
        RECT 69.070 69.120 77.120 69.260 ;
        RECT 69.070 69.060 69.390 69.120 ;
        RECT 60.330 68.780 63.320 68.920 ;
        RECT 68.575 68.920 68.865 68.965 ;
        RECT 70.465 68.920 70.755 68.965 ;
        RECT 73.585 68.920 73.875 68.965 ;
        RECT 68.575 68.780 73.875 68.920 ;
        RECT 26.290 68.720 26.610 68.780 ;
        RECT 42.850 68.720 43.170 68.780 ;
        RECT 60.330 68.720 60.650 68.780 ;
        RECT 68.575 68.735 68.865 68.780 ;
        RECT 70.465 68.735 70.755 68.780 ;
        RECT 73.585 68.735 73.875 68.780 ;
        RECT 12.965 68.580 13.255 68.625 ;
        RECT 11.570 68.440 13.255 68.580 ;
        RECT 11.570 68.380 11.890 68.440 ;
        RECT 12.965 68.395 13.255 68.440 ;
        RECT 18.025 68.395 18.315 68.625 ;
        RECT 20.325 68.580 20.615 68.625 ;
        RECT 21.230 68.580 21.550 68.640 ;
        RECT 20.325 68.440 21.550 68.580 ;
        RECT 20.325 68.395 20.615 68.440 ;
        RECT 21.230 68.380 21.550 68.440 ;
        RECT 28.590 68.580 28.910 68.640 ;
        RECT 31.825 68.580 32.115 68.625 ;
        RECT 28.590 68.440 32.115 68.580 ;
        RECT 28.590 68.380 28.910 68.440 ;
        RECT 31.825 68.395 32.115 68.440 ;
        RECT 35.490 68.580 35.810 68.640 ;
        RECT 36.885 68.580 37.175 68.625 ;
        RECT 35.490 68.440 37.175 68.580 ;
        RECT 35.490 68.380 35.810 68.440 ;
        RECT 36.885 68.395 37.175 68.440 ;
        RECT 50.670 68.380 50.990 68.640 ;
        RECT 58.490 68.580 58.810 68.640 ;
        RECT 78.360 68.580 78.500 69.460 ;
        RECT 90.245 69.415 90.535 69.460 ;
        RECT 90.690 69.400 91.010 69.460 ;
        RECT 91.165 69.415 91.455 69.645 ;
        RECT 78.745 69.260 79.035 69.305 ;
        RECT 81.950 69.260 82.270 69.320 ;
        RECT 78.745 69.120 82.270 69.260 ;
        RECT 91.240 69.260 91.380 69.415 ;
        RECT 91.610 69.400 91.930 69.660 ;
        RECT 92.160 69.645 92.300 69.800 ;
        RECT 92.085 69.600 92.375 69.645 ;
        RECT 92.530 69.600 92.850 69.660 ;
        RECT 96.210 69.600 96.530 69.660 ;
        RECT 92.085 69.460 96.530 69.600 ;
        RECT 92.085 69.415 92.375 69.460 ;
        RECT 92.530 69.400 92.850 69.460 ;
        RECT 96.210 69.400 96.530 69.460 ;
        RECT 98.970 69.600 99.290 69.660 ;
        RECT 99.905 69.600 100.195 69.645 ;
        RECT 98.970 69.460 100.195 69.600 ;
        RECT 98.970 69.400 99.290 69.460 ;
        RECT 99.905 69.415 100.195 69.460 ;
        RECT 103.125 69.600 103.415 69.645 ;
        RECT 104.490 69.600 104.810 69.660 ;
        RECT 103.125 69.460 104.810 69.600 ;
        RECT 103.125 69.415 103.415 69.460 ;
        RECT 104.490 69.400 104.810 69.460 ;
        RECT 105.885 69.415 106.175 69.645 ;
        RECT 98.510 69.260 98.830 69.320 ;
        RECT 91.240 69.120 98.830 69.260 ;
        RECT 78.745 69.075 79.035 69.120 ;
        RECT 81.950 69.060 82.270 69.120 ;
        RECT 98.510 69.060 98.830 69.120 ;
        RECT 94.370 68.920 94.690 68.980 ;
        RECT 105.960 68.920 106.100 69.415 ;
        RECT 109.550 68.920 109.870 68.980 ;
        RECT 94.370 68.780 109.870 68.920 ;
        RECT 94.370 68.720 94.690 68.780 ;
        RECT 109.550 68.720 109.870 68.780 ;
        RECT 58.490 68.440 78.500 68.580 ;
        RECT 79.205 68.580 79.495 68.625 ;
        RECT 82.870 68.580 83.190 68.640 ;
        RECT 79.205 68.440 83.190 68.580 ;
        RECT 58.490 68.380 58.810 68.440 ;
        RECT 79.205 68.395 79.495 68.440 ;
        RECT 82.870 68.380 83.190 68.440 ;
        RECT 90.690 68.580 91.010 68.640 ;
        RECT 95.750 68.580 96.070 68.640 ;
        RECT 90.690 68.440 96.070 68.580 ;
        RECT 90.690 68.380 91.010 68.440 ;
        RECT 95.750 68.380 96.070 68.440 ;
        RECT 100.825 68.580 101.115 68.625 ;
        RECT 101.730 68.580 102.050 68.640 ;
        RECT 100.825 68.440 102.050 68.580 ;
        RECT 100.825 68.395 101.115 68.440 ;
        RECT 101.730 68.380 102.050 68.440 ;
        RECT 104.030 68.380 104.350 68.640 ;
        RECT 105.410 68.380 105.730 68.640 ;
        RECT 5.520 67.760 113.620 68.240 ;
        RECT 23.530 67.560 23.850 67.620 ;
        RECT 24.925 67.560 25.215 67.605 ;
        RECT 23.530 67.420 25.215 67.560 ;
        RECT 23.530 67.360 23.850 67.420 ;
        RECT 24.925 67.375 25.215 67.420 ;
        RECT 30.905 67.560 31.195 67.605 ;
        RECT 33.190 67.560 33.510 67.620 ;
        RECT 30.905 67.420 33.510 67.560 ;
        RECT 30.905 67.375 31.195 67.420 ;
        RECT 33.190 67.360 33.510 67.420 ;
        RECT 42.850 67.360 43.170 67.620 ;
        RECT 53.430 67.560 53.750 67.620 ;
        RECT 53.905 67.560 54.195 67.605 ;
        RECT 53.430 67.420 54.195 67.560 ;
        RECT 53.430 67.360 53.750 67.420 ;
        RECT 53.905 67.375 54.195 67.420 ;
        RECT 54.810 67.360 55.130 67.620 ;
        RECT 58.030 67.360 58.350 67.620 ;
        RECT 72.750 67.560 73.070 67.620 ;
        RECT 73.225 67.560 73.515 67.605 ;
        RECT 72.750 67.420 73.515 67.560 ;
        RECT 72.750 67.360 73.070 67.420 ;
        RECT 73.225 67.375 73.515 67.420 ;
        RECT 86.550 67.560 86.870 67.620 ;
        RECT 87.485 67.560 87.775 67.605 ;
        RECT 86.550 67.420 87.775 67.560 ;
        RECT 86.550 67.360 86.870 67.420 ;
        RECT 87.485 67.375 87.775 67.420 ;
        RECT 93.925 67.560 94.215 67.605 ;
        RECT 95.290 67.560 95.610 67.620 ;
        RECT 97.590 67.560 97.910 67.620 ;
        RECT 93.925 67.420 95.610 67.560 ;
        RECT 93.925 67.375 94.215 67.420 ;
        RECT 95.290 67.360 95.610 67.420 ;
        RECT 96.530 67.420 97.910 67.560 ;
        RECT 14.345 67.220 14.635 67.265 ;
        RECT 34.995 67.220 35.285 67.265 ;
        RECT 36.885 67.220 37.175 67.265 ;
        RECT 40.005 67.220 40.295 67.265 ;
        RECT 13.730 67.080 14.635 67.220 ;
        RECT 13.730 66.880 13.870 67.080 ;
        RECT 14.345 67.035 14.635 67.080 ;
        RECT 21.780 67.080 24.220 67.220 ;
        RECT 12.120 66.740 13.870 66.880 ;
        RECT 10.665 66.540 10.955 66.585 ;
        RECT 11.570 66.540 11.890 66.600 ;
        RECT 12.120 66.585 12.260 66.740 ;
        RECT 16.630 66.680 16.950 66.940 ;
        RECT 17.550 66.680 17.870 66.940 ;
        RECT 21.780 66.600 21.920 67.080 ;
        RECT 22.150 66.880 22.470 66.940 ;
        RECT 22.150 66.740 23.760 66.880 ;
        RECT 22.150 66.680 22.470 66.740 ;
        RECT 10.665 66.400 11.890 66.540 ;
        RECT 10.665 66.355 10.955 66.400 ;
        RECT 11.570 66.340 11.890 66.400 ;
        RECT 12.045 66.355 12.335 66.585 ;
        RECT 13.410 66.340 13.730 66.600 ;
        RECT 21.690 66.340 22.010 66.600 ;
        RECT 22.625 66.355 22.915 66.585 ;
        RECT 21.230 66.200 21.550 66.260 ;
        RECT 22.700 66.200 22.840 66.355 ;
        RECT 23.070 66.340 23.390 66.600 ;
        RECT 23.620 66.585 23.760 66.740 ;
        RECT 23.545 66.355 23.835 66.585 ;
        RECT 24.080 66.540 24.220 67.080 ;
        RECT 34.995 67.080 40.295 67.220 ;
        RECT 34.995 67.035 35.285 67.080 ;
        RECT 36.885 67.035 37.175 67.080 ;
        RECT 40.005 67.035 40.295 67.080 ;
        RECT 50.670 67.220 50.990 67.280 ;
        RECT 52.510 67.220 52.830 67.280 ;
        RECT 59.870 67.220 60.190 67.280 ;
        RECT 50.670 67.080 52.830 67.220 ;
        RECT 50.670 67.020 50.990 67.080 ;
        RECT 52.510 67.020 52.830 67.080 ;
        RECT 55.360 67.080 60.190 67.220 ;
        RECT 26.750 66.880 27.070 66.940 ;
        RECT 33.190 66.880 33.510 66.940 ;
        RECT 26.750 66.740 33.510 66.880 ;
        RECT 26.750 66.680 27.070 66.740 ;
        RECT 27.685 66.540 27.975 66.585 ;
        RECT 24.080 66.400 27.975 66.540 ;
        RECT 27.685 66.355 27.975 66.400 ;
        RECT 21.230 66.060 22.840 66.200 ;
        RECT 21.230 66.000 21.550 66.060 ;
        RECT 8.810 65.860 9.130 65.920 ;
        RECT 9.745 65.860 10.035 65.905 ;
        RECT 8.810 65.720 10.035 65.860 ;
        RECT 8.810 65.660 9.130 65.720 ;
        RECT 9.745 65.675 10.035 65.720 ;
        RECT 11.125 65.860 11.415 65.905 ;
        RECT 11.570 65.860 11.890 65.920 ;
        RECT 11.125 65.720 11.890 65.860 ;
        RECT 11.125 65.675 11.415 65.720 ;
        RECT 11.570 65.660 11.890 65.720 ;
        RECT 12.950 65.660 13.270 65.920 ;
        RECT 16.185 65.860 16.475 65.905 ;
        RECT 26.290 65.860 26.610 65.920 ;
        RECT 16.185 65.720 26.610 65.860 ;
        RECT 27.760 65.860 27.900 66.355 ;
        RECT 28.590 66.340 28.910 66.600 ;
        RECT 29.140 66.585 29.280 66.740 ;
        RECT 33.190 66.680 33.510 66.740 ;
        RECT 35.490 66.680 35.810 66.940 ;
        RECT 35.950 66.880 36.270 66.940 ;
        RECT 53.890 66.880 54.210 66.940 ;
        RECT 55.360 66.925 55.500 67.080 ;
        RECT 59.870 67.020 60.190 67.080 ;
        RECT 60.790 67.220 61.110 67.280 ;
        RECT 91.610 67.220 91.930 67.280 ;
        RECT 96.530 67.220 96.670 67.420 ;
        RECT 97.590 67.360 97.910 67.420 ;
        RECT 98.050 67.560 98.370 67.620 ;
        RECT 99.445 67.560 99.735 67.605 ;
        RECT 105.870 67.560 106.190 67.620 ;
        RECT 98.050 67.420 99.735 67.560 ;
        RECT 98.050 67.360 98.370 67.420 ;
        RECT 99.445 67.375 99.735 67.420 ;
        RECT 99.980 67.420 106.190 67.560 ;
        RECT 99.980 67.220 100.120 67.420 ;
        RECT 105.870 67.360 106.190 67.420 ;
        RECT 60.790 67.080 96.670 67.220 ;
        RECT 97.450 67.080 100.120 67.220 ;
        RECT 100.370 67.220 100.660 67.265 ;
        RECT 102.230 67.220 102.520 67.265 ;
        RECT 105.010 67.220 105.300 67.265 ;
        RECT 100.370 67.080 105.300 67.220 ;
        RECT 60.790 67.020 61.110 67.080 ;
        RECT 35.950 66.740 54.210 66.880 ;
        RECT 35.950 66.680 36.270 66.740 ;
        RECT 53.890 66.680 54.210 66.740 ;
        RECT 55.285 66.695 55.575 66.925 ;
        RECT 55.745 66.880 56.035 66.925 ;
        RECT 60.330 66.880 60.650 66.940 ;
        RECT 63.090 66.880 63.410 66.940 ;
        RECT 55.745 66.740 63.410 66.880 ;
        RECT 55.745 66.695 56.035 66.740 ;
        RECT 60.330 66.680 60.650 66.740 ;
        RECT 63.090 66.680 63.410 66.740 ;
        RECT 68.150 66.680 68.470 66.940 ;
        RECT 29.065 66.355 29.355 66.585 ;
        RECT 29.525 66.540 29.815 66.585 ;
        RECT 29.970 66.540 30.290 66.600 ;
        RECT 29.525 66.400 30.290 66.540 ;
        RECT 29.525 66.355 29.815 66.400 ;
        RECT 29.970 66.340 30.290 66.400 ;
        RECT 32.730 66.540 33.050 66.600 ;
        RECT 34.125 66.540 34.415 66.585 ;
        RECT 32.730 66.400 34.415 66.540 ;
        RECT 32.730 66.340 33.050 66.400 ;
        RECT 34.125 66.355 34.415 66.400 ;
        RECT 34.590 66.540 34.880 66.585 ;
        RECT 36.425 66.540 36.715 66.585 ;
        RECT 40.005 66.540 40.295 66.585 ;
        RECT 34.590 66.400 40.295 66.540 ;
        RECT 34.590 66.355 34.880 66.400 ;
        RECT 36.425 66.355 36.715 66.400 ;
        RECT 40.005 66.355 40.295 66.400 ;
        RECT 37.785 66.200 38.435 66.245 ;
        RECT 39.170 66.200 39.490 66.260 ;
        RECT 41.085 66.245 41.375 66.560 ;
        RECT 50.210 66.540 50.530 66.600 ;
        RECT 50.685 66.540 50.975 66.585 ;
        RECT 50.210 66.400 50.975 66.540 ;
        RECT 50.210 66.340 50.530 66.400 ;
        RECT 50.685 66.355 50.975 66.400 ;
        RECT 51.605 66.355 51.895 66.585 ;
        RECT 52.065 66.355 52.355 66.585 ;
        RECT 41.085 66.200 41.675 66.245 ;
        RECT 37.785 66.060 41.675 66.200 ;
        RECT 37.785 66.015 38.435 66.060 ;
        RECT 39.170 66.000 39.490 66.060 ;
        RECT 41.385 66.015 41.675 66.060 ;
        RECT 48.830 66.200 49.150 66.260 ;
        RECT 51.680 66.200 51.820 66.355 ;
        RECT 48.830 66.060 51.820 66.200 ;
        RECT 48.830 66.000 49.150 66.060 ;
        RECT 35.950 65.860 36.270 65.920 ;
        RECT 27.760 65.720 36.270 65.860 ;
        RECT 52.140 65.860 52.280 66.355 ;
        RECT 52.510 66.340 52.830 66.600 ;
        RECT 56.650 66.340 56.970 66.600 ;
        RECT 57.125 66.540 57.415 66.585 ;
        RECT 58.490 66.540 58.810 66.600 ;
        RECT 57.125 66.400 58.810 66.540 ;
        RECT 57.125 66.355 57.415 66.400 ;
        RECT 58.490 66.340 58.810 66.400 ;
        RECT 58.965 66.355 59.255 66.585 ;
        RECT 56.740 66.200 56.880 66.340 ;
        RECT 59.040 66.200 59.180 66.355 ;
        RECT 59.410 66.340 59.730 66.600 ;
        RECT 67.230 66.540 67.550 66.600 ;
        RECT 72.765 66.540 73.055 66.585 ;
        RECT 67.230 66.400 73.055 66.540 ;
        RECT 67.230 66.340 67.550 66.400 ;
        RECT 72.765 66.355 73.055 66.400 ;
        RECT 82.870 66.540 83.190 66.600 ;
        RECT 85.720 66.585 85.860 67.080 ;
        RECT 91.610 67.020 91.930 67.080 ;
        RECT 97.450 66.880 97.590 67.080 ;
        RECT 100.370 67.035 100.660 67.080 ;
        RECT 102.230 67.035 102.520 67.080 ;
        RECT 105.010 67.035 105.300 67.080 ;
        RECT 93.080 66.740 97.590 66.880 ;
        RECT 84.265 66.540 84.555 66.585 ;
        RECT 85.080 66.540 85.370 66.585 ;
        RECT 82.870 66.400 84.555 66.540 ;
        RECT 82.870 66.340 83.190 66.400 ;
        RECT 84.265 66.355 84.555 66.400 ;
        RECT 84.800 66.400 85.370 66.540 ;
        RECT 56.740 66.060 59.180 66.200 ;
        RECT 83.790 66.200 84.110 66.260 ;
        RECT 84.800 66.200 84.940 66.400 ;
        RECT 85.080 66.355 85.370 66.400 ;
        RECT 85.645 66.355 85.935 66.585 ;
        RECT 86.090 66.340 86.410 66.600 ;
        RECT 90.690 66.340 91.010 66.600 ;
        RECT 91.610 66.340 91.930 66.600 ;
        RECT 92.085 66.355 92.375 66.585 ;
        RECT 83.790 66.060 84.940 66.200 ;
        RECT 91.150 66.200 91.470 66.260 ;
        RECT 92.160 66.200 92.300 66.355 ;
        RECT 92.530 66.340 92.850 66.600 ;
        RECT 91.150 66.060 92.300 66.200 ;
        RECT 83.790 66.000 84.110 66.060 ;
        RECT 91.150 66.000 91.470 66.060 ;
        RECT 52.510 65.860 52.830 65.920 ;
        RECT 52.140 65.720 52.830 65.860 ;
        RECT 16.185 65.675 16.475 65.720 ;
        RECT 26.290 65.660 26.610 65.720 ;
        RECT 35.950 65.660 36.270 65.720 ;
        RECT 52.510 65.660 52.830 65.720 ;
        RECT 64.010 65.860 64.330 65.920 ;
        RECT 85.630 65.860 85.950 65.920 ;
        RECT 64.010 65.720 85.950 65.860 ;
        RECT 64.010 65.660 64.330 65.720 ;
        RECT 85.630 65.660 85.950 65.720 ;
        RECT 91.610 65.860 91.930 65.920 ;
        RECT 93.080 65.860 93.220 66.740 ;
        RECT 101.730 66.680 102.050 66.940 ;
        RECT 94.370 66.340 94.690 66.600 ;
        RECT 95.750 66.540 96.070 66.600 ;
        RECT 96.225 66.540 96.515 66.585 ;
        RECT 95.750 66.400 96.515 66.540 ;
        RECT 95.750 66.340 96.070 66.400 ;
        RECT 96.225 66.355 96.515 66.400 ;
        RECT 96.670 66.540 96.990 66.600 ;
        RECT 97.145 66.540 97.435 66.585 ;
        RECT 96.670 66.400 97.435 66.540 ;
        RECT 96.670 66.340 96.990 66.400 ;
        RECT 97.145 66.355 97.435 66.400 ;
        RECT 97.590 66.340 97.910 66.600 ;
        RECT 98.065 66.355 98.355 66.585 ;
        RECT 98.140 66.200 98.280 66.355 ;
        RECT 99.890 66.340 100.210 66.600 ;
        RECT 105.010 66.540 105.300 66.585 ;
        RECT 102.765 66.400 105.300 66.540 ;
        RECT 102.765 66.245 102.980 66.400 ;
        RECT 105.010 66.355 105.300 66.400 ;
        RECT 109.550 66.340 109.870 66.600 ;
        RECT 97.680 66.060 98.280 66.200 ;
        RECT 100.830 66.200 101.120 66.245 ;
        RECT 102.690 66.200 102.980 66.245 ;
        RECT 100.830 66.060 102.980 66.200 ;
        RECT 91.610 65.720 93.220 65.860 ;
        RECT 94.845 65.860 95.135 65.905 ;
        RECT 95.290 65.860 95.610 65.920 ;
        RECT 94.845 65.720 95.610 65.860 ;
        RECT 91.610 65.660 91.930 65.720 ;
        RECT 94.845 65.675 95.135 65.720 ;
        RECT 95.290 65.660 95.610 65.720 ;
        RECT 96.210 65.860 96.530 65.920 ;
        RECT 97.680 65.860 97.820 66.060 ;
        RECT 100.830 66.015 101.120 66.060 ;
        RECT 102.690 66.015 102.980 66.060 ;
        RECT 103.610 66.200 103.900 66.245 ;
        RECT 105.410 66.200 105.730 66.260 ;
        RECT 106.870 66.200 107.160 66.245 ;
        RECT 103.610 66.060 107.160 66.200 ;
        RECT 103.610 66.015 103.900 66.060 ;
        RECT 105.410 66.000 105.730 66.060 ;
        RECT 106.870 66.015 107.160 66.060 ;
        RECT 96.210 65.720 97.820 65.860 ;
        RECT 103.110 65.860 103.430 65.920 ;
        RECT 108.875 65.860 109.165 65.905 ;
        RECT 103.110 65.720 109.165 65.860 ;
        RECT 96.210 65.660 96.530 65.720 ;
        RECT 103.110 65.660 103.430 65.720 ;
        RECT 108.875 65.675 109.165 65.720 ;
        RECT 110.010 65.660 110.330 65.920 ;
        RECT 5.520 65.040 113.620 65.520 ;
        RECT 15.250 64.840 15.570 64.900 ;
        RECT 15.955 64.840 16.245 64.885 ;
        RECT 15.250 64.700 16.245 64.840 ;
        RECT 15.250 64.640 15.570 64.700 ;
        RECT 15.955 64.655 16.245 64.700 ;
        RECT 20.770 64.640 21.090 64.900 ;
        RECT 21.690 64.840 22.010 64.900 ;
        RECT 24.450 64.840 24.770 64.900 ;
        RECT 21.690 64.700 24.770 64.840 ;
        RECT 21.690 64.640 22.010 64.700 ;
        RECT 24.450 64.640 24.770 64.700 ;
        RECT 27.670 64.640 27.990 64.900 ;
        RECT 31.825 64.840 32.115 64.885 ;
        RECT 33.650 64.840 33.970 64.900 ;
        RECT 31.825 64.700 33.970 64.840 ;
        RECT 31.825 64.655 32.115 64.700 ;
        RECT 33.650 64.640 33.970 64.700 ;
        RECT 39.170 64.840 39.490 64.900 ;
        RECT 39.645 64.840 39.935 64.885 ;
        RECT 39.170 64.700 39.935 64.840 ;
        RECT 39.170 64.640 39.490 64.700 ;
        RECT 39.645 64.655 39.935 64.700 ;
        RECT 50.685 64.840 50.975 64.885 ;
        RECT 51.590 64.840 51.910 64.900 ;
        RECT 64.485 64.840 64.775 64.885 ;
        RECT 50.685 64.700 51.910 64.840 ;
        RECT 50.685 64.655 50.975 64.700 ;
        RECT 51.590 64.640 51.910 64.700 ;
        RECT 53.980 64.700 64.775 64.840 ;
        RECT 7.910 64.500 8.200 64.545 ;
        RECT 9.770 64.500 10.060 64.545 ;
        RECT 7.910 64.360 10.060 64.500 ;
        RECT 7.910 64.315 8.200 64.360 ;
        RECT 9.770 64.315 10.060 64.360 ;
        RECT 10.690 64.500 10.980 64.545 ;
        RECT 12.950 64.500 13.270 64.560 ;
        RECT 13.950 64.500 14.240 64.545 ;
        RECT 50.210 64.500 50.530 64.560 ;
        RECT 53.980 64.500 54.120 64.700 ;
        RECT 64.485 64.655 64.775 64.700 ;
        RECT 73.685 64.840 73.975 64.885 ;
        RECT 77.810 64.840 78.130 64.900 ;
        RECT 73.685 64.700 78.130 64.840 ;
        RECT 73.685 64.655 73.975 64.700 ;
        RECT 64.560 64.500 64.700 64.655 ;
        RECT 77.810 64.640 78.130 64.700 ;
        RECT 83.330 64.640 83.650 64.900 ;
        RECT 98.970 64.840 99.290 64.900 ;
        RECT 99.890 64.840 100.210 64.900 ;
        RECT 89.860 64.700 100.210 64.840 ;
        RECT 68.610 64.500 68.930 64.560 ;
        RECT 77.350 64.500 77.670 64.560 ;
        RECT 10.690 64.360 14.240 64.500 ;
        RECT 10.690 64.315 10.980 64.360 ;
        RECT 8.810 63.960 9.130 64.220 ;
        RECT 9.845 64.160 10.060 64.315 ;
        RECT 12.950 64.300 13.270 64.360 ;
        RECT 13.950 64.315 14.240 64.360 ;
        RECT 17.640 64.360 39.400 64.500 ;
        RECT 12.090 64.160 12.380 64.205 ;
        RECT 9.845 64.020 12.380 64.160 ;
        RECT 12.090 63.975 12.380 64.020 ;
        RECT 13.410 64.160 13.730 64.220 ;
        RECT 17.640 64.205 17.780 64.360 ;
        RECT 17.565 64.160 17.855 64.205 ;
        RECT 13.410 64.020 17.855 64.160 ;
        RECT 13.410 63.960 13.730 64.020 ;
        RECT 17.565 63.975 17.855 64.020 ;
        RECT 22.165 63.975 22.455 64.205 ;
        RECT 22.625 63.975 22.915 64.205 ;
        RECT 6.985 63.820 7.275 63.865 ;
        RECT 7.890 63.820 8.210 63.880 ;
        RECT 6.985 63.680 8.210 63.820 ;
        RECT 6.985 63.635 7.275 63.680 ;
        RECT 7.890 63.620 8.210 63.680 ;
        RECT 7.450 63.480 7.740 63.525 ;
        RECT 9.310 63.480 9.600 63.525 ;
        RECT 12.090 63.480 12.380 63.525 ;
        RECT 7.450 63.340 12.380 63.480 ;
        RECT 7.450 63.295 7.740 63.340 ;
        RECT 9.310 63.295 9.600 63.340 ;
        RECT 12.090 63.295 12.380 63.340 ;
        RECT 22.240 63.200 22.380 63.975 ;
        RECT 22.700 63.820 22.840 63.975 ;
        RECT 23.070 63.960 23.390 64.220 ;
        RECT 24.005 64.160 24.295 64.205 ;
        RECT 24.450 64.160 24.770 64.220 ;
        RECT 24.005 64.020 24.770 64.160 ;
        RECT 24.005 63.975 24.295 64.020 ;
        RECT 24.450 63.960 24.770 64.020 ;
        RECT 25.385 63.975 25.675 64.205 ;
        RECT 25.460 63.820 25.600 63.975 ;
        RECT 25.830 63.960 26.150 64.220 ;
        RECT 26.305 64.160 26.595 64.205 ;
        RECT 29.970 64.160 30.290 64.220 ;
        RECT 33.205 64.160 33.495 64.205 ;
        RECT 26.305 64.020 33.495 64.160 ;
        RECT 26.305 63.975 26.595 64.020 ;
        RECT 26.750 63.820 27.070 63.880 ;
        RECT 22.700 63.680 23.760 63.820 ;
        RECT 25.460 63.680 27.070 63.820 ;
        RECT 23.620 63.540 23.760 63.680 ;
        RECT 26.750 63.620 27.070 63.680 ;
        RECT 23.530 63.480 23.850 63.540 ;
        RECT 25.830 63.480 26.150 63.540 ;
        RECT 23.530 63.340 26.150 63.480 ;
        RECT 23.530 63.280 23.850 63.340 ;
        RECT 25.830 63.280 26.150 63.340 ;
        RECT 17.090 62.940 17.410 63.200 ;
        RECT 22.150 63.140 22.470 63.200 ;
        RECT 27.300 63.140 27.440 64.020 ;
        RECT 29.970 63.960 30.290 64.020 ;
        RECT 33.205 63.975 33.495 64.020 ;
        RECT 33.280 63.820 33.420 63.975 ;
        RECT 33.650 63.960 33.970 64.220 ;
        RECT 34.110 63.960 34.430 64.220 ;
        RECT 35.045 64.160 35.335 64.205 ;
        RECT 35.950 64.160 36.270 64.220 ;
        RECT 39.260 64.205 39.400 64.360 ;
        RECT 50.210 64.360 54.120 64.500 ;
        RECT 50.210 64.300 50.530 64.360 ;
        RECT 53.980 64.220 54.120 64.360 ;
        RECT 59.500 64.360 61.940 64.500 ;
        RECT 64.560 64.360 68.380 64.500 ;
        RECT 35.045 64.020 36.270 64.160 ;
        RECT 35.045 63.975 35.335 64.020 ;
        RECT 35.950 63.960 36.270 64.020 ;
        RECT 39.185 64.160 39.475 64.205 ;
        RECT 43.770 64.160 44.090 64.220 ;
        RECT 39.185 64.020 44.090 64.160 ;
        RECT 39.185 63.975 39.475 64.020 ;
        RECT 43.770 63.960 44.090 64.020 ;
        RECT 50.670 64.160 50.990 64.220 ;
        RECT 52.065 64.160 52.355 64.205 ;
        RECT 50.670 64.020 52.355 64.160 ;
        RECT 50.670 63.960 50.990 64.020 ;
        RECT 52.065 63.975 52.355 64.020 ;
        RECT 52.510 63.960 52.830 64.220 ;
        RECT 52.985 64.160 53.275 64.205 ;
        RECT 53.430 64.160 53.750 64.220 ;
        RECT 52.985 64.020 53.750 64.160 ;
        RECT 52.985 63.975 53.275 64.020 ;
        RECT 53.430 63.960 53.750 64.020 ;
        RECT 53.890 63.960 54.210 64.220 ;
        RECT 56.665 64.160 56.955 64.205 ;
        RECT 57.110 64.160 57.430 64.220 ;
        RECT 56.665 64.020 57.430 64.160 ;
        RECT 56.665 63.975 56.955 64.020 ;
        RECT 57.110 63.960 57.430 64.020 ;
        RECT 58.490 64.160 58.810 64.220 ;
        RECT 59.500 64.205 59.640 64.360 ;
        RECT 59.425 64.160 59.715 64.205 ;
        RECT 58.490 64.020 59.715 64.160 ;
        RECT 58.490 63.960 58.810 64.020 ;
        RECT 59.425 63.975 59.715 64.020 ;
        RECT 59.870 63.960 60.190 64.220 ;
        RECT 61.800 64.205 61.940 64.360 ;
        RECT 61.725 63.975 62.015 64.205 ;
        RECT 63.565 63.975 63.855 64.205 ;
        RECT 51.590 63.820 51.910 63.880 ;
        RECT 52.600 63.820 52.740 63.960 ;
        RECT 33.280 63.680 33.880 63.820 ;
        RECT 33.740 63.480 33.880 63.680 ;
        RECT 51.590 63.680 52.740 63.820 ;
        RECT 54.350 63.820 54.670 63.880 ;
        RECT 58.030 63.820 58.350 63.880 ;
        RECT 59.960 63.820 60.100 63.960 ;
        RECT 63.640 63.820 63.780 63.975 ;
        RECT 66.310 63.960 66.630 64.220 ;
        RECT 68.240 64.160 68.380 64.360 ;
        RECT 68.610 64.360 85.400 64.500 ;
        RECT 68.610 64.300 68.930 64.360 ;
        RECT 70.465 64.160 70.755 64.205 ;
        RECT 68.240 64.020 70.755 64.160 ;
        RECT 70.465 63.975 70.755 64.020 ;
        RECT 54.350 63.680 59.640 63.820 ;
        RECT 59.960 63.680 63.780 63.820 ;
        RECT 70.540 63.820 70.680 63.975 ;
        RECT 71.370 63.960 71.690 64.220 ;
        RECT 71.920 64.205 72.060 64.360 ;
        RECT 77.350 64.300 77.670 64.360 ;
        RECT 71.845 63.975 72.135 64.205 ;
        RECT 72.290 63.960 72.610 64.220 ;
        RECT 81.030 64.160 81.350 64.220 ;
        RECT 85.260 64.205 85.400 64.360 ;
        RECT 84.725 64.160 85.015 64.205 ;
        RECT 81.030 64.020 85.015 64.160 ;
        RECT 81.030 63.960 81.350 64.020 ;
        RECT 84.725 63.975 85.015 64.020 ;
        RECT 85.185 63.975 85.475 64.205 ;
        RECT 85.630 63.960 85.950 64.220 ;
        RECT 86.550 63.960 86.870 64.220 ;
        RECT 89.860 64.205 90.000 64.700 ;
        RECT 98.970 64.640 99.290 64.700 ;
        RECT 99.890 64.640 100.210 64.700 ;
        RECT 103.585 64.840 103.875 64.885 ;
        RECT 104.490 64.840 104.810 64.900 ;
        RECT 103.585 64.700 104.810 64.840 ;
        RECT 103.585 64.655 103.875 64.700 ;
        RECT 104.490 64.640 104.810 64.700 ;
        RECT 105.870 64.640 106.190 64.900 ;
        RECT 90.710 64.500 91.000 64.545 ;
        RECT 92.570 64.500 92.860 64.545 ;
        RECT 90.710 64.360 92.860 64.500 ;
        RECT 90.710 64.315 91.000 64.360 ;
        RECT 92.570 64.315 92.860 64.360 ;
        RECT 93.490 64.500 93.780 64.545 ;
        RECT 95.290 64.500 95.610 64.560 ;
        RECT 96.750 64.500 97.040 64.545 ;
        RECT 93.490 64.360 97.040 64.500 ;
        RECT 93.490 64.315 93.780 64.360 ;
        RECT 88.405 63.975 88.695 64.205 ;
        RECT 89.785 63.975 90.075 64.205 ;
        RECT 92.645 64.160 92.860 64.315 ;
        RECT 95.290 64.300 95.610 64.360 ;
        RECT 96.750 64.315 97.040 64.360 ;
        RECT 98.510 64.500 98.830 64.560 ;
        RECT 101.745 64.500 102.035 64.545 ;
        RECT 103.110 64.500 103.430 64.560 ;
        RECT 105.425 64.500 105.715 64.545 ;
        RECT 98.510 64.360 105.715 64.500 ;
        RECT 98.510 64.300 98.830 64.360 ;
        RECT 101.745 64.315 102.035 64.360 ;
        RECT 103.110 64.300 103.430 64.360 ;
        RECT 105.425 64.315 105.715 64.360 ;
        RECT 94.890 64.160 95.180 64.205 ;
        RECT 92.645 64.020 95.180 64.160 ;
        RECT 94.890 63.975 95.180 64.020 ;
        RECT 101.285 63.975 101.575 64.205 ;
        RECT 75.970 63.820 76.290 63.880 ;
        RECT 70.540 63.680 76.290 63.820 ;
        RECT 51.590 63.620 51.910 63.680 ;
        RECT 54.350 63.620 54.670 63.680 ;
        RECT 58.030 63.620 58.350 63.680 ;
        RECT 52.510 63.480 52.830 63.540 ;
        RECT 33.740 63.340 52.830 63.480 ;
        RECT 52.510 63.280 52.830 63.340 ;
        RECT 58.505 63.480 58.795 63.525 ;
        RECT 58.950 63.480 59.270 63.540 ;
        RECT 58.505 63.340 59.270 63.480 ;
        RECT 59.500 63.480 59.640 63.680 ;
        RECT 75.970 63.620 76.290 63.680 ;
        RECT 60.805 63.480 61.095 63.525 ;
        RECT 59.500 63.340 61.095 63.480 ;
        RECT 58.505 63.295 58.795 63.340 ;
        RECT 58.950 63.280 59.270 63.340 ;
        RECT 60.805 63.295 61.095 63.340 ;
        RECT 62.170 63.480 62.490 63.540 ;
        RECT 65.405 63.480 65.695 63.525 ;
        RECT 62.170 63.340 65.695 63.480 ;
        RECT 62.170 63.280 62.490 63.340 ;
        RECT 65.405 63.295 65.695 63.340 ;
        RECT 22.150 63.000 27.440 63.140 ;
        RECT 33.650 63.140 33.970 63.200 ;
        RECT 55.270 63.140 55.590 63.200 ;
        RECT 33.650 63.000 55.590 63.140 ;
        RECT 22.150 62.940 22.470 63.000 ;
        RECT 33.650 62.940 33.970 63.000 ;
        RECT 55.270 62.940 55.590 63.000 ;
        RECT 55.730 62.940 56.050 63.200 ;
        RECT 62.645 63.140 62.935 63.185 ;
        RECT 64.470 63.140 64.790 63.200 ;
        RECT 78.270 63.140 78.590 63.200 ;
        RECT 62.645 63.000 78.590 63.140 ;
        RECT 88.480 63.140 88.620 63.975 ;
        RECT 91.625 63.820 91.915 63.865 ;
        RECT 89.400 63.680 91.915 63.820 ;
        RECT 89.400 63.525 89.540 63.680 ;
        RECT 91.625 63.635 91.915 63.680 ;
        RECT 92.990 63.820 93.310 63.880 ;
        RECT 98.755 63.820 99.045 63.865 ;
        RECT 101.360 63.820 101.500 63.975 ;
        RECT 92.990 63.680 101.500 63.820 ;
        RECT 92.990 63.620 93.310 63.680 ;
        RECT 98.755 63.635 99.045 63.680 ;
        RECT 102.665 63.635 102.955 63.865 ;
        RECT 106.345 63.635 106.635 63.865 ;
        RECT 89.325 63.295 89.615 63.525 ;
        RECT 90.250 63.480 90.540 63.525 ;
        RECT 92.110 63.480 92.400 63.525 ;
        RECT 94.890 63.480 95.180 63.525 ;
        RECT 90.250 63.340 95.180 63.480 ;
        RECT 90.250 63.295 90.540 63.340 ;
        RECT 92.110 63.295 92.400 63.340 ;
        RECT 94.890 63.295 95.180 63.340 ;
        RECT 99.430 63.280 99.750 63.540 ;
        RECT 102.190 63.480 102.510 63.540 ;
        RECT 102.740 63.480 102.880 63.635 ;
        RECT 106.420 63.480 106.560 63.635 ;
        RECT 102.190 63.340 106.560 63.480 ;
        RECT 102.190 63.280 102.510 63.340 ;
        RECT 89.770 63.140 90.090 63.200 ;
        RECT 88.480 63.000 90.090 63.140 ;
        RECT 62.645 62.955 62.935 63.000 ;
        RECT 64.470 62.940 64.790 63.000 ;
        RECT 78.270 62.940 78.590 63.000 ;
        RECT 89.770 62.940 90.090 63.000 ;
        RECT 5.520 62.320 113.620 62.800 ;
        RECT 16.630 61.920 16.950 62.180 ;
        RECT 24.465 62.120 24.755 62.165 ;
        RECT 27.210 62.120 27.530 62.180 ;
        RECT 24.465 61.980 27.530 62.120 ;
        RECT 24.465 61.935 24.755 61.980 ;
        RECT 27.210 61.920 27.530 61.980 ;
        RECT 52.970 62.120 53.290 62.180 ;
        RECT 54.365 62.120 54.655 62.165 ;
        RECT 52.970 61.980 54.655 62.120 ;
        RECT 52.970 61.920 53.290 61.980 ;
        RECT 54.365 61.935 54.655 61.980 ;
        RECT 55.270 62.120 55.590 62.180 ;
        RECT 60.790 62.120 61.110 62.180 ;
        RECT 55.270 61.980 61.110 62.120 ;
        RECT 55.270 61.920 55.590 61.980 ;
        RECT 60.790 61.920 61.110 61.980 ;
        RECT 64.485 62.120 64.775 62.165 ;
        RECT 66.310 62.120 66.630 62.180 ;
        RECT 64.485 61.980 66.630 62.120 ;
        RECT 64.485 61.935 64.775 61.980 ;
        RECT 66.310 61.920 66.630 61.980 ;
        RECT 79.205 62.120 79.495 62.165 ;
        RECT 79.650 62.120 79.970 62.180 ;
        RECT 79.205 61.980 79.970 62.120 ;
        RECT 79.205 61.935 79.495 61.980 ;
        RECT 79.650 61.920 79.970 61.980 ;
        RECT 83.790 62.120 84.110 62.180 ;
        RECT 90.230 62.120 90.550 62.180 ;
        RECT 90.705 62.120 90.995 62.165 ;
        RECT 83.790 61.980 90.000 62.120 ;
        RECT 83.790 61.920 84.110 61.980 ;
        RECT 8.775 61.780 9.065 61.825 ;
        RECT 10.665 61.780 10.955 61.825 ;
        RECT 13.785 61.780 14.075 61.825 ;
        RECT 8.775 61.640 14.075 61.780 ;
        RECT 8.775 61.595 9.065 61.640 ;
        RECT 10.665 61.595 10.955 61.640 ;
        RECT 13.785 61.595 14.075 61.640 ;
        RECT 45.170 61.780 45.460 61.825 ;
        RECT 47.030 61.780 47.320 61.825 ;
        RECT 49.810 61.780 50.100 61.825 ;
        RECT 45.170 61.640 50.100 61.780 ;
        RECT 45.170 61.595 45.460 61.640 ;
        RECT 47.030 61.595 47.320 61.640 ;
        RECT 49.810 61.595 50.100 61.640 ;
        RECT 53.890 61.780 54.210 61.840 ;
        RECT 75.970 61.780 76.290 61.840 ;
        RECT 82.870 61.780 83.190 61.840 ;
        RECT 86.550 61.780 86.870 61.840 ;
        RECT 53.890 61.640 57.340 61.780 ;
        RECT 53.890 61.580 54.210 61.640 ;
        RECT 9.285 61.440 9.575 61.485 ;
        RECT 11.570 61.440 11.890 61.500 ;
        RECT 23.530 61.440 23.850 61.500 ;
        RECT 9.285 61.300 11.890 61.440 ;
        RECT 9.285 61.255 9.575 61.300 ;
        RECT 11.570 61.240 11.890 61.300 ;
        RECT 22.700 61.300 23.850 61.440 ;
        RECT 7.890 60.900 8.210 61.160 ;
        RECT 8.370 61.100 8.660 61.145 ;
        RECT 10.205 61.100 10.495 61.145 ;
        RECT 13.785 61.100 14.075 61.145 ;
        RECT 8.370 60.960 14.075 61.100 ;
        RECT 8.370 60.915 8.660 60.960 ;
        RECT 10.205 60.915 10.495 60.960 ;
        RECT 13.785 60.915 14.075 60.960 ;
        RECT 14.865 60.805 15.155 61.120 ;
        RECT 21.245 61.100 21.535 61.145 ;
        RECT 21.690 61.100 22.010 61.160 ;
        RECT 22.700 61.145 22.840 61.300 ;
        RECT 23.530 61.240 23.850 61.300 ;
        RECT 51.590 61.440 51.910 61.500 ;
        RECT 51.590 61.300 56.420 61.440 ;
        RECT 51.590 61.240 51.910 61.300 ;
        RECT 21.245 60.960 22.010 61.100 ;
        RECT 21.245 60.915 21.535 60.960 ;
        RECT 21.690 60.900 22.010 60.960 ;
        RECT 22.165 60.915 22.455 61.145 ;
        RECT 22.625 60.915 22.915 61.145 ;
        RECT 23.085 60.915 23.375 61.145 ;
        RECT 11.565 60.760 12.215 60.805 ;
        RECT 14.865 60.760 15.455 60.805 ;
        RECT 17.090 60.760 17.410 60.820 ;
        RECT 11.565 60.620 17.410 60.760 ;
        RECT 11.565 60.575 12.215 60.620 ;
        RECT 15.165 60.575 15.455 60.620 ;
        RECT 17.090 60.560 17.410 60.620 ;
        RECT 17.550 60.760 17.870 60.820 ;
        RECT 22.240 60.760 22.380 60.915 ;
        RECT 17.550 60.620 22.380 60.760 ;
        RECT 17.550 60.560 17.870 60.620 ;
        RECT 22.150 60.420 22.470 60.480 ;
        RECT 23.160 60.420 23.300 60.915 ;
        RECT 44.690 60.900 45.010 61.160 ;
        RECT 46.545 61.100 46.835 61.145 ;
        RECT 49.810 61.100 50.100 61.145 ;
        RECT 45.240 60.960 46.835 61.100 ;
        RECT 43.310 60.760 43.630 60.820 ;
        RECT 45.240 60.760 45.380 60.960 ;
        RECT 46.545 60.915 46.835 60.960 ;
        RECT 47.565 60.960 50.100 61.100 ;
        RECT 47.565 60.805 47.780 60.960 ;
        RECT 49.810 60.915 50.100 60.960 ;
        RECT 50.670 61.100 50.990 61.160 ;
        RECT 56.280 61.145 56.420 61.300 ;
        RECT 55.745 61.100 56.035 61.145 ;
        RECT 50.670 60.960 56.035 61.100 ;
        RECT 50.670 60.900 50.990 60.960 ;
        RECT 55.745 60.915 56.035 60.960 ;
        RECT 56.205 60.915 56.495 61.145 ;
        RECT 56.665 60.915 56.955 61.145 ;
        RECT 57.200 61.100 57.340 61.640 ;
        RECT 75.970 61.640 86.870 61.780 ;
        RECT 75.970 61.580 76.290 61.640 ;
        RECT 82.870 61.580 83.190 61.640 ;
        RECT 86.550 61.580 86.870 61.640 ;
        RECT 64.470 61.440 64.790 61.500 ;
        RECT 67.245 61.440 67.535 61.485 ;
        RECT 72.290 61.440 72.610 61.500 ;
        RECT 79.665 61.440 79.955 61.485 ;
        RECT 80.110 61.440 80.430 61.500 ;
        RECT 64.470 61.300 67.535 61.440 ;
        RECT 64.470 61.240 64.790 61.300 ;
        RECT 67.245 61.255 67.535 61.300 ;
        RECT 68.240 61.300 78.040 61.440 ;
        RECT 57.585 61.100 57.875 61.145 ;
        RECT 57.200 60.960 57.875 61.100 ;
        RECT 57.585 60.915 57.875 60.960 ;
        RECT 59.410 61.100 59.730 61.160 ;
        RECT 59.885 61.100 60.175 61.145 ;
        RECT 59.410 60.960 60.175 61.100 ;
        RECT 43.310 60.620 45.380 60.760 ;
        RECT 45.630 60.760 45.920 60.805 ;
        RECT 47.490 60.760 47.780 60.805 ;
        RECT 48.410 60.760 48.700 60.805 ;
        RECT 51.670 60.760 51.960 60.805 ;
        RECT 45.630 60.620 47.780 60.760 ;
        RECT 43.310 60.560 43.630 60.620 ;
        RECT 45.630 60.575 45.920 60.620 ;
        RECT 47.490 60.575 47.780 60.620 ;
        RECT 48.000 60.620 51.960 60.760 ;
        RECT 22.150 60.280 23.300 60.420 ;
        RECT 44.230 60.420 44.550 60.480 ;
        RECT 48.000 60.420 48.140 60.620 ;
        RECT 48.410 60.575 48.700 60.620 ;
        RECT 51.670 60.575 51.960 60.620 ;
        RECT 44.230 60.280 48.140 60.420 ;
        RECT 48.830 60.420 49.150 60.480 ;
        RECT 53.675 60.420 53.965 60.465 ;
        RECT 48.830 60.280 53.965 60.420 ;
        RECT 55.820 60.420 55.960 60.915 ;
        RECT 56.740 60.760 56.880 60.915 ;
        RECT 59.410 60.900 59.730 60.960 ;
        RECT 59.885 60.915 60.175 60.960 ;
        RECT 61.710 60.900 62.030 61.160 ;
        RECT 68.240 61.100 68.380 61.300 ;
        RECT 72.290 61.240 72.610 61.300 ;
        RECT 62.720 60.960 68.380 61.100 ;
        RECT 68.625 61.100 68.915 61.145 ;
        RECT 69.530 61.100 69.850 61.160 ;
        RECT 68.625 60.960 69.850 61.100 ;
        RECT 58.030 60.760 58.350 60.820 ;
        RECT 56.740 60.620 58.350 60.760 ;
        RECT 58.030 60.560 58.350 60.620 ;
        RECT 62.720 60.465 62.860 60.960 ;
        RECT 68.625 60.915 68.915 60.960 ;
        RECT 69.530 60.900 69.850 60.960 ;
        RECT 75.970 60.900 76.290 61.160 ;
        RECT 76.890 60.900 77.210 61.160 ;
        RECT 77.350 60.900 77.670 61.160 ;
        RECT 77.900 61.145 78.040 61.300 ;
        RECT 79.665 61.300 80.430 61.440 ;
        RECT 79.665 61.255 79.955 61.300 ;
        RECT 80.110 61.240 80.430 61.300 ;
        RECT 77.825 61.100 78.115 61.145 ;
        RECT 77.825 61.085 80.800 61.100 ;
        RECT 81.030 61.085 81.350 61.160 ;
        RECT 77.825 60.960 81.350 61.085 ;
        RECT 77.825 60.915 78.115 60.960 ;
        RECT 80.660 60.945 81.350 60.960 ;
        RECT 81.030 60.900 81.350 60.945 ;
        RECT 81.505 60.915 81.795 61.145 ;
        RECT 81.965 61.100 82.255 61.145 ;
        RECT 82.410 61.100 82.730 61.160 ;
        RECT 82.960 61.145 83.100 61.580 ;
        RECT 83.330 61.240 83.650 61.500 ;
        RECT 81.965 60.960 82.730 61.100 ;
        RECT 81.965 60.915 82.255 60.960 ;
        RECT 66.785 60.760 67.075 60.805 ;
        RECT 71.370 60.760 71.690 60.820 ;
        RECT 66.785 60.620 71.690 60.760 ;
        RECT 77.440 60.760 77.580 60.900 ;
        RECT 81.580 60.760 81.720 60.915 ;
        RECT 82.410 60.900 82.730 60.960 ;
        RECT 82.885 60.915 83.175 61.145 ;
        RECT 83.790 61.100 84.110 61.160 ;
        RECT 84.495 61.100 84.785 61.145 ;
        RECT 83.790 60.960 84.785 61.100 ;
        RECT 83.790 60.900 84.110 60.960 ;
        RECT 84.495 60.915 84.785 60.960 ;
        RECT 85.185 60.915 85.475 61.145 ;
        RECT 85.645 61.100 85.935 61.145 ;
        RECT 86.090 61.100 86.410 61.160 ;
        RECT 86.640 61.145 86.780 61.580 ;
        RECT 89.860 61.440 90.000 61.980 ;
        RECT 90.230 61.980 90.995 62.120 ;
        RECT 90.230 61.920 90.550 61.980 ;
        RECT 90.705 61.935 90.995 61.980 ;
        RECT 96.670 62.120 96.990 62.180 ;
        RECT 97.590 62.120 97.910 62.180 ;
        RECT 96.670 61.980 97.910 62.120 ;
        RECT 96.670 61.920 96.990 61.980 ;
        RECT 97.590 61.920 97.910 61.980 ;
        RECT 105.870 62.120 106.190 62.180 ;
        RECT 111.175 62.120 111.465 62.165 ;
        RECT 105.870 61.980 111.465 62.120 ;
        RECT 105.870 61.920 106.190 61.980 ;
        RECT 111.175 61.935 111.465 61.980 ;
        RECT 102.190 61.580 102.510 61.840 ;
        RECT 102.670 61.780 102.960 61.825 ;
        RECT 104.530 61.780 104.820 61.825 ;
        RECT 107.310 61.780 107.600 61.825 ;
        RECT 102.670 61.640 107.600 61.780 ;
        RECT 102.670 61.595 102.960 61.640 ;
        RECT 104.530 61.595 104.820 61.640 ;
        RECT 107.310 61.595 107.600 61.640 ;
        RECT 92.990 61.440 93.310 61.500 ;
        RECT 89.860 61.300 93.310 61.440 ;
        RECT 92.990 61.240 93.310 61.300 ;
        RECT 93.925 61.440 94.215 61.485 ;
        RECT 96.670 61.440 96.990 61.500 ;
        RECT 102.280 61.440 102.420 61.580 ;
        RECT 93.925 61.300 102.420 61.440 ;
        RECT 93.925 61.255 94.215 61.300 ;
        RECT 96.670 61.240 96.990 61.300 ;
        RECT 104.030 61.240 104.350 61.500 ;
        RECT 85.645 60.960 86.410 61.100 ;
        RECT 85.645 60.915 85.935 60.960 ;
        RECT 83.330 60.760 83.650 60.820 ;
        RECT 77.440 60.620 83.650 60.760 ;
        RECT 66.785 60.575 67.075 60.620 ;
        RECT 71.370 60.560 71.690 60.620 ;
        RECT 83.330 60.560 83.650 60.620 ;
        RECT 62.645 60.420 62.935 60.465 ;
        RECT 55.820 60.280 62.935 60.420 ;
        RECT 22.150 60.220 22.470 60.280 ;
        RECT 44.230 60.220 44.550 60.280 ;
        RECT 48.830 60.220 49.150 60.280 ;
        RECT 53.675 60.235 53.965 60.280 ;
        RECT 62.645 60.235 62.935 60.280 ;
        RECT 66.325 60.420 66.615 60.465 ;
        RECT 69.070 60.420 69.390 60.480 ;
        RECT 66.325 60.280 69.390 60.420 ;
        RECT 66.325 60.235 66.615 60.280 ;
        RECT 69.070 60.220 69.390 60.280 ;
        RECT 69.545 60.420 69.835 60.465 ;
        RECT 71.830 60.420 72.150 60.480 ;
        RECT 69.545 60.280 72.150 60.420 ;
        RECT 83.420 60.420 83.560 60.560 ;
        RECT 85.260 60.420 85.400 60.915 ;
        RECT 86.090 60.900 86.410 60.960 ;
        RECT 86.565 60.915 86.855 61.145 ;
        RECT 98.970 61.100 99.290 61.160 ;
        RECT 102.205 61.100 102.495 61.145 ;
        RECT 107.310 61.100 107.600 61.145 ;
        RECT 98.970 60.960 102.495 61.100 ;
        RECT 98.970 60.900 99.290 60.960 ;
        RECT 102.205 60.915 102.495 60.960 ;
        RECT 105.065 60.960 107.600 61.100 ;
        RECT 105.065 60.805 105.280 60.960 ;
        RECT 107.310 60.915 107.600 60.960 ;
        RECT 103.130 60.760 103.420 60.805 ;
        RECT 104.990 60.760 105.280 60.805 ;
        RECT 103.130 60.620 105.280 60.760 ;
        RECT 103.130 60.575 103.420 60.620 ;
        RECT 104.990 60.575 105.280 60.620 ;
        RECT 105.910 60.760 106.200 60.805 ;
        RECT 109.170 60.760 109.460 60.805 ;
        RECT 110.010 60.760 110.330 60.820 ;
        RECT 105.910 60.620 110.330 60.760 ;
        RECT 105.910 60.575 106.200 60.620 ;
        RECT 109.170 60.575 109.460 60.620 ;
        RECT 110.010 60.560 110.330 60.620 ;
        RECT 83.420 60.280 85.400 60.420 ;
        RECT 85.630 60.420 85.950 60.480 ;
        RECT 92.530 60.420 92.850 60.480 ;
        RECT 85.630 60.280 92.850 60.420 ;
        RECT 69.545 60.235 69.835 60.280 ;
        RECT 71.830 60.220 72.150 60.280 ;
        RECT 85.630 60.220 85.950 60.280 ;
        RECT 92.530 60.220 92.850 60.280 ;
        RECT 5.520 59.600 113.620 60.080 ;
        RECT 26.750 59.400 27.070 59.460 ;
        RECT 28.145 59.400 28.435 59.445 ;
        RECT 26.750 59.260 28.435 59.400 ;
        RECT 26.750 59.200 27.070 59.260 ;
        RECT 28.145 59.215 28.435 59.260 ;
        RECT 28.605 59.400 28.895 59.445 ;
        RECT 34.110 59.400 34.430 59.460 ;
        RECT 36.425 59.400 36.715 59.445 ;
        RECT 28.605 59.260 36.715 59.400 ;
        RECT 28.605 59.215 28.895 59.260 ;
        RECT 34.110 59.200 34.430 59.260 ;
        RECT 36.425 59.215 36.715 59.260 ;
        RECT 43.310 59.200 43.630 59.460 ;
        RECT 44.230 59.200 44.550 59.460 ;
        RECT 45.165 59.215 45.455 59.445 ;
        RECT 47.465 59.400 47.755 59.445 ;
        RECT 48.830 59.400 49.150 59.460 ;
        RECT 47.465 59.260 49.150 59.400 ;
        RECT 47.465 59.215 47.755 59.260 ;
        RECT 14.805 59.060 15.095 59.105 ;
        RECT 15.250 59.060 15.570 59.120 ;
        RECT 45.240 59.060 45.380 59.215 ;
        RECT 48.830 59.200 49.150 59.260 ;
        RECT 49.290 59.400 49.610 59.460 ;
        RECT 49.765 59.400 50.055 59.445 ;
        RECT 49.290 59.260 50.055 59.400 ;
        RECT 49.290 59.200 49.610 59.260 ;
        RECT 49.765 59.215 50.055 59.260 ;
        RECT 54.350 59.400 54.670 59.460 ;
        RECT 58.030 59.400 58.350 59.460 ;
        RECT 54.350 59.260 58.350 59.400 ;
        RECT 54.350 59.200 54.670 59.260 ;
        RECT 58.030 59.200 58.350 59.260 ;
        RECT 58.965 59.400 59.255 59.445 ;
        RECT 68.610 59.400 68.930 59.460 ;
        RECT 58.965 59.260 68.930 59.400 ;
        RECT 58.965 59.215 59.255 59.260 ;
        RECT 14.805 58.920 15.570 59.060 ;
        RECT 14.805 58.875 15.095 58.920 ;
        RECT 15.250 58.860 15.570 58.920 ;
        RECT 42.480 58.920 45.380 59.060 ;
        RECT 50.670 59.060 50.990 59.120 ;
        RECT 59.040 59.060 59.180 59.215 ;
        RECT 68.610 59.200 68.930 59.260 ;
        RECT 69.085 59.215 69.375 59.445 ;
        RECT 50.670 58.920 51.360 59.060 ;
        RECT 16.170 58.520 16.490 58.780 ;
        RECT 42.480 58.765 42.620 58.920 ;
        RECT 50.670 58.860 50.990 58.920 ;
        RECT 29.140 58.580 37.560 58.720 ;
        RECT 22.150 58.380 22.470 58.440 ;
        RECT 29.140 58.425 29.280 58.580 ;
        RECT 29.065 58.380 29.355 58.425 ;
        RECT 22.150 58.240 29.355 58.380 ;
        RECT 22.150 58.180 22.470 58.240 ;
        RECT 29.065 58.195 29.355 58.240 ;
        RECT 36.870 58.180 37.190 58.440 ;
        RECT 37.420 58.425 37.560 58.580 ;
        RECT 42.405 58.535 42.695 58.765 ;
        RECT 43.770 58.520 44.090 58.780 ;
        RECT 46.990 58.720 47.310 58.780 ;
        RECT 51.220 58.765 51.360 58.920 ;
        RECT 51.680 58.920 59.180 59.060 ;
        RECT 61.725 59.060 62.015 59.105 ;
        RECT 62.170 59.060 62.490 59.120 ;
        RECT 61.725 58.920 62.490 59.060 ;
        RECT 51.680 58.780 51.820 58.920 ;
        RECT 61.725 58.875 62.015 58.920 ;
        RECT 62.170 58.860 62.490 58.920 ;
        RECT 64.005 59.060 64.655 59.105 ;
        RECT 65.390 59.060 65.710 59.120 ;
        RECT 67.605 59.060 67.895 59.105 ;
        RECT 64.005 58.920 67.895 59.060 ;
        RECT 69.160 59.060 69.300 59.215 ;
        RECT 69.530 59.200 69.850 59.460 ;
        RECT 71.370 59.400 71.690 59.460 ;
        RECT 70.080 59.260 71.690 59.400 ;
        RECT 70.080 59.060 70.220 59.260 ;
        RECT 71.370 59.200 71.690 59.260 ;
        RECT 86.565 59.400 86.855 59.445 ;
        RECT 87.010 59.400 87.330 59.460 ;
        RECT 86.565 59.260 87.330 59.400 ;
        RECT 86.565 59.215 86.855 59.260 ;
        RECT 87.010 59.200 87.330 59.260 ;
        RECT 102.665 59.400 102.955 59.445 ;
        RECT 105.870 59.400 106.190 59.460 ;
        RECT 102.665 59.260 106.190 59.400 ;
        RECT 102.665 59.215 102.955 59.260 ;
        RECT 105.870 59.200 106.190 59.260 ;
        RECT 69.160 58.920 70.220 59.060 ;
        RECT 73.670 59.060 73.990 59.120 ;
        RECT 75.525 59.060 75.815 59.105 ;
        RECT 73.670 58.920 75.815 59.060 ;
        RECT 64.005 58.875 64.655 58.920 ;
        RECT 65.390 58.860 65.710 58.920 ;
        RECT 67.305 58.875 67.895 58.920 ;
        RECT 46.990 58.580 50.900 58.720 ;
        RECT 46.990 58.520 47.310 58.580 ;
        RECT 37.345 58.380 37.635 58.425 ;
        RECT 47.925 58.380 48.215 58.425 ;
        RECT 49.750 58.380 50.070 58.440 ;
        RECT 37.345 58.240 50.070 58.380 ;
        RECT 50.760 58.380 50.900 58.580 ;
        RECT 51.145 58.535 51.435 58.765 ;
        RECT 51.590 58.520 51.910 58.780 ;
        RECT 52.065 58.535 52.355 58.765 ;
        RECT 52.985 58.720 53.275 58.765 ;
        RECT 53.890 58.720 54.210 58.780 ;
        RECT 52.985 58.580 54.210 58.720 ;
        RECT 52.985 58.535 53.275 58.580 ;
        RECT 52.140 58.380 52.280 58.535 ;
        RECT 53.890 58.520 54.210 58.580 ;
        RECT 59.410 58.720 59.730 58.780 ;
        RECT 59.885 58.720 60.175 58.765 ;
        RECT 59.410 58.580 60.175 58.720 ;
        RECT 59.410 58.520 59.730 58.580 ;
        RECT 59.885 58.535 60.175 58.580 ;
        RECT 60.810 58.720 61.100 58.765 ;
        RECT 62.645 58.720 62.935 58.765 ;
        RECT 66.225 58.720 66.515 58.765 ;
        RECT 60.810 58.580 66.515 58.720 ;
        RECT 60.810 58.535 61.100 58.580 ;
        RECT 62.645 58.535 62.935 58.580 ;
        RECT 66.225 58.535 66.515 58.580 ;
        RECT 67.305 58.560 67.595 58.875 ;
        RECT 73.670 58.860 73.990 58.920 ;
        RECT 75.525 58.875 75.815 58.920 ;
        RECT 81.030 59.060 81.350 59.120 ;
        RECT 83.790 59.060 84.110 59.120 ;
        RECT 81.030 58.920 85.400 59.060 ;
        RECT 81.030 58.860 81.350 58.920 ;
        RECT 83.790 58.860 84.110 58.920 ;
        RECT 71.845 58.720 72.135 58.765 ;
        RECT 75.985 58.720 76.275 58.765 ;
        RECT 76.890 58.720 77.210 58.780 ;
        RECT 79.190 58.720 79.510 58.780 ;
        RECT 71.845 58.580 79.510 58.720 ;
        RECT 71.845 58.535 72.135 58.580 ;
        RECT 75.985 58.535 76.275 58.580 ;
        RECT 76.890 58.520 77.210 58.580 ;
        RECT 79.190 58.520 79.510 58.580 ;
        RECT 82.870 58.720 83.190 58.780 ;
        RECT 83.345 58.720 83.635 58.765 ;
        RECT 82.870 58.580 83.635 58.720 ;
        RECT 82.870 58.520 83.190 58.580 ;
        RECT 83.345 58.535 83.635 58.580 ;
        RECT 84.265 58.535 84.555 58.765 ;
        RECT 50.760 58.240 52.280 58.380 ;
        RECT 37.345 58.195 37.635 58.240 ;
        RECT 47.925 58.195 48.215 58.240 ;
        RECT 49.750 58.180 50.070 58.240 ;
        RECT 60.345 58.195 60.635 58.425 ;
        RECT 64.470 58.380 64.790 58.440 ;
        RECT 72.305 58.380 72.595 58.425 ;
        RECT 74.590 58.380 74.910 58.440 ;
        RECT 64.470 58.240 74.910 58.380 ;
        RECT 84.340 58.380 84.480 58.535 ;
        RECT 84.710 58.520 85.030 58.780 ;
        RECT 85.260 58.765 85.400 58.920 ;
        RECT 85.185 58.535 85.475 58.765 ;
        RECT 102.190 58.720 102.510 58.780 ;
        RECT 105.885 58.720 106.175 58.765 ;
        RECT 109.550 58.720 109.870 58.780 ;
        RECT 102.190 58.580 103.800 58.720 ;
        RECT 102.190 58.520 102.510 58.580 ;
        RECT 103.110 58.380 103.430 58.440 ;
        RECT 103.660 58.425 103.800 58.580 ;
        RECT 105.885 58.580 109.870 58.720 ;
        RECT 105.885 58.535 106.175 58.580 ;
        RECT 109.550 58.520 109.870 58.580 ;
        RECT 84.340 58.240 103.430 58.380 ;
        RECT 26.305 57.700 26.595 57.745 ;
        RECT 28.130 57.700 28.450 57.760 ;
        RECT 26.305 57.560 28.450 57.700 ;
        RECT 26.305 57.515 26.595 57.560 ;
        RECT 28.130 57.500 28.450 57.560 ;
        RECT 34.585 57.700 34.875 57.745 ;
        RECT 35.490 57.700 35.810 57.760 ;
        RECT 34.585 57.560 35.810 57.700 ;
        RECT 60.420 57.700 60.560 58.195 ;
        RECT 64.470 58.180 64.790 58.240 ;
        RECT 72.305 58.195 72.595 58.240 ;
        RECT 74.590 58.180 74.910 58.240 ;
        RECT 103.110 58.180 103.430 58.240 ;
        RECT 103.585 58.195 103.875 58.425 ;
        RECT 61.215 58.040 61.505 58.085 ;
        RECT 63.105 58.040 63.395 58.085 ;
        RECT 66.225 58.040 66.515 58.085 ;
        RECT 97.590 58.040 97.910 58.100 ;
        RECT 61.215 57.900 66.515 58.040 ;
        RECT 61.215 57.855 61.505 57.900 ;
        RECT 63.105 57.855 63.395 57.900 ;
        RECT 66.225 57.855 66.515 57.900 ;
        RECT 77.440 57.900 97.910 58.040 ;
        RECT 67.690 57.700 68.010 57.760 ;
        RECT 68.610 57.700 68.930 57.760 ;
        RECT 60.420 57.560 68.930 57.700 ;
        RECT 34.585 57.515 34.875 57.560 ;
        RECT 35.490 57.500 35.810 57.560 ;
        RECT 67.690 57.500 68.010 57.560 ;
        RECT 68.610 57.500 68.930 57.560 ;
        RECT 69.070 57.700 69.390 57.760 ;
        RECT 77.440 57.700 77.580 57.900 ;
        RECT 97.590 57.840 97.910 57.900 ;
        RECT 69.070 57.560 77.580 57.700 ;
        RECT 77.825 57.700 78.115 57.745 ;
        RECT 80.570 57.700 80.890 57.760 ;
        RECT 77.825 57.560 80.890 57.700 ;
        RECT 69.070 57.500 69.390 57.560 ;
        RECT 77.825 57.515 78.115 57.560 ;
        RECT 80.570 57.500 80.890 57.560 ;
        RECT 98.510 57.700 98.830 57.760 ;
        RECT 100.825 57.700 101.115 57.745 ;
        RECT 98.510 57.560 101.115 57.700 ;
        RECT 98.510 57.500 98.830 57.560 ;
        RECT 100.825 57.515 101.115 57.560 ;
        RECT 105.410 57.500 105.730 57.760 ;
        RECT 5.520 56.880 113.620 57.360 ;
        RECT 32.055 56.680 32.345 56.725 ;
        RECT 34.110 56.680 34.430 56.740 ;
        RECT 32.055 56.540 34.430 56.680 ;
        RECT 32.055 56.495 32.345 56.540 ;
        RECT 34.110 56.480 34.430 56.540 ;
        RECT 36.870 56.680 37.190 56.740 ;
        RECT 41.715 56.680 42.005 56.725 ;
        RECT 46.990 56.680 47.310 56.740 ;
        RECT 36.870 56.540 47.310 56.680 ;
        RECT 36.870 56.480 37.190 56.540 ;
        RECT 41.715 56.495 42.005 56.540 ;
        RECT 46.990 56.480 47.310 56.540 ;
        RECT 52.510 56.680 52.830 56.740 ;
        RECT 60.805 56.680 61.095 56.725 ;
        RECT 64.010 56.680 64.330 56.740 ;
        RECT 52.510 56.540 64.330 56.680 ;
        RECT 52.510 56.480 52.830 56.540 ;
        RECT 60.805 56.495 61.095 56.540 ;
        RECT 64.010 56.480 64.330 56.540 ;
        RECT 65.390 56.480 65.710 56.740 ;
        RECT 79.190 56.480 79.510 56.740 ;
        RECT 96.670 56.680 96.990 56.740 ;
        RECT 81.580 56.540 90.000 56.680 ;
        RECT 18.945 56.155 19.235 56.385 ;
        RECT 23.550 56.340 23.840 56.385 ;
        RECT 25.410 56.340 25.700 56.385 ;
        RECT 28.190 56.340 28.480 56.385 ;
        RECT 23.550 56.200 28.480 56.340 ;
        RECT 23.550 56.155 23.840 56.200 ;
        RECT 25.410 56.155 25.700 56.200 ;
        RECT 28.190 56.155 28.480 56.200 ;
        RECT 33.210 56.340 33.500 56.385 ;
        RECT 35.070 56.340 35.360 56.385 ;
        RECT 37.850 56.340 38.140 56.385 ;
        RECT 33.210 56.200 38.140 56.340 ;
        RECT 33.210 56.155 33.500 56.200 ;
        RECT 35.070 56.155 35.360 56.200 ;
        RECT 37.850 56.155 38.140 56.200 ;
        RECT 48.385 56.155 48.675 56.385 ;
        RECT 71.335 56.340 71.625 56.385 ;
        RECT 73.225 56.340 73.515 56.385 ;
        RECT 76.345 56.340 76.635 56.385 ;
        RECT 71.335 56.200 76.635 56.340 ;
        RECT 71.335 56.155 71.625 56.200 ;
        RECT 73.225 56.155 73.515 56.200 ;
        RECT 76.345 56.155 76.635 56.200 ;
        RECT 13.410 56.000 13.730 56.060 ;
        RECT 13.885 56.000 14.175 56.045 ;
        RECT 13.410 55.860 14.175 56.000 ;
        RECT 13.410 55.800 13.730 55.860 ;
        RECT 13.885 55.815 14.175 55.860 ;
        RECT 12.045 55.475 12.335 55.705 ;
        RECT 12.950 55.660 13.270 55.720 ;
        RECT 16.170 55.660 16.490 55.720 ;
        RECT 17.105 55.660 17.395 55.705 ;
        RECT 19.020 55.660 19.160 56.155 ;
        RECT 22.150 55.800 22.470 56.060 ;
        RECT 24.925 56.000 25.215 56.045 ;
        RECT 27.210 56.000 27.530 56.060 ;
        RECT 24.925 55.860 27.530 56.000 ;
        RECT 24.925 55.815 25.215 55.860 ;
        RECT 27.210 55.800 27.530 55.860 ;
        RECT 32.730 55.800 33.050 56.060 ;
        RECT 12.950 55.520 16.860 55.660 ;
        RECT 12.120 55.320 12.260 55.475 ;
        RECT 12.950 55.460 13.270 55.520 ;
        RECT 16.170 55.460 16.490 55.520 ;
        RECT 13.870 55.320 14.190 55.380 ;
        RECT 12.120 55.180 14.190 55.320 ;
        RECT 16.720 55.320 16.860 55.520 ;
        RECT 17.105 55.520 19.160 55.660 ;
        RECT 20.770 55.660 21.090 55.720 ;
        RECT 23.085 55.660 23.375 55.705 ;
        RECT 28.190 55.660 28.480 55.705 ;
        RECT 20.770 55.520 23.375 55.660 ;
        RECT 17.105 55.475 17.395 55.520 ;
        RECT 20.770 55.460 21.090 55.520 ;
        RECT 23.085 55.475 23.375 55.520 ;
        RECT 25.945 55.520 28.480 55.660 ;
        RECT 19.390 55.320 19.710 55.380 ;
        RECT 21.690 55.320 22.010 55.380 ;
        RECT 25.945 55.365 26.160 55.520 ;
        RECT 28.190 55.475 28.480 55.520 ;
        RECT 34.570 55.460 34.890 55.720 ;
        RECT 37.850 55.660 38.140 55.705 ;
        RECT 35.605 55.520 38.140 55.660 ;
        RECT 29.970 55.365 30.290 55.380 ;
        RECT 35.605 55.365 35.820 55.520 ;
        RECT 37.850 55.475 38.140 55.520 ;
        RECT 47.925 55.660 48.215 55.705 ;
        RECT 48.460 55.660 48.600 56.155 ;
        RECT 49.750 56.000 50.070 56.060 ;
        RECT 51.145 56.000 51.435 56.045 ;
        RECT 52.970 56.000 53.290 56.060 ;
        RECT 55.285 56.000 55.575 56.045 ;
        RECT 49.750 55.860 55.575 56.000 ;
        RECT 49.750 55.800 50.070 55.860 ;
        RECT 51.145 55.815 51.435 55.860 ;
        RECT 52.970 55.800 53.290 55.860 ;
        RECT 55.285 55.815 55.575 55.860 ;
        RECT 67.230 55.800 67.550 56.060 ;
        RECT 68.610 56.000 68.930 56.060 ;
        RECT 70.465 56.000 70.755 56.045 ;
        RECT 72.290 56.000 72.610 56.060 ;
        RECT 68.610 55.860 72.610 56.000 ;
        RECT 68.610 55.800 68.930 55.860 ;
        RECT 70.465 55.815 70.755 55.860 ;
        RECT 72.290 55.800 72.610 55.860 ;
        RECT 74.590 56.000 74.910 56.060 ;
        RECT 81.580 56.045 81.720 56.540 ;
        RECT 84.725 56.155 85.015 56.385 ;
        RECT 89.325 56.155 89.615 56.385 ;
        RECT 81.505 56.000 81.795 56.045 ;
        RECT 74.590 55.860 81.795 56.000 ;
        RECT 74.590 55.800 74.910 55.860 ;
        RECT 81.505 55.815 81.795 55.860 ;
        RECT 47.925 55.520 48.600 55.660 ;
        RECT 48.830 55.660 49.150 55.720 ;
        RECT 50.225 55.660 50.515 55.705 ;
        RECT 48.830 55.520 50.515 55.660 ;
        RECT 47.925 55.475 48.215 55.520 ;
        RECT 48.830 55.460 49.150 55.520 ;
        RECT 50.225 55.475 50.515 55.520 ;
        RECT 50.685 55.660 50.975 55.705 ;
        RECT 54.350 55.660 54.670 55.720 ;
        RECT 50.685 55.520 54.670 55.660 ;
        RECT 50.685 55.475 50.975 55.520 ;
        RECT 54.350 55.460 54.670 55.520 ;
        RECT 59.870 55.660 60.190 55.720 ;
        RECT 61.710 55.660 62.030 55.720 ;
        RECT 59.870 55.520 62.030 55.660 ;
        RECT 59.870 55.460 60.190 55.520 ;
        RECT 61.710 55.460 62.030 55.520 ;
        RECT 65.850 55.460 66.170 55.720 ;
        RECT 66.310 55.460 66.630 55.720 ;
        RECT 70.930 55.660 71.220 55.705 ;
        RECT 72.765 55.660 73.055 55.705 ;
        RECT 76.345 55.660 76.635 55.705 ;
        RECT 70.930 55.520 76.635 55.660 ;
        RECT 70.930 55.475 71.220 55.520 ;
        RECT 72.765 55.475 73.055 55.520 ;
        RECT 76.345 55.475 76.635 55.520 ;
        RECT 16.720 55.180 19.710 55.320 ;
        RECT 13.870 55.120 14.190 55.180 ;
        RECT 19.390 55.120 19.710 55.180 ;
        RECT 20.860 55.180 22.010 55.320 ;
        RECT 11.110 54.780 11.430 55.040 ;
        RECT 18.010 54.780 18.330 55.040 ;
        RECT 20.860 55.025 21.000 55.180 ;
        RECT 21.690 55.120 22.010 55.180 ;
        RECT 24.010 55.320 24.300 55.365 ;
        RECT 25.870 55.320 26.160 55.365 ;
        RECT 24.010 55.180 26.160 55.320 ;
        RECT 24.010 55.135 24.300 55.180 ;
        RECT 25.870 55.135 26.160 55.180 ;
        RECT 26.790 55.320 27.080 55.365 ;
        RECT 29.970 55.320 30.340 55.365 ;
        RECT 26.790 55.180 30.340 55.320 ;
        RECT 26.790 55.135 27.080 55.180 ;
        RECT 29.970 55.135 30.340 55.180 ;
        RECT 33.670 55.320 33.960 55.365 ;
        RECT 35.530 55.320 35.820 55.365 ;
        RECT 33.670 55.180 35.820 55.320 ;
        RECT 33.670 55.135 33.960 55.180 ;
        RECT 35.530 55.135 35.820 55.180 ;
        RECT 36.450 55.320 36.740 55.365 ;
        RECT 37.330 55.320 37.650 55.380 ;
        RECT 39.710 55.320 40.000 55.365 ;
        RECT 36.450 55.180 40.000 55.320 ;
        RECT 36.450 55.135 36.740 55.180 ;
        RECT 29.970 55.120 30.290 55.135 ;
        RECT 37.330 55.120 37.650 55.180 ;
        RECT 39.710 55.135 40.000 55.180 ;
        RECT 71.830 55.120 72.150 55.380 ;
        RECT 74.590 55.365 74.910 55.380 ;
        RECT 74.125 55.320 74.910 55.365 ;
        RECT 77.425 55.365 77.715 55.680 ;
        RECT 80.570 55.460 80.890 55.720 ;
        RECT 82.410 55.460 82.730 55.720 ;
        RECT 84.800 55.660 84.940 56.155 ;
        RECT 86.105 55.660 86.395 55.705 ;
        RECT 84.800 55.520 86.395 55.660 ;
        RECT 86.105 55.475 86.395 55.520 ;
        RECT 86.550 55.460 86.870 55.720 ;
        RECT 88.865 55.660 89.155 55.705 ;
        RECT 89.400 55.660 89.540 56.155 ;
        RECT 89.860 56.000 90.000 56.540 ;
        RECT 92.160 56.540 96.990 56.680 ;
        RECT 92.160 56.045 92.300 56.540 ;
        RECT 96.670 56.480 96.990 56.540 ;
        RECT 103.110 56.680 103.430 56.740 ;
        RECT 108.875 56.680 109.165 56.725 ;
        RECT 103.110 56.540 109.165 56.680 ;
        RECT 103.110 56.480 103.430 56.540 ;
        RECT 108.875 56.495 109.165 56.540 ;
        RECT 99.445 56.155 99.735 56.385 ;
        RECT 100.370 56.340 100.660 56.385 ;
        RECT 102.230 56.340 102.520 56.385 ;
        RECT 105.010 56.340 105.300 56.385 ;
        RECT 100.370 56.200 105.300 56.340 ;
        RECT 100.370 56.155 100.660 56.200 ;
        RECT 102.230 56.155 102.520 56.200 ;
        RECT 105.010 56.155 105.300 56.200 ;
        RECT 92.085 56.000 92.375 56.045 ;
        RECT 89.860 55.860 92.375 56.000 ;
        RECT 99.520 56.000 99.660 56.155 ;
        RECT 101.745 56.000 102.035 56.045 ;
        RECT 99.520 55.860 102.035 56.000 ;
        RECT 92.085 55.815 92.375 55.860 ;
        RECT 101.745 55.815 102.035 55.860 ;
        RECT 88.865 55.520 89.540 55.660 ;
        RECT 88.865 55.475 89.155 55.520 ;
        RECT 97.130 55.460 97.450 55.720 ;
        RECT 98.510 55.460 98.830 55.720 ;
        RECT 98.970 55.660 99.290 55.720 ;
        RECT 99.905 55.660 100.195 55.705 ;
        RECT 105.010 55.660 105.300 55.705 ;
        RECT 98.970 55.520 100.195 55.660 ;
        RECT 98.970 55.460 99.290 55.520 ;
        RECT 99.905 55.475 100.195 55.520 ;
        RECT 102.765 55.520 105.300 55.660 ;
        RECT 77.425 55.320 78.015 55.365 ;
        RECT 82.500 55.320 82.640 55.460 ;
        RECT 82.885 55.320 83.175 55.365 ;
        RECT 86.640 55.320 86.780 55.460 ;
        RECT 102.765 55.365 102.980 55.520 ;
        RECT 105.010 55.475 105.300 55.520 ;
        RECT 109.550 55.460 109.870 55.720 ;
        RECT 100.830 55.320 101.120 55.365 ;
        RECT 102.690 55.320 102.980 55.365 ;
        RECT 74.125 55.180 78.015 55.320 ;
        RECT 74.125 55.135 74.910 55.180 ;
        RECT 77.725 55.135 78.015 55.180 ;
        RECT 78.360 55.180 83.175 55.320 ;
        RECT 74.590 55.120 74.910 55.135 ;
        RECT 20.785 54.795 21.075 55.025 ;
        RECT 21.245 54.980 21.535 55.025 ;
        RECT 26.290 54.980 26.610 55.040 ;
        RECT 21.245 54.840 26.610 54.980 ;
        RECT 21.245 54.795 21.535 54.840 ;
        RECT 26.290 54.780 26.610 54.840 ;
        RECT 46.990 54.780 47.310 55.040 ;
        RECT 52.510 54.780 52.830 55.040 ;
        RECT 53.430 54.980 53.750 55.040 ;
        RECT 54.825 54.980 55.115 55.025 ;
        RECT 53.430 54.840 55.115 54.980 ;
        RECT 53.430 54.780 53.750 54.840 ;
        RECT 54.825 54.795 55.115 54.840 ;
        RECT 58.030 54.980 58.350 55.040 ;
        RECT 58.950 54.980 59.270 55.040 ;
        RECT 58.030 54.840 59.270 54.980 ;
        RECT 58.030 54.780 58.350 54.840 ;
        RECT 58.950 54.780 59.270 54.840 ;
        RECT 73.670 54.980 73.990 55.040 ;
        RECT 78.360 54.980 78.500 55.180 ;
        RECT 82.885 55.135 83.175 55.180 ;
        RECT 84.800 55.180 91.380 55.320 ;
        RECT 73.670 54.840 78.500 54.980 ;
        RECT 73.670 54.780 73.990 54.840 ;
        RECT 79.650 54.780 79.970 55.040 ;
        RECT 82.425 54.980 82.715 55.025 ;
        RECT 84.800 54.980 84.940 55.180 ;
        RECT 91.240 55.040 91.380 55.180 ;
        RECT 100.830 55.180 102.980 55.320 ;
        RECT 100.830 55.135 101.120 55.180 ;
        RECT 102.690 55.135 102.980 55.180 ;
        RECT 103.610 55.320 103.900 55.365 ;
        RECT 105.410 55.320 105.730 55.380 ;
        RECT 106.870 55.320 107.160 55.365 ;
        RECT 103.610 55.180 107.160 55.320 ;
        RECT 103.610 55.135 103.900 55.180 ;
        RECT 105.410 55.120 105.730 55.180 ;
        RECT 106.870 55.135 107.160 55.180 ;
        RECT 82.425 54.840 84.940 54.980 ;
        RECT 85.185 54.980 85.475 55.025 ;
        RECT 86.550 54.980 86.870 55.040 ;
        RECT 85.185 54.840 86.870 54.980 ;
        RECT 82.425 54.795 82.715 54.840 ;
        RECT 85.185 54.795 85.475 54.840 ;
        RECT 86.550 54.780 86.870 54.840 ;
        RECT 87.930 54.780 88.250 55.040 ;
        RECT 91.150 54.780 91.470 55.040 ;
        RECT 91.625 54.980 91.915 55.025 ;
        RECT 92.530 54.980 92.850 55.040 ;
        RECT 94.370 54.980 94.690 55.040 ;
        RECT 91.625 54.840 94.690 54.980 ;
        RECT 91.625 54.795 91.915 54.840 ;
        RECT 92.530 54.780 92.850 54.840 ;
        RECT 94.370 54.780 94.690 54.840 ;
        RECT 98.050 54.780 98.370 55.040 ;
        RECT 110.010 54.780 110.330 55.040 ;
        RECT 5.520 54.160 113.620 54.640 ;
        RECT 21.230 53.960 21.550 54.020 ;
        RECT 17.640 53.820 21.550 53.960 ;
        RECT 9.745 53.620 10.035 53.665 ;
        RECT 11.110 53.620 11.430 53.680 ;
        RECT 9.745 53.480 11.430 53.620 ;
        RECT 9.745 53.435 10.035 53.480 ;
        RECT 11.110 53.420 11.430 53.480 ;
        RECT 12.025 53.620 12.675 53.665 ;
        RECT 15.625 53.620 15.915 53.665 ;
        RECT 17.090 53.620 17.410 53.680 ;
        RECT 12.025 53.480 17.410 53.620 ;
        RECT 12.025 53.435 12.675 53.480 ;
        RECT 15.325 53.435 15.915 53.480 ;
        RECT 8.830 53.280 9.120 53.325 ;
        RECT 10.665 53.280 10.955 53.325 ;
        RECT 14.245 53.280 14.535 53.325 ;
        RECT 8.830 53.140 14.535 53.280 ;
        RECT 8.830 53.095 9.120 53.140 ;
        RECT 10.665 53.095 10.955 53.140 ;
        RECT 14.245 53.095 14.535 53.140 ;
        RECT 15.325 53.120 15.615 53.435 ;
        RECT 17.090 53.420 17.410 53.480 ;
        RECT 7.890 52.940 8.210 53.000 ;
        RECT 8.365 52.940 8.655 52.985 ;
        RECT 17.105 52.940 17.395 52.985 ;
        RECT 17.640 52.940 17.780 53.820 ;
        RECT 21.230 53.760 21.550 53.820 ;
        RECT 26.750 53.760 27.070 54.020 ;
        RECT 27.210 53.760 27.530 54.020 ;
        RECT 29.970 53.960 30.290 54.020 ;
        RECT 32.285 53.960 32.575 54.005 ;
        RECT 29.970 53.820 32.575 53.960 ;
        RECT 29.970 53.760 30.290 53.820 ;
        RECT 32.285 53.775 32.575 53.820 ;
        RECT 34.570 53.760 34.890 54.020 ;
        RECT 37.330 53.960 37.650 54.020 ;
        RECT 53.890 54.005 54.210 54.020 ;
        RECT 37.805 53.960 38.095 54.005 ;
        RECT 37.330 53.820 38.095 53.960 ;
        RECT 37.330 53.760 37.650 53.820 ;
        RECT 37.805 53.775 38.095 53.820 ;
        RECT 43.785 53.960 44.075 54.005 ;
        RECT 43.785 53.820 48.140 53.960 ;
        RECT 43.785 53.775 44.075 53.820 ;
        RECT 18.010 53.620 18.330 53.680 ;
        RECT 19.405 53.620 19.695 53.665 ;
        RECT 18.010 53.480 19.695 53.620 ;
        RECT 18.010 53.420 18.330 53.480 ;
        RECT 19.405 53.435 19.695 53.480 ;
        RECT 21.685 53.620 22.335 53.665 ;
        RECT 25.285 53.620 25.575 53.665 ;
        RECT 29.065 53.620 29.355 53.665 ;
        RECT 21.685 53.480 29.355 53.620 ;
        RECT 21.685 53.435 22.335 53.480 ;
        RECT 24.985 53.435 25.575 53.480 ;
        RECT 29.065 53.435 29.355 53.480 ;
        RECT 45.630 53.620 45.920 53.665 ;
        RECT 47.490 53.620 47.780 53.665 ;
        RECT 45.630 53.480 47.780 53.620 ;
        RECT 48.000 53.620 48.140 53.820 ;
        RECT 53.675 53.775 54.210 54.005 ;
        RECT 71.385 53.960 71.675 54.005 ;
        RECT 74.590 53.960 74.910 54.020 ;
        RECT 71.385 53.820 74.910 53.960 ;
        RECT 71.385 53.775 71.675 53.820 ;
        RECT 53.890 53.760 54.210 53.775 ;
        RECT 74.590 53.760 74.910 53.820 ;
        RECT 91.150 53.960 91.470 54.020 ;
        RECT 92.085 53.960 92.375 54.005 ;
        RECT 91.150 53.820 92.375 53.960 ;
        RECT 91.150 53.760 91.470 53.820 ;
        RECT 92.085 53.775 92.375 53.820 ;
        RECT 48.410 53.620 48.700 53.665 ;
        RECT 51.670 53.620 51.960 53.665 ;
        RECT 48.000 53.480 51.960 53.620 ;
        RECT 45.630 53.435 45.920 53.480 ;
        RECT 47.490 53.435 47.780 53.480 ;
        RECT 48.410 53.435 48.700 53.480 ;
        RECT 51.670 53.435 51.960 53.480 ;
        RECT 52.970 53.620 53.290 53.680 ;
        RECT 54.365 53.620 54.655 53.665 ;
        RECT 52.970 53.480 54.655 53.620 ;
        RECT 18.490 53.280 18.780 53.325 ;
        RECT 20.325 53.280 20.615 53.325 ;
        RECT 23.905 53.280 24.195 53.325 ;
        RECT 18.490 53.140 24.195 53.280 ;
        RECT 18.490 53.095 18.780 53.140 ;
        RECT 20.325 53.095 20.615 53.140 ;
        RECT 23.905 53.095 24.195 53.140 ;
        RECT 24.985 53.120 25.275 53.435 ;
        RECT 28.130 53.080 28.450 53.340 ;
        RECT 29.525 53.280 29.815 53.325 ;
        RECT 31.810 53.280 32.130 53.340 ;
        RECT 29.525 53.140 32.130 53.280 ;
        RECT 29.525 53.095 29.815 53.140 ;
        RECT 31.810 53.080 32.130 53.140 ;
        RECT 32.745 53.095 33.035 53.325 ;
        RECT 7.890 52.800 9.040 52.940 ;
        RECT 7.890 52.740 8.210 52.800 ;
        RECT 8.365 52.755 8.655 52.800 ;
        RECT 8.900 52.260 9.040 52.800 ;
        RECT 17.105 52.800 17.780 52.940 ;
        RECT 17.105 52.755 17.395 52.800 ;
        RECT 18.025 52.755 18.315 52.985 ;
        RECT 19.390 52.940 19.710 53.000 ;
        RECT 32.820 52.940 32.960 53.095 ;
        RECT 35.490 53.080 35.810 53.340 ;
        RECT 37.345 53.280 37.635 53.325 ;
        RECT 43.325 53.280 43.615 53.325 ;
        RECT 43.770 53.280 44.090 53.340 ;
        RECT 37.345 53.140 44.090 53.280 ;
        RECT 37.345 53.095 37.635 53.140 ;
        RECT 43.325 53.095 43.615 53.140 ;
        RECT 37.420 52.940 37.560 53.095 ;
        RECT 43.770 53.080 44.090 53.140 ;
        RECT 46.545 53.280 46.835 53.325 ;
        RECT 46.990 53.280 47.310 53.340 ;
        RECT 46.545 53.140 47.310 53.280 ;
        RECT 47.565 53.280 47.780 53.435 ;
        RECT 52.970 53.420 53.290 53.480 ;
        RECT 54.365 53.435 54.655 53.480 ;
        RECT 56.205 53.620 56.495 53.665 ;
        RECT 58.950 53.620 59.270 53.680 ;
        RECT 62.645 53.620 62.935 53.665 ;
        RECT 56.205 53.480 62.935 53.620 ;
        RECT 56.205 53.435 56.495 53.480 ;
        RECT 58.950 53.420 59.270 53.480 ;
        RECT 62.645 53.435 62.935 53.480 ;
        RECT 64.470 53.420 64.790 53.680 ;
        RECT 66.310 53.620 66.630 53.680 ;
        RECT 77.350 53.665 77.670 53.680 ;
        RECT 65.480 53.480 66.630 53.620 ;
        RECT 49.810 53.280 50.100 53.325 ;
        RECT 59.425 53.280 59.715 53.325 ;
        RECT 63.550 53.280 63.870 53.340 ;
        RECT 65.480 53.325 65.620 53.480 ;
        RECT 66.310 53.420 66.630 53.480 ;
        RECT 73.785 53.620 74.075 53.665 ;
        RECT 77.025 53.620 77.675 53.665 ;
        RECT 73.785 53.480 77.675 53.620 ;
        RECT 73.785 53.435 74.375 53.480 ;
        RECT 77.025 53.435 77.675 53.480 ;
        RECT 65.405 53.280 65.695 53.325 ;
        RECT 68.150 53.280 68.470 53.340 ;
        RECT 70.925 53.280 71.215 53.325 ;
        RECT 47.565 53.140 50.100 53.280 ;
        RECT 46.545 53.095 46.835 53.140 ;
        RECT 46.990 53.080 47.310 53.140 ;
        RECT 49.810 53.095 50.100 53.140 ;
        RECT 50.760 53.140 65.695 53.280 ;
        RECT 19.390 52.800 24.680 52.940 ;
        RECT 32.820 52.800 37.560 52.940 ;
        RECT 9.235 52.600 9.525 52.645 ;
        RECT 11.125 52.600 11.415 52.645 ;
        RECT 14.245 52.600 14.535 52.645 ;
        RECT 18.100 52.600 18.240 52.755 ;
        RECT 19.390 52.740 19.710 52.800 ;
        RECT 9.235 52.460 14.535 52.600 ;
        RECT 9.235 52.415 9.525 52.460 ;
        RECT 11.125 52.415 11.415 52.460 ;
        RECT 14.245 52.415 14.535 52.460 ;
        RECT 16.720 52.460 18.240 52.600 ;
        RECT 18.895 52.600 19.185 52.645 ;
        RECT 20.785 52.600 21.075 52.645 ;
        RECT 23.905 52.600 24.195 52.645 ;
        RECT 18.895 52.460 24.195 52.600 ;
        RECT 16.720 52.260 16.860 52.460 ;
        RECT 8.900 52.120 16.860 52.260 ;
        RECT 17.640 52.260 17.780 52.460 ;
        RECT 18.895 52.415 19.185 52.460 ;
        RECT 20.785 52.415 21.075 52.460 ;
        RECT 23.905 52.415 24.195 52.460 ;
        RECT 20.310 52.260 20.630 52.320 ;
        RECT 17.640 52.120 20.630 52.260 ;
        RECT 24.540 52.260 24.680 52.800 ;
        RECT 44.690 52.740 45.010 53.000 ;
        RECT 45.170 52.600 45.460 52.645 ;
        RECT 47.030 52.600 47.320 52.645 ;
        RECT 49.810 52.600 50.100 52.645 ;
        RECT 45.170 52.460 50.100 52.600 ;
        RECT 45.170 52.415 45.460 52.460 ;
        RECT 47.030 52.415 47.320 52.460 ;
        RECT 49.810 52.415 50.100 52.460 ;
        RECT 50.760 52.260 50.900 53.140 ;
        RECT 59.425 53.095 59.715 53.140 ;
        RECT 63.550 53.080 63.870 53.140 ;
        RECT 65.405 53.095 65.695 53.140 ;
        RECT 66.400 53.140 71.215 53.280 ;
        RECT 56.650 52.940 56.970 53.000 ;
        RECT 60.805 52.940 61.095 52.985 ;
        RECT 56.650 52.800 61.095 52.940 ;
        RECT 56.650 52.740 56.970 52.800 ;
        RECT 60.805 52.755 61.095 52.800 ;
        RECT 65.850 52.940 66.170 53.000 ;
        RECT 66.400 52.985 66.540 53.140 ;
        RECT 68.150 53.080 68.470 53.140 ;
        RECT 70.925 53.095 71.215 53.140 ;
        RECT 74.085 53.120 74.375 53.435 ;
        RECT 77.350 53.420 77.670 53.435 ;
        RECT 79.650 53.420 79.970 53.680 ;
        RECT 87.005 53.620 87.655 53.665 ;
        RECT 90.605 53.620 90.895 53.665 ;
        RECT 93.005 53.620 93.295 53.665 ;
        RECT 87.005 53.480 93.295 53.620 ;
        RECT 87.005 53.435 87.655 53.480 ;
        RECT 90.305 53.435 90.895 53.480 ;
        RECT 93.005 53.435 93.295 53.480 ;
        RECT 99.910 53.620 100.200 53.665 ;
        RECT 101.770 53.620 102.060 53.665 ;
        RECT 99.910 53.480 102.060 53.620 ;
        RECT 99.910 53.435 100.200 53.480 ;
        RECT 101.770 53.435 102.060 53.480 ;
        RECT 102.690 53.620 102.980 53.665 ;
        RECT 105.950 53.620 106.240 53.665 ;
        RECT 110.010 53.620 110.330 53.680 ;
        RECT 102.690 53.480 110.330 53.620 ;
        RECT 102.690 53.435 102.980 53.480 ;
        RECT 105.950 53.435 106.240 53.480 ;
        RECT 75.165 53.280 75.455 53.325 ;
        RECT 78.745 53.280 79.035 53.325 ;
        RECT 80.580 53.280 80.870 53.325 ;
        RECT 75.165 53.140 80.870 53.280 ;
        RECT 75.165 53.095 75.455 53.140 ;
        RECT 78.745 53.095 79.035 53.140 ;
        RECT 80.580 53.095 80.870 53.140 ;
        RECT 83.810 53.280 84.100 53.325 ;
        RECT 85.645 53.280 85.935 53.325 ;
        RECT 89.225 53.280 89.515 53.325 ;
        RECT 83.810 53.140 89.515 53.280 ;
        RECT 83.810 53.095 84.100 53.140 ;
        RECT 85.645 53.095 85.935 53.140 ;
        RECT 89.225 53.095 89.515 53.140 ;
        RECT 90.305 53.120 90.595 53.435 ;
        RECT 92.530 53.280 92.850 53.340 ;
        RECT 93.465 53.280 93.755 53.325 ;
        RECT 95.305 53.280 95.595 53.325 ;
        RECT 92.530 53.140 95.595 53.280 ;
        RECT 92.530 53.080 92.850 53.140 ;
        RECT 93.465 53.095 93.755 53.140 ;
        RECT 95.305 53.095 95.595 53.140 ;
        RECT 98.050 53.280 98.370 53.340 ;
        RECT 100.825 53.280 101.115 53.325 ;
        RECT 98.050 53.140 101.115 53.280 ;
        RECT 101.845 53.280 102.060 53.435 ;
        RECT 110.010 53.420 110.330 53.480 ;
        RECT 104.090 53.280 104.380 53.325 ;
        RECT 101.845 53.140 104.380 53.280 ;
        RECT 98.050 53.080 98.370 53.140 ;
        RECT 100.825 53.095 101.115 53.140 ;
        RECT 104.090 53.095 104.380 53.140 ;
        RECT 66.325 52.940 66.615 52.985 ;
        RECT 65.850 52.800 66.615 52.940 ;
        RECT 60.880 52.600 61.020 52.755 ;
        RECT 65.850 52.740 66.170 52.800 ;
        RECT 66.325 52.755 66.615 52.800 ;
        RECT 72.305 52.940 72.595 52.985 ;
        RECT 73.670 52.940 73.990 53.000 ;
        RECT 81.045 52.940 81.335 52.985 ;
        RECT 72.305 52.800 73.990 52.940 ;
        RECT 72.305 52.755 72.595 52.800 ;
        RECT 73.670 52.740 73.990 52.800 ;
        RECT 80.660 52.800 81.335 52.940 ;
        RECT 75.165 52.600 75.455 52.645 ;
        RECT 78.285 52.600 78.575 52.645 ;
        RECT 80.175 52.600 80.465 52.645 ;
        RECT 60.880 52.460 72.520 52.600 ;
        RECT 72.380 52.320 72.520 52.460 ;
        RECT 75.165 52.460 80.465 52.600 ;
        RECT 75.165 52.415 75.455 52.460 ;
        RECT 78.285 52.415 78.575 52.460 ;
        RECT 80.175 52.415 80.465 52.460 ;
        RECT 24.540 52.120 50.900 52.260 ;
        RECT 58.490 52.260 58.810 52.320 ;
        RECT 61.710 52.260 62.030 52.320 ;
        RECT 58.490 52.120 62.030 52.260 ;
        RECT 20.310 52.060 20.630 52.120 ;
        RECT 58.490 52.060 58.810 52.120 ;
        RECT 61.710 52.060 62.030 52.120 ;
        RECT 72.290 52.060 72.610 52.320 ;
        RECT 72.750 52.260 73.070 52.320 ;
        RECT 80.660 52.260 80.800 52.800 ;
        RECT 81.045 52.755 81.335 52.800 ;
        RECT 83.330 52.740 83.650 53.000 ;
        RECT 84.725 52.940 85.015 52.985 ;
        RECT 86.550 52.940 86.870 53.000 ;
        RECT 84.725 52.800 86.870 52.940 ;
        RECT 84.725 52.755 85.015 52.800 ;
        RECT 86.550 52.740 86.870 52.800 ;
        RECT 98.970 52.740 99.290 53.000 ;
        RECT 84.215 52.600 84.505 52.645 ;
        RECT 86.105 52.600 86.395 52.645 ;
        RECT 89.225 52.600 89.515 52.645 ;
        RECT 84.215 52.460 89.515 52.600 ;
        RECT 84.215 52.415 84.505 52.460 ;
        RECT 86.105 52.415 86.395 52.460 ;
        RECT 89.225 52.415 89.515 52.460 ;
        RECT 99.450 52.600 99.740 52.645 ;
        RECT 101.310 52.600 101.600 52.645 ;
        RECT 104.090 52.600 104.380 52.645 ;
        RECT 99.450 52.460 104.380 52.600 ;
        RECT 99.450 52.415 99.740 52.460 ;
        RECT 101.310 52.415 101.600 52.460 ;
        RECT 104.090 52.415 104.380 52.460 ;
        RECT 72.750 52.120 80.800 52.260 ;
        RECT 72.750 52.060 73.070 52.120 ;
        RECT 94.830 52.060 95.150 52.320 ;
        RECT 102.650 52.260 102.970 52.320 ;
        RECT 107.955 52.260 108.245 52.305 ;
        RECT 102.650 52.120 108.245 52.260 ;
        RECT 102.650 52.060 102.970 52.120 ;
        RECT 107.955 52.075 108.245 52.120 ;
        RECT 5.520 51.440 113.620 51.920 ;
        RECT 13.870 51.040 14.190 51.300 ;
        RECT 52.510 51.240 52.830 51.300 ;
        RECT 31.440 51.100 39.860 51.240 ;
        RECT 9.285 50.900 9.575 50.945 ;
        RECT 12.950 50.900 13.270 50.960 ;
        RECT 9.285 50.760 13.270 50.900 ;
        RECT 9.285 50.715 9.575 50.760 ;
        RECT 12.950 50.700 13.270 50.760 ;
        RECT 13.425 50.900 13.715 50.945 ;
        RECT 21.690 50.900 22.010 50.960 ;
        RECT 13.425 50.760 22.010 50.900 ;
        RECT 13.425 50.715 13.715 50.760 ;
        RECT 21.690 50.700 22.010 50.760 ;
        RECT 23.070 50.900 23.390 50.960 ;
        RECT 30.890 50.900 31.210 50.960 ;
        RECT 23.070 50.760 31.210 50.900 ;
        RECT 23.070 50.700 23.390 50.760 ;
        RECT 30.890 50.700 31.210 50.760 ;
        RECT 10.665 50.375 10.955 50.605 ;
        RECT 16.645 50.560 16.935 50.605 ;
        RECT 22.150 50.560 22.470 50.620 ;
        RECT 31.440 50.605 31.580 51.100 ;
        RECT 36.885 50.715 37.175 50.945 ;
        RECT 31.365 50.560 31.655 50.605 ;
        RECT 13.730 50.420 31.655 50.560 ;
        RECT 10.740 50.220 10.880 50.375 ;
        RECT 13.730 50.220 13.870 50.420 ;
        RECT 16.645 50.375 16.935 50.420 ;
        RECT 22.150 50.360 22.470 50.420 ;
        RECT 31.365 50.375 31.655 50.420 ;
        RECT 10.740 50.080 13.870 50.220 ;
        RECT 16.185 50.220 16.475 50.265 ;
        RECT 21.230 50.220 21.550 50.280 ;
        RECT 16.185 50.080 21.550 50.220 ;
        RECT 16.185 50.035 16.475 50.080 ;
        RECT 21.230 50.020 21.550 50.080 ;
        RECT 28.590 50.220 28.910 50.280 ;
        RECT 30.445 50.220 30.735 50.265 ;
        RECT 28.590 50.080 30.735 50.220 ;
        RECT 28.590 50.020 28.910 50.080 ;
        RECT 30.445 50.035 30.735 50.080 ;
        RECT 8.350 49.680 8.670 49.940 ;
        RECT 11.110 49.880 11.430 49.940 ;
        RECT 15.725 49.880 16.015 49.925 ;
        RECT 17.550 49.880 17.870 49.940 ;
        RECT 23.070 49.880 23.390 49.940 ;
        RECT 11.110 49.740 17.870 49.880 ;
        RECT 11.110 49.680 11.430 49.740 ;
        RECT 15.725 49.695 16.015 49.740 ;
        RECT 17.550 49.680 17.870 49.740 ;
        RECT 20.400 49.740 23.390 49.880 ;
        RECT 11.585 49.540 11.875 49.585 ;
        RECT 20.400 49.540 20.540 49.740 ;
        RECT 23.070 49.680 23.390 49.740 ;
        RECT 28.130 49.680 28.450 49.940 ;
        RECT 30.520 49.880 30.660 50.035 ;
        RECT 30.890 50.020 31.210 50.280 ;
        RECT 36.425 50.220 36.715 50.265 ;
        RECT 36.960 50.220 37.100 50.715 ;
        RECT 39.720 50.605 39.860 51.100 ;
        RECT 43.400 51.100 52.830 51.240 ;
        RECT 39.645 50.375 39.935 50.605 ;
        RECT 36.425 50.080 37.100 50.220 ;
        RECT 42.865 50.220 43.155 50.265 ;
        RECT 43.400 50.220 43.540 51.100 ;
        RECT 52.510 51.040 52.830 51.100 ;
        RECT 58.950 51.040 59.270 51.300 ;
        RECT 77.350 51.040 77.670 51.300 ;
        RECT 86.565 51.240 86.855 51.285 ;
        RECT 87.470 51.240 87.790 51.300 ;
        RECT 86.565 51.100 87.790 51.240 ;
        RECT 86.565 51.055 86.855 51.100 ;
        RECT 87.470 51.040 87.790 51.100 ;
        RECT 97.130 51.240 97.450 51.300 ;
        RECT 101.285 51.240 101.575 51.285 ;
        RECT 97.130 51.100 101.575 51.240 ;
        RECT 97.130 51.040 97.450 51.100 ;
        RECT 101.285 51.055 101.575 51.100 ;
        RECT 43.785 50.715 44.075 50.945 ;
        RECT 45.170 50.900 45.460 50.945 ;
        RECT 47.030 50.900 47.320 50.945 ;
        RECT 49.810 50.900 50.100 50.945 ;
        RECT 45.170 50.760 50.100 50.900 ;
        RECT 45.170 50.715 45.460 50.760 ;
        RECT 47.030 50.715 47.320 50.760 ;
        RECT 49.810 50.715 50.100 50.760 ;
        RECT 43.860 50.560 44.000 50.715 ;
        RECT 62.630 50.700 62.950 50.960 ;
        RECT 87.010 50.900 87.330 50.960 ;
        RECT 92.530 50.900 92.850 50.960 ;
        RECT 77.900 50.760 92.850 50.900 ;
        RECT 46.545 50.560 46.835 50.605 ;
        RECT 43.860 50.420 46.835 50.560 ;
        RECT 46.545 50.375 46.835 50.420 ;
        RECT 58.030 50.360 58.350 50.620 ;
        RECT 58.490 50.560 58.810 50.620 ;
        RECT 60.330 50.560 60.650 50.620 ;
        RECT 58.490 50.420 60.650 50.560 ;
        RECT 58.490 50.360 58.810 50.420 ;
        RECT 60.330 50.360 60.650 50.420 ;
        RECT 42.865 50.080 43.540 50.220 ;
        RECT 36.425 50.035 36.715 50.080 ;
        RECT 42.865 50.035 43.155 50.080 ;
        RECT 44.690 50.020 45.010 50.280 ;
        RECT 49.810 50.220 50.100 50.265 ;
        RECT 47.565 50.080 50.100 50.220 ;
        RECT 39.185 49.880 39.475 49.925 ;
        RECT 41.930 49.880 42.250 49.940 ;
        RECT 47.565 49.925 47.780 50.080 ;
        RECT 49.810 50.035 50.100 50.080 ;
        RECT 58.950 50.220 59.270 50.280 ;
        RECT 59.425 50.220 59.715 50.265 ;
        RECT 58.950 50.080 59.715 50.220 ;
        RECT 58.950 50.020 59.270 50.080 ;
        RECT 59.425 50.035 59.715 50.080 ;
        RECT 59.870 50.020 60.190 50.280 ;
        RECT 63.550 50.020 63.870 50.280 ;
        RECT 68.150 50.220 68.470 50.280 ;
        RECT 77.900 50.265 78.040 50.760 ;
        RECT 87.010 50.700 87.330 50.760 ;
        RECT 92.530 50.700 92.850 50.760 ;
        RECT 90.690 50.560 91.010 50.620 ;
        RECT 84.340 50.420 91.010 50.560 ;
        RECT 84.340 50.265 84.480 50.420 ;
        RECT 90.690 50.360 91.010 50.420 ;
        RECT 102.190 50.560 102.510 50.620 ;
        RECT 104.045 50.560 104.335 50.605 ;
        RECT 102.190 50.420 104.335 50.560 ;
        RECT 102.190 50.360 102.510 50.420 ;
        RECT 104.045 50.375 104.335 50.420 ;
        RECT 77.825 50.220 78.115 50.265 ;
        RECT 68.150 50.080 78.115 50.220 ;
        RECT 68.150 50.020 68.470 50.080 ;
        RECT 77.825 50.035 78.115 50.080 ;
        RECT 83.345 50.035 83.635 50.265 ;
        RECT 84.265 50.035 84.555 50.265 ;
        RECT 84.725 50.035 85.015 50.265 ;
        RECT 85.185 50.220 85.475 50.265 ;
        RECT 86.550 50.220 86.870 50.280 ;
        RECT 85.185 50.080 86.870 50.220 ;
        RECT 85.185 50.035 85.475 50.080 ;
        RECT 30.520 49.740 42.250 49.880 ;
        RECT 39.185 49.695 39.475 49.740 ;
        RECT 41.930 49.680 42.250 49.740 ;
        RECT 45.630 49.880 45.920 49.925 ;
        RECT 47.490 49.880 47.780 49.925 ;
        RECT 45.630 49.740 47.780 49.880 ;
        RECT 45.630 49.695 45.920 49.740 ;
        RECT 47.490 49.695 47.780 49.740 ;
        RECT 48.410 49.880 48.700 49.925 ;
        RECT 49.290 49.880 49.610 49.940 ;
        RECT 51.670 49.880 51.960 49.925 ;
        RECT 48.410 49.740 51.960 49.880 ;
        RECT 48.410 49.695 48.700 49.740 ;
        RECT 49.290 49.680 49.610 49.740 ;
        RECT 51.670 49.695 51.960 49.740 ;
        RECT 68.610 49.880 68.930 49.940 ;
        RECT 83.420 49.880 83.560 50.035 ;
        RECT 68.610 49.740 83.560 49.880 ;
        RECT 83.790 49.880 84.110 49.940 ;
        RECT 84.800 49.880 84.940 50.035 ;
        RECT 86.550 50.020 86.870 50.080 ;
        RECT 103.110 50.020 103.430 50.280 ;
        RECT 83.790 49.740 84.940 49.880 ;
        RECT 97.590 49.880 97.910 49.940 ;
        RECT 102.650 49.880 102.970 49.940 ;
        RECT 103.585 49.880 103.875 49.925 ;
        RECT 97.590 49.740 103.875 49.880 ;
        RECT 68.610 49.680 68.930 49.740 ;
        RECT 83.790 49.680 84.110 49.740 ;
        RECT 97.590 49.680 97.910 49.740 ;
        RECT 102.650 49.680 102.970 49.740 ;
        RECT 103.585 49.695 103.875 49.740 ;
        RECT 11.585 49.400 20.540 49.540 ;
        RECT 11.585 49.355 11.875 49.400 ;
        RECT 20.770 49.340 21.090 49.600 ;
        RECT 21.230 49.540 21.550 49.600 ;
        RECT 28.605 49.540 28.895 49.585 ;
        RECT 21.230 49.400 28.895 49.540 ;
        RECT 21.230 49.340 21.550 49.400 ;
        RECT 28.605 49.355 28.895 49.400 ;
        RECT 34.570 49.540 34.890 49.600 ;
        RECT 53.430 49.585 53.750 49.600 ;
        RECT 35.505 49.540 35.795 49.585 ;
        RECT 34.570 49.400 35.795 49.540 ;
        RECT 34.570 49.340 34.890 49.400 ;
        RECT 35.505 49.355 35.795 49.400 ;
        RECT 38.725 49.540 39.015 49.585 ;
        RECT 53.430 49.540 53.965 49.585 ;
        RECT 38.725 49.400 53.965 49.540 ;
        RECT 38.725 49.355 39.015 49.400 ;
        RECT 53.430 49.355 53.965 49.400 ;
        RECT 53.430 49.340 53.750 49.355 ;
        RECT 5.520 48.720 113.620 49.200 ;
        RECT 8.365 48.520 8.655 48.565 ;
        RECT 11.110 48.520 11.430 48.580 ;
        RECT 8.365 48.380 11.430 48.520 ;
        RECT 8.365 48.335 8.655 48.380 ;
        RECT 11.110 48.320 11.430 48.380 ;
        RECT 59.885 48.520 60.175 48.565 ;
        RECT 64.930 48.520 65.250 48.580 ;
        RECT 68.610 48.520 68.930 48.580 ;
        RECT 59.885 48.380 68.930 48.520 ;
        RECT 59.885 48.335 60.175 48.380 ;
        RECT 64.930 48.320 65.250 48.380 ;
        RECT 68.610 48.320 68.930 48.380 ;
        RECT 9.845 48.180 10.135 48.225 ;
        RECT 13.085 48.180 13.735 48.225 ;
        RECT 17.550 48.180 17.870 48.240 ;
        RECT 21.230 48.180 21.550 48.240 ;
        RECT 35.950 48.180 36.270 48.240 ;
        RECT 9.845 48.040 17.870 48.180 ;
        RECT 9.845 47.995 10.435 48.040 ;
        RECT 13.085 47.995 13.735 48.040 ;
        RECT 10.145 47.680 10.435 47.995 ;
        RECT 17.550 47.980 17.870 48.040 ;
        RECT 18.100 48.040 21.550 48.180 ;
        RECT 18.100 47.885 18.240 48.040 ;
        RECT 21.230 47.980 21.550 48.040 ;
        RECT 33.280 48.040 36.270 48.180 ;
        RECT 11.225 47.840 11.515 47.885 ;
        RECT 14.805 47.840 15.095 47.885 ;
        RECT 16.640 47.840 16.930 47.885 ;
        RECT 11.225 47.700 16.930 47.840 ;
        RECT 11.225 47.655 11.515 47.700 ;
        RECT 14.805 47.655 15.095 47.700 ;
        RECT 16.640 47.655 16.930 47.700 ;
        RECT 18.025 47.655 18.315 47.885 ;
        RECT 19.405 47.840 19.695 47.885 ;
        RECT 32.730 47.840 33.050 47.900 ;
        RECT 33.280 47.885 33.420 48.040 ;
        RECT 35.950 47.980 36.270 48.040 ;
        RECT 36.865 48.180 37.515 48.225 ;
        RECT 40.465 48.180 40.755 48.225 ;
        RECT 42.865 48.180 43.155 48.225 ;
        RECT 36.865 48.040 43.155 48.180 ;
        RECT 36.865 47.995 37.515 48.040 ;
        RECT 40.165 47.995 40.755 48.040 ;
        RECT 42.865 47.995 43.155 48.040 ;
        RECT 48.845 48.180 49.135 48.225 ;
        RECT 49.290 48.180 49.610 48.240 ;
        RECT 48.845 48.040 49.610 48.180 ;
        RECT 48.845 47.995 49.135 48.040 ;
        RECT 33.205 47.840 33.495 47.885 ;
        RECT 19.405 47.700 19.805 47.840 ;
        RECT 32.730 47.700 33.495 47.840 ;
        RECT 19.405 47.655 19.695 47.700 ;
        RECT 15.710 47.300 16.030 47.560 ;
        RECT 17.105 47.500 17.395 47.545 ;
        RECT 19.480 47.500 19.620 47.655 ;
        RECT 32.730 47.640 33.050 47.700 ;
        RECT 33.205 47.655 33.495 47.700 ;
        RECT 33.670 47.840 33.960 47.885 ;
        RECT 35.505 47.840 35.795 47.885 ;
        RECT 39.085 47.840 39.375 47.885 ;
        RECT 33.670 47.700 39.375 47.840 ;
        RECT 33.670 47.655 33.960 47.700 ;
        RECT 35.505 47.655 35.795 47.700 ;
        RECT 39.085 47.655 39.375 47.700 ;
        RECT 40.165 47.680 40.455 47.995 ;
        RECT 49.290 47.980 49.610 48.040 ;
        RECT 54.350 48.180 54.670 48.240 ;
        RECT 62.630 48.180 62.950 48.240 ;
        RECT 64.470 48.180 64.790 48.240 ;
        RECT 54.350 48.040 64.790 48.180 ;
        RECT 54.350 47.980 54.670 48.040 ;
        RECT 62.630 47.980 62.950 48.040 ;
        RECT 64.470 47.980 64.790 48.040 ;
        RECT 78.730 47.980 79.050 48.240 ;
        RECT 87.485 48.180 87.775 48.225 ;
        RECT 87.930 48.180 88.250 48.240 ;
        RECT 87.485 48.040 88.250 48.180 ;
        RECT 87.485 47.995 87.775 48.040 ;
        RECT 87.930 47.980 88.250 48.040 ;
        RECT 89.765 48.180 90.415 48.225 ;
        RECT 93.365 48.180 93.655 48.225 ;
        RECT 94.830 48.180 95.150 48.240 ;
        RECT 89.765 48.040 95.150 48.180 ;
        RECT 89.765 47.995 90.415 48.040 ;
        RECT 93.065 47.995 93.655 48.040 ;
        RECT 43.310 47.640 43.630 47.900 ;
        RECT 43.770 47.840 44.090 47.900 ;
        RECT 48.385 47.840 48.675 47.885 ;
        RECT 43.770 47.700 48.675 47.840 ;
        RECT 43.770 47.640 44.090 47.700 ;
        RECT 48.385 47.655 48.675 47.700 ;
        RECT 58.030 47.840 58.350 47.900 ;
        RECT 60.805 47.840 61.095 47.885 ;
        RECT 61.265 47.840 61.555 47.885 ;
        RECT 58.030 47.700 61.555 47.840 ;
        RECT 58.030 47.640 58.350 47.700 ;
        RECT 60.805 47.655 61.095 47.700 ;
        RECT 61.265 47.655 61.555 47.700 ;
        RECT 69.070 47.840 69.390 47.900 ;
        RECT 72.750 47.840 73.070 47.900 ;
        RECT 69.070 47.700 73.070 47.840 ;
        RECT 69.070 47.640 69.390 47.700 ;
        RECT 72.750 47.640 73.070 47.700 ;
        RECT 75.510 47.640 75.830 47.900 ;
        RECT 75.970 47.840 76.290 47.900 ;
        RECT 76.445 47.840 76.735 47.885 ;
        RECT 75.970 47.700 76.735 47.840 ;
        RECT 75.970 47.640 76.290 47.700 ;
        RECT 76.445 47.655 76.735 47.700 ;
        RECT 76.905 47.655 77.195 47.885 ;
        RECT 20.770 47.500 21.090 47.560 ;
        RECT 23.530 47.500 23.850 47.560 ;
        RECT 17.105 47.360 23.850 47.500 ;
        RECT 17.105 47.315 17.395 47.360 ;
        RECT 20.770 47.300 21.090 47.360 ;
        RECT 23.530 47.300 23.850 47.360 ;
        RECT 34.570 47.300 34.890 47.560 ;
        RECT 41.930 47.300 42.250 47.560 ;
        RECT 53.430 47.500 53.750 47.560 ;
        RECT 63.090 47.500 63.410 47.560 ;
        RECT 76.980 47.500 77.120 47.655 ;
        RECT 77.350 47.640 77.670 47.900 ;
        RECT 86.570 47.840 86.860 47.885 ;
        RECT 88.405 47.840 88.695 47.885 ;
        RECT 91.985 47.840 92.275 47.885 ;
        RECT 86.570 47.700 92.275 47.840 ;
        RECT 86.570 47.655 86.860 47.700 ;
        RECT 88.405 47.655 88.695 47.700 ;
        RECT 91.985 47.655 92.275 47.700 ;
        RECT 93.065 47.680 93.355 47.995 ;
        RECT 94.830 47.980 95.150 48.040 ;
        RECT 96.225 47.840 96.515 47.885 ;
        RECT 98.970 47.840 99.290 47.900 ;
        RECT 96.225 47.700 99.290 47.840 ;
        RECT 96.225 47.655 96.515 47.700 ;
        RECT 81.030 47.500 81.350 47.560 ;
        RECT 53.430 47.360 81.350 47.500 ;
        RECT 53.430 47.300 53.750 47.360 ;
        RECT 63.090 47.300 63.410 47.360 ;
        RECT 81.030 47.300 81.350 47.360 ;
        RECT 83.330 47.500 83.650 47.560 ;
        RECT 86.090 47.500 86.410 47.560 ;
        RECT 83.330 47.360 86.410 47.500 ;
        RECT 83.330 47.300 83.650 47.360 ;
        RECT 86.090 47.300 86.410 47.360 ;
        RECT 94.830 47.300 95.150 47.560 ;
        RECT 11.225 47.160 11.515 47.205 ;
        RECT 14.345 47.160 14.635 47.205 ;
        RECT 16.235 47.160 16.525 47.205 ;
        RECT 11.225 47.020 16.525 47.160 ;
        RECT 11.225 46.975 11.515 47.020 ;
        RECT 14.345 46.975 14.635 47.020 ;
        RECT 16.235 46.975 16.525 47.020 ;
        RECT 34.075 47.160 34.365 47.205 ;
        RECT 35.965 47.160 36.255 47.205 ;
        RECT 39.085 47.160 39.375 47.205 ;
        RECT 34.075 47.020 39.375 47.160 ;
        RECT 34.075 46.975 34.365 47.020 ;
        RECT 35.965 46.975 36.255 47.020 ;
        RECT 39.085 46.975 39.375 47.020 ;
        RECT 42.390 47.160 42.710 47.220 ;
        RECT 62.185 47.160 62.475 47.205 ;
        RECT 82.870 47.160 83.190 47.220 ;
        RECT 42.390 47.020 83.190 47.160 ;
        RECT 42.390 46.960 42.710 47.020 ;
        RECT 62.185 46.975 62.475 47.020 ;
        RECT 82.870 46.960 83.190 47.020 ;
        RECT 86.975 47.160 87.265 47.205 ;
        RECT 88.865 47.160 89.155 47.205 ;
        RECT 91.985 47.160 92.275 47.205 ;
        RECT 86.975 47.020 92.275 47.160 ;
        RECT 86.975 46.975 87.265 47.020 ;
        RECT 88.865 46.975 89.155 47.020 ;
        RECT 91.985 46.975 92.275 47.020 ;
        RECT 18.930 46.620 19.250 46.880 ;
        RECT 33.650 46.820 33.970 46.880 ;
        RECT 56.650 46.820 56.970 46.880 ;
        RECT 33.650 46.680 56.970 46.820 ;
        RECT 33.650 46.620 33.970 46.680 ;
        RECT 56.650 46.620 56.970 46.680 ;
        RECT 86.090 46.820 86.410 46.880 ;
        RECT 87.470 46.820 87.790 46.880 ;
        RECT 96.300 46.820 96.440 47.655 ;
        RECT 98.970 47.640 99.290 47.700 ;
        RECT 86.090 46.680 96.440 46.820 ;
        RECT 86.090 46.620 86.410 46.680 ;
        RECT 87.470 46.620 87.790 46.680 ;
        RECT 5.520 46.000 113.620 46.480 ;
        RECT 17.550 45.600 17.870 45.860 ;
        RECT 18.930 45.800 19.250 45.860 ;
        RECT 22.990 45.800 23.280 45.845 ;
        RECT 18.930 45.660 23.280 45.800 ;
        RECT 18.930 45.600 19.250 45.660 ;
        RECT 22.990 45.615 23.280 45.660 ;
        RECT 30.445 45.800 30.735 45.845 ;
        RECT 30.890 45.800 31.210 45.860 ;
        RECT 30.445 45.660 31.210 45.800 ;
        RECT 30.445 45.615 30.735 45.660 ;
        RECT 30.890 45.600 31.210 45.660 ;
        RECT 51.130 45.600 51.450 45.860 ;
        RECT 61.250 45.800 61.570 45.860 ;
        RECT 51.680 45.660 61.570 45.800 ;
        RECT 15.710 45.460 16.030 45.520 ;
        RECT 20.325 45.460 20.615 45.505 ;
        RECT 15.710 45.320 20.615 45.460 ;
        RECT 15.710 45.260 16.030 45.320 ;
        RECT 20.325 45.275 20.615 45.320 ;
        RECT 22.575 45.460 22.865 45.505 ;
        RECT 24.465 45.460 24.755 45.505 ;
        RECT 27.585 45.460 27.875 45.505 ;
        RECT 22.575 45.320 27.875 45.460 ;
        RECT 22.575 45.275 22.865 45.320 ;
        RECT 24.465 45.275 24.755 45.320 ;
        RECT 27.585 45.275 27.875 45.320 ;
        RECT 33.190 45.460 33.510 45.520 ;
        RECT 51.680 45.460 51.820 45.660 ;
        RECT 61.250 45.600 61.570 45.660 ;
        RECT 63.090 45.600 63.410 45.860 ;
        RECT 81.950 45.600 82.270 45.860 ;
        RECT 83.330 45.800 83.650 45.860 ;
        RECT 85.170 45.800 85.490 45.860 ;
        RECT 83.330 45.660 85.490 45.800 ;
        RECT 83.330 45.600 83.650 45.660 ;
        RECT 85.170 45.600 85.490 45.660 ;
        RECT 85.630 45.600 85.950 45.860 ;
        RECT 88.850 45.800 89.170 45.860 ;
        RECT 89.325 45.800 89.615 45.845 ;
        RECT 88.850 45.660 89.615 45.800 ;
        RECT 88.850 45.600 89.170 45.660 ;
        RECT 89.325 45.615 89.615 45.660 ;
        RECT 98.970 45.800 99.290 45.860 ;
        RECT 102.650 45.800 102.970 45.860 ;
        RECT 98.970 45.660 102.970 45.800 ;
        RECT 98.970 45.600 99.290 45.660 ;
        RECT 102.650 45.600 102.970 45.660 ;
        RECT 33.190 45.320 51.820 45.460 ;
        RECT 56.650 45.460 56.970 45.520 ;
        RECT 57.125 45.460 57.415 45.505 ;
        RECT 60.805 45.460 61.095 45.505 ;
        RECT 77.350 45.460 77.670 45.520 ;
        RECT 56.650 45.320 57.415 45.460 ;
        RECT 33.190 45.260 33.510 45.320 ;
        RECT 56.650 45.260 56.970 45.320 ;
        RECT 57.125 45.275 57.415 45.320 ;
        RECT 57.660 45.320 77.670 45.460 ;
        RECT 17.090 45.120 17.410 45.180 ;
        RECT 19.405 45.120 19.695 45.165 ;
        RECT 17.090 44.980 19.695 45.120 ;
        RECT 17.090 44.920 17.410 44.980 ;
        RECT 19.405 44.935 19.695 44.980 ;
        RECT 21.705 45.120 21.995 45.165 ;
        RECT 23.530 45.120 23.850 45.180 ;
        RECT 54.350 45.120 54.670 45.180 ;
        RECT 21.705 44.980 23.850 45.120 ;
        RECT 21.705 44.935 21.995 44.980 ;
        RECT 23.530 44.920 23.850 44.980 ;
        RECT 47.080 44.980 54.670 45.120 ;
        RECT 18.025 44.780 18.315 44.825 ;
        RECT 19.865 44.780 20.155 44.825 ;
        RECT 18.025 44.640 20.155 44.780 ;
        RECT 18.025 44.595 18.315 44.640 ;
        RECT 19.865 44.595 20.155 44.640 ;
        RECT 19.940 44.100 20.080 44.595 ;
        RECT 21.230 44.580 21.550 44.840 ;
        RECT 22.170 44.780 22.460 44.825 ;
        RECT 24.005 44.780 24.295 44.825 ;
        RECT 27.585 44.780 27.875 44.825 ;
        RECT 22.170 44.640 27.875 44.780 ;
        RECT 22.170 44.595 22.460 44.640 ;
        RECT 24.005 44.595 24.295 44.640 ;
        RECT 27.585 44.595 27.875 44.640 ;
        RECT 28.665 44.485 28.955 44.800 ;
        RECT 31.810 44.580 32.130 44.840 ;
        RECT 35.950 44.780 36.270 44.840 ;
        RECT 38.250 44.780 38.570 44.840 ;
        RECT 44.690 44.780 45.010 44.840 ;
        RECT 47.080 44.825 47.220 44.980 ;
        RECT 54.350 44.920 54.670 44.980 ;
        RECT 35.950 44.640 45.010 44.780 ;
        RECT 35.950 44.580 36.270 44.640 ;
        RECT 38.250 44.580 38.570 44.640 ;
        RECT 44.690 44.580 45.010 44.640 ;
        RECT 47.005 44.595 47.295 44.825 ;
        RECT 47.925 44.595 48.215 44.825 ;
        RECT 25.365 44.440 26.015 44.485 ;
        RECT 28.665 44.440 29.255 44.485 ;
        RECT 31.365 44.440 31.655 44.485 ;
        RECT 25.365 44.300 31.655 44.440 ;
        RECT 25.365 44.255 26.015 44.300 ;
        RECT 28.965 44.255 29.255 44.300 ;
        RECT 31.365 44.255 31.655 44.300 ;
        RECT 31.900 44.440 32.040 44.580 ;
        RECT 43.310 44.440 43.630 44.500 ;
        RECT 45.625 44.440 45.915 44.485 ;
        RECT 47.450 44.440 47.770 44.500 ;
        RECT 31.900 44.300 47.770 44.440 ;
        RECT 48.000 44.440 48.140 44.595 ;
        RECT 48.830 44.580 49.150 44.840 ;
        RECT 49.290 44.580 49.610 44.840 ;
        RECT 49.765 44.780 50.055 44.825 ;
        RECT 53.890 44.780 54.210 44.840 ;
        RECT 57.660 44.780 57.800 45.320 ;
        RECT 60.805 45.275 61.095 45.320 ;
        RECT 77.350 45.260 77.670 45.320 ;
        RECT 85.260 45.320 89.080 45.460 ;
        RECT 62.630 45.120 62.950 45.180 ;
        RECT 58.120 44.980 62.950 45.120 ;
        RECT 58.120 44.825 58.260 44.980 ;
        RECT 49.765 44.640 57.800 44.780 ;
        RECT 49.765 44.595 50.055 44.640 ;
        RECT 53.890 44.580 54.210 44.640 ;
        RECT 58.045 44.595 58.335 44.825 ;
        RECT 58.505 44.780 58.795 44.825 ;
        RECT 59.410 44.780 59.730 44.840 ;
        RECT 62.260 44.825 62.400 44.980 ;
        RECT 62.630 44.920 62.950 44.980 ;
        RECT 75.510 45.120 75.830 45.180 ;
        RECT 81.490 45.120 81.810 45.180 ;
        RECT 85.260 45.120 85.400 45.320 ;
        RECT 75.510 44.980 85.400 45.120 ;
        RECT 75.510 44.920 75.830 44.980 ;
        RECT 81.490 44.920 81.810 44.980 ;
        RECT 61.725 44.780 62.015 44.825 ;
        RECT 58.505 44.640 59.180 44.780 ;
        RECT 58.505 44.595 58.795 44.640 ;
        RECT 48.370 44.440 48.690 44.500 ;
        RECT 48.000 44.300 48.690 44.440 ;
        RECT 31.900 44.100 32.040 44.300 ;
        RECT 43.310 44.240 43.630 44.300 ;
        RECT 45.625 44.255 45.915 44.300 ;
        RECT 47.450 44.240 47.770 44.300 ;
        RECT 48.370 44.240 48.690 44.300 ;
        RECT 19.940 43.960 32.040 44.100 ;
        RECT 56.650 44.100 56.970 44.160 ;
        RECT 58.030 44.100 58.350 44.160 ;
        RECT 59.040 44.100 59.180 44.640 ;
        RECT 59.410 44.640 62.015 44.780 ;
        RECT 59.410 44.580 59.730 44.640 ;
        RECT 61.725 44.595 62.015 44.640 ;
        RECT 62.185 44.780 62.475 44.825 ;
        RECT 62.185 44.640 62.585 44.780 ;
        RECT 62.185 44.595 62.475 44.640 ;
        RECT 64.025 44.595 64.315 44.825 ;
        RECT 61.800 44.440 61.940 44.595 ;
        RECT 64.100 44.440 64.240 44.595 ;
        RECT 72.750 44.580 73.070 44.840 ;
        RECT 75.600 44.440 75.740 44.920 ;
        RECT 77.350 44.780 77.670 44.840 ;
        RECT 83.330 44.780 83.650 44.840 ;
        RECT 77.350 44.640 83.650 44.780 ;
        RECT 77.350 44.580 77.670 44.640 ;
        RECT 83.330 44.580 83.650 44.640 ;
        RECT 83.790 44.580 84.110 44.840 ;
        RECT 85.260 44.825 85.400 44.980 ;
        RECT 86.550 44.920 86.870 45.180 ;
        RECT 88.940 45.120 89.080 45.320 ;
        RECT 88.940 44.980 92.760 45.120 ;
        RECT 84.265 44.595 84.555 44.825 ;
        RECT 85.185 44.595 85.475 44.825 ;
        RECT 85.630 44.780 85.950 44.840 ;
        RECT 86.640 44.780 86.780 44.920 ;
        RECT 87.025 44.780 87.315 44.825 ;
        RECT 85.630 44.640 87.315 44.780 ;
        RECT 61.800 44.300 64.240 44.440 ;
        RECT 64.560 44.300 75.740 44.440 ;
        RECT 81.030 44.440 81.350 44.500 ;
        RECT 83.880 44.440 84.020 44.580 ;
        RECT 81.030 44.300 84.020 44.440 ;
        RECT 84.340 44.440 84.480 44.595 ;
        RECT 85.630 44.580 85.950 44.640 ;
        RECT 87.025 44.595 87.315 44.640 ;
        RECT 87.485 44.595 87.775 44.825 ;
        RECT 86.550 44.440 86.870 44.500 ;
        RECT 84.340 44.300 86.870 44.440 ;
        RECT 56.650 43.960 59.180 44.100 ;
        RECT 59.425 44.100 59.715 44.145 ;
        RECT 60.790 44.100 61.110 44.160 ;
        RECT 64.560 44.100 64.700 44.300 ;
        RECT 81.030 44.240 81.350 44.300 ;
        RECT 59.425 43.960 64.700 44.100 ;
        RECT 56.650 43.900 56.970 43.960 ;
        RECT 58.030 43.900 58.350 43.960 ;
        RECT 59.425 43.915 59.715 43.960 ;
        RECT 60.790 43.900 61.110 43.960 ;
        RECT 64.930 43.900 65.250 44.160 ;
        RECT 69.070 44.100 69.390 44.160 ;
        RECT 79.205 44.100 79.495 44.145 ;
        RECT 83.330 44.100 83.650 44.160 ;
        RECT 69.070 43.960 83.650 44.100 ;
        RECT 83.880 44.100 84.020 44.300 ;
        RECT 86.550 44.240 86.870 44.300 ;
        RECT 87.560 44.100 87.700 44.595 ;
        RECT 87.930 44.580 88.250 44.840 ;
        RECT 88.940 44.825 89.080 44.980 ;
        RECT 88.865 44.595 89.155 44.825 ;
        RECT 90.705 44.595 90.995 44.825 ;
        RECT 90.780 44.440 90.920 44.595 ;
        RECT 91.150 44.580 91.470 44.840 ;
        RECT 91.610 44.580 91.930 44.840 ;
        RECT 92.620 44.825 92.760 44.980 ;
        RECT 92.545 44.595 92.835 44.825 ;
        RECT 96.210 44.580 96.530 44.840 ;
        RECT 90.780 44.300 91.380 44.440 ;
        RECT 91.240 44.160 91.380 44.300 ;
        RECT 83.880 43.960 87.700 44.100 ;
        RECT 69.070 43.900 69.390 43.960 ;
        RECT 79.205 43.915 79.495 43.960 ;
        RECT 83.330 43.900 83.650 43.960 ;
        RECT 91.150 43.900 91.470 44.160 ;
        RECT 5.520 43.280 113.620 43.760 ;
        RECT 20.325 43.080 20.615 43.125 ;
        RECT 22.610 43.080 22.930 43.140 ;
        RECT 20.325 42.940 22.930 43.080 ;
        RECT 20.325 42.895 20.615 42.940 ;
        RECT 22.610 42.880 22.930 42.940 ;
        RECT 24.005 43.080 24.295 43.125 ;
        RECT 29.050 43.080 29.370 43.140 ;
        RECT 24.005 42.940 29.370 43.080 ;
        RECT 24.005 42.895 24.295 42.940 ;
        RECT 29.050 42.880 29.370 42.940 ;
        RECT 29.510 42.880 29.830 43.140 ;
        RECT 31.825 43.080 32.115 43.125 ;
        RECT 32.270 43.080 32.590 43.140 ;
        RECT 42.390 43.080 42.710 43.140 ;
        RECT 31.825 42.940 32.590 43.080 ;
        RECT 31.825 42.895 32.115 42.940 ;
        RECT 32.270 42.880 32.590 42.940 ;
        RECT 35.120 42.940 42.710 43.080 ;
        RECT 20.400 42.600 28.360 42.740 ;
        RECT 17.105 42.215 17.395 42.445 ;
        RECT 17.180 42.060 17.320 42.215 ;
        RECT 18.010 42.200 18.330 42.460 ;
        RECT 18.485 42.215 18.775 42.445 ;
        RECT 18.945 42.400 19.235 42.445 ;
        RECT 20.400 42.400 20.540 42.600 ;
        RECT 18.945 42.260 20.540 42.400 ;
        RECT 18.945 42.215 19.235 42.260 ;
        RECT 17.180 41.920 18.240 42.060 ;
        RECT 18.100 41.380 18.240 41.920 ;
        RECT 18.560 41.720 18.700 42.215 ;
        RECT 20.770 42.200 21.090 42.460 ;
        RECT 22.700 42.445 22.840 42.600 ;
        RECT 28.220 42.460 28.360 42.600 ;
        RECT 21.705 42.215 21.995 42.445 ;
        RECT 22.165 42.215 22.455 42.445 ;
        RECT 22.625 42.215 22.915 42.445 ;
        RECT 19.390 42.060 19.710 42.120 ;
        RECT 21.780 42.060 21.920 42.215 ;
        RECT 19.390 41.920 21.920 42.060 ;
        RECT 19.390 41.860 19.710 41.920 ;
        RECT 22.240 41.720 22.380 42.215 ;
        RECT 26.290 42.200 26.610 42.460 ;
        RECT 27.225 42.215 27.515 42.445 ;
        RECT 27.685 42.215 27.975 42.445 ;
        RECT 28.130 42.400 28.450 42.460 ;
        RECT 33.190 42.400 33.510 42.460 ;
        RECT 28.130 42.260 33.510 42.400 ;
        RECT 23.530 42.060 23.850 42.120 ;
        RECT 27.300 42.060 27.440 42.215 ;
        RECT 23.530 41.920 27.440 42.060 ;
        RECT 27.760 42.060 27.900 42.215 ;
        RECT 28.130 42.200 28.450 42.260 ;
        RECT 33.190 42.200 33.510 42.260 ;
        RECT 33.650 42.200 33.970 42.460 ;
        RECT 34.110 42.200 34.430 42.460 ;
        RECT 35.120 42.445 35.260 42.940 ;
        RECT 42.390 42.880 42.710 42.940 ;
        RECT 51.605 43.080 51.895 43.125 ;
        RECT 52.050 43.080 52.370 43.140 ;
        RECT 51.605 42.940 52.370 43.080 ;
        RECT 51.605 42.895 51.895 42.940 ;
        RECT 52.050 42.880 52.370 42.940 ;
        RECT 55.285 43.080 55.575 43.125 ;
        RECT 57.570 43.080 57.890 43.140 ;
        RECT 55.285 42.940 57.890 43.080 ;
        RECT 55.285 42.895 55.575 42.940 ;
        RECT 57.570 42.880 57.890 42.940 ;
        RECT 58.030 43.080 58.350 43.140 ;
        RECT 61.250 43.080 61.570 43.140 ;
        RECT 64.930 43.080 65.250 43.140 ;
        RECT 91.150 43.080 91.470 43.140 ;
        RECT 58.030 42.940 58.720 43.080 ;
        RECT 58.030 42.880 58.350 42.940 ;
        RECT 38.250 42.540 38.570 42.800 ;
        RECT 46.990 42.540 47.310 42.800 ;
        RECT 50.670 42.740 50.990 42.800 ;
        RECT 58.580 42.740 58.720 42.940 ;
        RECT 61.250 42.940 91.470 43.080 ;
        RECT 61.250 42.880 61.570 42.940 ;
        RECT 64.930 42.880 65.250 42.940 ;
        RECT 91.150 42.880 91.470 42.940 ;
        RECT 92.070 43.080 92.390 43.140 ;
        RECT 92.545 43.080 92.835 43.125 ;
        RECT 104.965 43.080 105.255 43.125 ;
        RECT 92.070 42.940 92.835 43.080 ;
        RECT 92.070 42.880 92.390 42.940 ;
        RECT 92.545 42.895 92.835 42.940 ;
        RECT 95.380 42.940 105.255 43.080 ;
        RECT 62.185 42.740 62.475 42.785 ;
        RECT 50.300 42.600 54.120 42.740 ;
        RECT 58.580 42.600 62.475 42.740 ;
        RECT 35.045 42.215 35.335 42.445 ;
        RECT 35.505 42.400 35.795 42.445 ;
        RECT 43.310 42.400 43.630 42.460 ;
        RECT 35.505 42.260 43.630 42.400 ;
        RECT 35.505 42.215 35.795 42.260 ;
        RECT 29.050 42.060 29.370 42.120 ;
        RECT 33.740 42.060 33.880 42.200 ;
        RECT 27.760 41.920 33.880 42.060 ;
        RECT 23.530 41.860 23.850 41.920 ;
        RECT 27.760 41.720 27.900 41.920 ;
        RECT 29.050 41.860 29.370 41.920 ;
        RECT 18.560 41.580 27.900 41.720 ;
        RECT 29.510 41.720 29.830 41.780 ;
        RECT 35.120 41.720 35.260 42.215 ;
        RECT 43.310 42.200 43.630 42.260 ;
        RECT 48.370 42.200 48.690 42.460 ;
        RECT 49.290 42.200 49.610 42.460 ;
        RECT 49.750 42.200 50.070 42.460 ;
        RECT 50.300 42.445 50.440 42.600 ;
        RECT 50.670 42.540 50.990 42.600 ;
        RECT 53.980 42.460 54.120 42.600 ;
        RECT 62.185 42.555 62.475 42.600 ;
        RECT 66.310 42.540 66.630 42.800 ;
        RECT 68.605 42.740 69.255 42.785 ;
        RECT 72.205 42.740 72.495 42.785 ;
        RECT 68.605 42.600 72.495 42.740 ;
        RECT 68.605 42.555 69.255 42.600 ;
        RECT 71.905 42.555 72.495 42.600 ;
        RECT 77.350 42.740 77.670 42.800 ;
        RECT 81.030 42.740 81.350 42.800 ;
        RECT 77.350 42.600 79.880 42.740 ;
        RECT 71.905 42.460 72.195 42.555 ;
        RECT 77.350 42.540 77.670 42.600 ;
        RECT 79.740 42.460 79.880 42.600 ;
        RECT 80.200 42.600 81.350 42.740 ;
        RECT 50.225 42.215 50.515 42.445 ;
        RECT 52.050 42.200 52.370 42.460 ;
        RECT 52.985 42.215 53.275 42.445 ;
        RECT 46.990 42.060 47.310 42.120 ;
        RECT 53.060 42.060 53.200 42.215 ;
        RECT 53.430 42.200 53.750 42.460 ;
        RECT 53.890 42.200 54.210 42.460 ;
        RECT 58.490 42.200 58.810 42.460 ;
        RECT 59.410 42.400 59.730 42.460 ;
        RECT 59.885 42.400 60.175 42.445 ;
        RECT 59.410 42.260 60.175 42.400 ;
        RECT 59.410 42.200 59.730 42.260 ;
        RECT 59.885 42.215 60.175 42.260 ;
        RECT 65.410 42.400 65.700 42.445 ;
        RECT 67.245 42.400 67.535 42.445 ;
        RECT 70.825 42.400 71.115 42.445 ;
        RECT 65.410 42.260 71.115 42.400 ;
        RECT 65.410 42.215 65.700 42.260 ;
        RECT 67.245 42.215 67.535 42.260 ;
        RECT 70.825 42.215 71.115 42.260 ;
        RECT 71.830 42.240 72.195 42.460 ;
        RECT 71.830 42.200 72.150 42.240 ;
        RECT 75.970 42.200 76.290 42.460 ;
        RECT 76.445 42.400 76.735 42.445 ;
        RECT 76.445 42.260 77.580 42.400 ;
        RECT 76.445 42.215 76.735 42.260 ;
        RECT 46.990 41.920 53.200 42.060 ;
        RECT 46.990 41.860 47.310 41.920 ;
        RECT 29.510 41.580 35.260 41.720 ;
        RECT 35.490 41.720 35.810 41.780 ;
        RECT 35.965 41.720 36.255 41.765 ;
        RECT 35.490 41.580 36.255 41.720 ;
        RECT 29.510 41.520 29.830 41.580 ;
        RECT 35.490 41.520 35.810 41.580 ;
        RECT 35.965 41.535 36.255 41.580 ;
        RECT 49.750 41.720 50.070 41.780 ;
        RECT 53.520 41.720 53.660 42.200 ;
        RECT 56.650 42.060 56.970 42.120 ;
        RECT 58.045 42.060 58.335 42.105 ;
        RECT 61.250 42.060 61.570 42.120 ;
        RECT 56.650 41.920 61.570 42.060 ;
        RECT 56.650 41.860 56.970 41.920 ;
        RECT 58.045 41.875 58.335 41.920 ;
        RECT 61.250 41.860 61.570 41.920 ;
        RECT 64.945 42.060 65.235 42.105 ;
        RECT 69.070 42.060 69.390 42.120 ;
        RECT 64.945 41.920 69.390 42.060 ;
        RECT 64.945 41.875 65.235 41.920 ;
        RECT 69.070 41.860 69.390 41.920 ;
        RECT 73.670 42.060 73.990 42.120 ;
        RECT 76.520 42.060 76.660 42.215 ;
        RECT 73.670 41.920 76.660 42.060 ;
        RECT 73.670 41.860 73.990 41.920 ;
        RECT 76.905 41.875 77.195 42.105 ;
        RECT 77.440 42.060 77.580 42.260 ;
        RECT 79.650 42.200 79.970 42.460 ;
        RECT 80.200 42.445 80.340 42.600 ;
        RECT 81.030 42.540 81.350 42.600 ;
        RECT 87.005 42.740 87.655 42.785 ;
        RECT 89.770 42.740 90.090 42.800 ;
        RECT 90.605 42.740 90.895 42.785 ;
        RECT 87.005 42.600 90.895 42.740 ;
        RECT 87.005 42.555 87.655 42.600 ;
        RECT 89.770 42.540 90.090 42.600 ;
        RECT 90.305 42.555 90.895 42.600 ;
        RECT 80.125 42.215 80.415 42.445 ;
        RECT 80.585 42.215 80.875 42.445 ;
        RECT 80.660 42.060 80.800 42.215 ;
        RECT 81.490 42.200 81.810 42.460 ;
        RECT 83.330 42.200 83.650 42.460 ;
        RECT 83.810 42.400 84.100 42.445 ;
        RECT 85.645 42.400 85.935 42.445 ;
        RECT 89.225 42.400 89.515 42.445 ;
        RECT 83.810 42.260 89.515 42.400 ;
        RECT 83.810 42.215 84.100 42.260 ;
        RECT 85.645 42.215 85.935 42.260 ;
        RECT 89.225 42.215 89.515 42.260 ;
        RECT 90.305 42.240 90.595 42.555 ;
        RECT 91.240 42.400 91.380 42.880 ;
        RECT 93.925 42.400 94.215 42.445 ;
        RECT 91.240 42.260 94.215 42.400 ;
        RECT 93.925 42.215 94.215 42.260 ;
        RECT 94.370 42.200 94.690 42.460 ;
        RECT 94.830 42.400 95.150 42.460 ;
        RECT 95.380 42.400 95.520 42.940 ;
        RECT 104.965 42.895 105.255 42.940 ;
        RECT 99.885 42.740 100.535 42.785 ;
        RECT 103.485 42.740 103.775 42.785 ;
        RECT 105.885 42.740 106.175 42.785 ;
        RECT 99.885 42.600 106.175 42.740 ;
        RECT 99.885 42.555 100.535 42.600 ;
        RECT 103.185 42.555 103.775 42.600 ;
        RECT 105.885 42.555 106.175 42.600 ;
        RECT 94.830 42.260 95.520 42.400 ;
        RECT 94.830 42.200 95.150 42.260 ;
        RECT 95.750 42.200 96.070 42.460 ;
        RECT 96.690 42.400 96.980 42.445 ;
        RECT 98.525 42.400 98.815 42.445 ;
        RECT 102.105 42.400 102.395 42.445 ;
        RECT 96.690 42.260 102.395 42.400 ;
        RECT 96.690 42.215 96.980 42.260 ;
        RECT 98.525 42.215 98.815 42.260 ;
        RECT 102.105 42.215 102.395 42.260 ;
        RECT 103.185 42.240 103.475 42.555 ;
        RECT 105.425 42.215 105.715 42.445 ;
        RECT 77.440 41.920 80.800 42.060 ;
        RECT 49.750 41.580 53.660 41.720 ;
        RECT 59.425 41.720 59.715 41.765 ;
        RECT 62.630 41.720 62.950 41.780 ;
        RECT 59.425 41.580 62.950 41.720 ;
        RECT 49.750 41.520 50.070 41.580 ;
        RECT 59.425 41.535 59.715 41.580 ;
        RECT 62.630 41.520 62.950 41.580 ;
        RECT 63.565 41.720 63.855 41.765 ;
        RECT 65.815 41.720 66.105 41.765 ;
        RECT 67.705 41.720 67.995 41.765 ;
        RECT 70.825 41.720 71.115 41.765 ;
        RECT 76.980 41.720 77.120 41.875 ;
        RECT 63.565 41.580 65.620 41.720 ;
        RECT 63.565 41.535 63.855 41.580 ;
        RECT 20.770 41.380 21.090 41.440 ;
        RECT 22.610 41.380 22.930 41.440 ;
        RECT 26.290 41.380 26.610 41.440 ;
        RECT 29.600 41.380 29.740 41.520 ;
        RECT 18.100 41.240 29.740 41.380 ;
        RECT 48.370 41.380 48.690 41.440 ;
        RECT 52.050 41.380 52.370 41.440 ;
        RECT 60.790 41.380 61.110 41.440 ;
        RECT 48.370 41.240 61.110 41.380 ;
        RECT 65.480 41.380 65.620 41.580 ;
        RECT 65.815 41.580 71.115 41.720 ;
        RECT 65.815 41.535 66.105 41.580 ;
        RECT 67.705 41.535 67.995 41.580 ;
        RECT 70.825 41.535 71.115 41.580 ;
        RECT 73.300 41.580 77.120 41.720 ;
        RECT 78.730 41.720 79.050 41.780 ;
        RECT 81.580 41.720 81.720 42.200 ;
        RECT 84.710 41.860 85.030 42.120 ;
        RECT 87.470 42.060 87.790 42.120 ;
        RECT 96.225 42.060 96.515 42.105 ;
        RECT 87.470 41.920 96.515 42.060 ;
        RECT 87.470 41.860 87.790 41.920 ;
        RECT 96.225 41.875 96.515 41.920 ;
        RECT 97.590 41.860 97.910 42.120 ;
        RECT 105.500 42.060 105.640 42.215 ;
        RECT 103.200 41.920 105.640 42.060 ;
        RECT 103.200 41.780 103.340 41.920 ;
        RECT 78.730 41.580 81.720 41.720 ;
        RECT 84.215 41.720 84.505 41.765 ;
        RECT 86.105 41.720 86.395 41.765 ;
        RECT 89.225 41.720 89.515 41.765 ;
        RECT 95.750 41.720 96.070 41.780 ;
        RECT 84.215 41.580 89.515 41.720 ;
        RECT 73.300 41.440 73.440 41.580 ;
        RECT 78.730 41.520 79.050 41.580 ;
        RECT 84.215 41.535 84.505 41.580 ;
        RECT 86.105 41.535 86.395 41.580 ;
        RECT 89.225 41.535 89.515 41.580 ;
        RECT 91.700 41.580 96.070 41.720 ;
        RECT 73.210 41.380 73.530 41.440 ;
        RECT 65.480 41.240 73.530 41.380 ;
        RECT 20.770 41.180 21.090 41.240 ;
        RECT 22.610 41.180 22.930 41.240 ;
        RECT 26.290 41.180 26.610 41.240 ;
        RECT 48.370 41.180 48.690 41.240 ;
        RECT 52.050 41.180 52.370 41.240 ;
        RECT 60.790 41.180 61.110 41.240 ;
        RECT 73.210 41.180 73.530 41.240 ;
        RECT 74.130 41.180 74.450 41.440 ;
        RECT 78.270 41.180 78.590 41.440 ;
        RECT 82.870 41.380 83.190 41.440 ;
        RECT 88.390 41.380 88.710 41.440 ;
        RECT 91.700 41.380 91.840 41.580 ;
        RECT 95.750 41.520 96.070 41.580 ;
        RECT 97.095 41.720 97.385 41.765 ;
        RECT 98.985 41.720 99.275 41.765 ;
        RECT 102.105 41.720 102.395 41.765 ;
        RECT 97.095 41.580 102.395 41.720 ;
        RECT 97.095 41.535 97.385 41.580 ;
        RECT 98.985 41.535 99.275 41.580 ;
        RECT 102.105 41.535 102.395 41.580 ;
        RECT 103.110 41.520 103.430 41.780 ;
        RECT 82.870 41.240 91.840 41.380 ;
        RECT 82.870 41.180 83.190 41.240 ;
        RECT 88.390 41.180 88.710 41.240 ;
        RECT 92.070 41.180 92.390 41.440 ;
        RECT 5.520 40.560 113.620 41.040 ;
        RECT 23.070 40.360 23.390 40.420 ;
        RECT 25.845 40.360 26.135 40.405 ;
        RECT 23.070 40.220 26.135 40.360 ;
        RECT 23.070 40.160 23.390 40.220 ;
        RECT 25.845 40.175 26.135 40.220 ;
        RECT 52.050 40.160 52.370 40.420 ;
        RECT 59.870 40.360 60.190 40.420 ;
        RECT 60.805 40.360 61.095 40.405 ;
        RECT 59.870 40.220 61.095 40.360 ;
        RECT 59.870 40.160 60.190 40.220 ;
        RECT 60.805 40.175 61.095 40.220 ;
        RECT 61.250 40.360 61.570 40.420 ;
        RECT 65.405 40.360 65.695 40.405 ;
        RECT 61.250 40.220 65.695 40.360 ;
        RECT 61.250 40.160 61.570 40.220 ;
        RECT 65.405 40.175 65.695 40.220 ;
        RECT 66.310 40.360 66.630 40.420 ;
        RECT 67.705 40.360 67.995 40.405 ;
        RECT 66.310 40.220 67.995 40.360 ;
        RECT 66.310 40.160 66.630 40.220 ;
        RECT 67.705 40.175 67.995 40.220 ;
        RECT 70.925 40.360 71.215 40.405 ;
        RECT 71.830 40.360 72.150 40.420 ;
        RECT 70.925 40.220 72.150 40.360 ;
        RECT 70.925 40.175 71.215 40.220 ;
        RECT 71.830 40.160 72.150 40.220 ;
        RECT 81.490 40.160 81.810 40.420 ;
        RECT 84.710 40.360 85.030 40.420 ;
        RECT 86.565 40.360 86.855 40.405 ;
        RECT 84.710 40.220 86.855 40.360 ;
        RECT 84.710 40.160 85.030 40.220 ;
        RECT 86.565 40.175 86.855 40.220 ;
        RECT 91.165 40.360 91.455 40.405 ;
        RECT 96.670 40.360 96.990 40.420 ;
        RECT 91.165 40.220 96.990 40.360 ;
        RECT 91.165 40.175 91.455 40.220 ;
        RECT 96.670 40.160 96.990 40.220 ;
        RECT 19.850 40.020 20.170 40.080 ;
        RECT 26.305 40.020 26.595 40.065 ;
        RECT 19.850 39.880 26.595 40.020 ;
        RECT 19.850 39.820 20.170 39.880 ;
        RECT 26.305 39.835 26.595 39.880 ;
        RECT 31.315 40.020 31.605 40.065 ;
        RECT 33.205 40.020 33.495 40.065 ;
        RECT 36.325 40.020 36.615 40.065 ;
        RECT 72.305 40.020 72.595 40.065 ;
        RECT 31.315 39.880 36.615 40.020 ;
        RECT 31.315 39.835 31.605 39.880 ;
        RECT 33.205 39.835 33.495 39.880 ;
        RECT 36.325 39.835 36.615 39.880 ;
        RECT 66.400 39.880 72.595 40.020 ;
        RECT 29.050 39.680 29.370 39.740 ;
        RECT 24.080 39.540 29.370 39.680 ;
        RECT 12.505 39.340 12.795 39.385 ;
        RECT 13.410 39.340 13.730 39.400 ;
        RECT 12.505 39.200 13.730 39.340 ;
        RECT 12.505 39.155 12.795 39.200 ;
        RECT 13.410 39.140 13.730 39.200 ;
        RECT 13.870 39.140 14.190 39.400 ;
        RECT 15.265 39.340 15.555 39.385 ;
        RECT 16.645 39.340 16.935 39.385 ;
        RECT 17.550 39.340 17.870 39.400 ;
        RECT 15.265 39.200 17.870 39.340 ;
        RECT 15.265 39.155 15.555 39.200 ;
        RECT 16.645 39.155 16.935 39.200 ;
        RECT 17.550 39.140 17.870 39.200 ;
        RECT 22.610 39.140 22.930 39.400 ;
        RECT 24.080 39.385 24.220 39.540 ;
        RECT 23.545 39.155 23.835 39.385 ;
        RECT 24.005 39.155 24.295 39.385 ;
        RECT 24.465 39.340 24.755 39.385 ;
        RECT 27.670 39.340 27.990 39.400 ;
        RECT 28.220 39.385 28.360 39.540 ;
        RECT 29.050 39.480 29.370 39.540 ;
        RECT 30.445 39.680 30.735 39.725 ;
        RECT 38.250 39.680 38.570 39.740 ;
        RECT 30.445 39.540 38.570 39.680 ;
        RECT 30.445 39.495 30.735 39.540 ;
        RECT 38.250 39.480 38.570 39.540 ;
        RECT 39.260 39.540 46.760 39.680 ;
        RECT 24.465 39.200 27.990 39.340 ;
        RECT 24.465 39.155 24.755 39.200 ;
        RECT 21.230 39.000 21.550 39.060 ;
        RECT 23.620 39.000 23.760 39.155 ;
        RECT 27.670 39.140 27.990 39.200 ;
        RECT 28.145 39.155 28.435 39.385 ;
        RECT 28.605 39.155 28.895 39.385 ;
        RECT 21.230 38.860 23.760 39.000 ;
        RECT 27.210 39.000 27.530 39.060 ;
        RECT 28.680 39.000 28.820 39.155 ;
        RECT 29.510 39.140 29.830 39.400 ;
        RECT 30.910 39.340 31.200 39.385 ;
        RECT 32.745 39.340 33.035 39.385 ;
        RECT 36.325 39.340 36.615 39.385 ;
        RECT 30.910 39.200 36.615 39.340 ;
        RECT 30.910 39.155 31.200 39.200 ;
        RECT 32.745 39.155 33.035 39.200 ;
        RECT 36.325 39.155 36.615 39.200 ;
        RECT 27.210 38.860 28.820 39.000 ;
        RECT 29.970 39.000 30.290 39.060 ;
        RECT 31.825 39.000 32.115 39.045 ;
        RECT 29.970 38.860 32.115 39.000 ;
        RECT 21.230 38.800 21.550 38.860 ;
        RECT 27.210 38.800 27.530 38.860 ;
        RECT 29.970 38.800 30.290 38.860 ;
        RECT 31.825 38.815 32.115 38.860 ;
        RECT 34.105 39.000 34.755 39.045 ;
        RECT 35.490 39.000 35.810 39.060 ;
        RECT 37.405 39.045 37.695 39.360 ;
        RECT 37.405 39.000 37.995 39.045 ;
        RECT 34.105 38.860 37.995 39.000 ;
        RECT 34.105 38.815 34.755 38.860 ;
        RECT 35.490 38.800 35.810 38.860 ;
        RECT 37.705 38.815 37.995 38.860 ;
        RECT 39.260 38.720 39.400 39.540 ;
        RECT 46.620 39.385 46.760 39.540 ;
        RECT 46.990 39.480 47.310 39.740 ;
        RECT 47.925 39.680 48.215 39.725 ;
        RECT 51.130 39.680 51.450 39.740 ;
        RECT 52.985 39.680 53.275 39.725 ;
        RECT 47.925 39.540 53.275 39.680 ;
        RECT 47.925 39.495 48.215 39.540 ;
        RECT 51.130 39.480 51.450 39.540 ;
        RECT 52.985 39.495 53.275 39.540 ;
        RECT 57.570 39.680 57.890 39.740 ;
        RECT 58.965 39.680 59.255 39.725 ;
        RECT 57.570 39.540 59.255 39.680 ;
        RECT 57.570 39.480 57.890 39.540 ;
        RECT 58.965 39.495 59.255 39.540 ;
        RECT 59.425 39.680 59.715 39.725 ;
        RECT 61.250 39.680 61.570 39.740 ;
        RECT 59.425 39.540 61.020 39.680 ;
        RECT 59.425 39.495 59.715 39.540 ;
        RECT 41.485 39.340 41.775 39.385 ;
        RECT 41.485 39.200 44.920 39.340 ;
        RECT 41.485 39.155 41.775 39.200 ;
        RECT 9.730 38.660 10.050 38.720 ;
        RECT 11.585 38.660 11.875 38.705 ;
        RECT 9.730 38.520 11.875 38.660 ;
        RECT 9.730 38.460 10.050 38.520 ;
        RECT 11.585 38.475 11.875 38.520 ;
        RECT 12.950 38.460 13.270 38.720 ;
        RECT 14.790 38.460 15.110 38.720 ;
        RECT 15.710 38.660 16.030 38.720 ;
        RECT 16.185 38.660 16.475 38.705 ;
        RECT 15.710 38.520 16.475 38.660 ;
        RECT 15.710 38.460 16.030 38.520 ;
        RECT 16.185 38.475 16.475 38.520 ;
        RECT 39.170 38.460 39.490 38.720 ;
        RECT 39.630 38.660 39.950 38.720 ;
        RECT 44.780 38.705 44.920 39.200 ;
        RECT 46.545 39.155 46.835 39.385 ;
        RECT 48.370 39.340 48.690 39.400 ;
        RECT 48.845 39.340 49.135 39.385 ;
        RECT 48.370 39.200 49.135 39.340 ;
        RECT 46.620 39.000 46.760 39.155 ;
        RECT 48.370 39.140 48.690 39.200 ;
        RECT 48.845 39.155 49.135 39.200 ;
        RECT 49.765 39.155 50.055 39.385 ;
        RECT 49.840 39.000 49.980 39.155 ;
        RECT 50.210 39.140 50.530 39.400 ;
        RECT 50.670 39.140 50.990 39.400 ;
        RECT 54.365 39.340 54.655 39.385 ;
        RECT 58.030 39.340 58.350 39.400 ;
        RECT 54.365 39.200 58.350 39.340 ;
        RECT 54.365 39.155 54.655 39.200 ;
        RECT 58.030 39.140 58.350 39.200 ;
        RECT 58.490 39.140 58.810 39.400 ;
        RECT 59.870 39.140 60.190 39.400 ;
        RECT 60.880 39.340 61.020 39.540 ;
        RECT 61.250 39.540 66.080 39.680 ;
        RECT 61.250 39.480 61.570 39.540 ;
        RECT 62.170 39.340 62.490 39.400 ;
        RECT 60.880 39.200 62.490 39.340 ;
        RECT 62.170 39.140 62.490 39.200 ;
        RECT 64.470 39.140 64.790 39.400 ;
        RECT 65.940 39.385 66.080 39.540 ;
        RECT 66.400 39.385 66.540 39.880 ;
        RECT 72.305 39.835 72.595 39.880 ;
        RECT 73.210 40.020 73.530 40.080 ;
        RECT 73.210 39.880 83.100 40.020 ;
        RECT 73.210 39.820 73.530 39.880 ;
        RECT 75.140 39.740 75.280 39.880 ;
        RECT 74.130 39.680 74.450 39.740 ;
        RECT 68.700 39.540 74.450 39.680 ;
        RECT 68.700 39.385 68.840 39.540 ;
        RECT 74.130 39.480 74.450 39.540 ;
        RECT 75.050 39.480 75.370 39.740 ;
        RECT 81.030 39.680 81.350 39.740 ;
        RECT 82.960 39.725 83.100 39.880 ;
        RECT 86.090 39.820 86.410 40.080 ;
        RECT 99.545 40.020 99.835 40.065 ;
        RECT 102.665 40.020 102.955 40.065 ;
        RECT 104.555 40.020 104.845 40.065 ;
        RECT 99.545 39.880 104.845 40.020 ;
        RECT 99.545 39.835 99.835 39.880 ;
        RECT 102.665 39.835 102.955 39.880 ;
        RECT 104.555 39.835 104.845 39.880 ;
        RECT 79.740 39.540 81.350 39.680 ;
        RECT 65.865 39.155 66.155 39.385 ;
        RECT 66.325 39.155 66.615 39.385 ;
        RECT 68.625 39.155 68.915 39.385 ;
        RECT 71.385 39.340 71.675 39.385 ;
        RECT 72.290 39.340 72.610 39.400 ;
        RECT 71.385 39.200 72.610 39.340 ;
        RECT 71.385 39.155 71.675 39.200 ;
        RECT 72.290 39.140 72.610 39.200 ;
        RECT 78.285 39.340 78.575 39.385 ;
        RECT 78.730 39.340 79.050 39.400 ;
        RECT 79.740 39.385 79.880 39.540 ;
        RECT 81.030 39.480 81.350 39.540 ;
        RECT 82.885 39.495 83.175 39.725 ;
        RECT 83.805 39.680 84.095 39.725 ;
        RECT 83.805 39.540 91.840 39.680 ;
        RECT 83.805 39.495 84.095 39.540 ;
        RECT 78.285 39.200 79.050 39.340 ;
        RECT 78.285 39.155 78.575 39.200 ;
        RECT 78.730 39.140 79.050 39.200 ;
        RECT 79.205 39.155 79.495 39.385 ;
        RECT 79.665 39.155 79.955 39.385 ;
        RECT 46.620 38.860 49.980 39.000 ;
        RECT 63.090 38.800 63.410 39.060 ;
        RECT 73.670 39.000 73.990 39.060 ;
        RECT 74.145 39.000 74.435 39.045 ;
        RECT 79.280 39.000 79.420 39.155 ;
        RECT 80.110 39.140 80.430 39.400 ;
        RECT 86.090 39.340 86.410 39.400 ;
        RECT 87.485 39.340 87.775 39.385 ;
        RECT 86.090 39.200 87.775 39.340 ;
        RECT 86.090 39.140 86.410 39.200 ;
        RECT 87.485 39.155 87.775 39.200 ;
        RECT 87.945 39.340 88.235 39.385 ;
        RECT 88.390 39.340 88.710 39.400 ;
        RECT 87.945 39.200 88.710 39.340 ;
        RECT 87.945 39.155 88.235 39.200 ;
        RECT 88.390 39.140 88.710 39.200 ;
        RECT 88.850 39.140 89.170 39.400 ;
        RECT 89.310 39.140 89.630 39.400 ;
        RECT 89.785 39.340 90.075 39.385 ;
        RECT 91.150 39.340 91.470 39.400 ;
        RECT 89.785 39.200 91.470 39.340 ;
        RECT 91.700 39.340 91.840 39.540 ;
        RECT 92.530 39.480 92.850 39.740 ;
        RECT 93.005 39.680 93.295 39.725 ;
        RECT 94.830 39.680 95.150 39.740 ;
        RECT 93.005 39.540 95.150 39.680 ;
        RECT 93.005 39.495 93.295 39.540 ;
        RECT 94.830 39.480 95.150 39.540 ;
        RECT 102.190 39.680 102.510 39.740 ;
        RECT 105.425 39.680 105.715 39.725 ;
        RECT 102.190 39.540 105.715 39.680 ;
        RECT 102.190 39.480 102.510 39.540 ;
        RECT 105.425 39.495 105.715 39.540 ;
        RECT 92.070 39.340 92.390 39.400 ;
        RECT 93.465 39.340 93.755 39.385 ;
        RECT 91.700 39.200 93.755 39.340 ;
        RECT 89.785 39.155 90.075 39.200 ;
        RECT 91.150 39.140 91.470 39.200 ;
        RECT 92.070 39.140 92.390 39.200 ;
        RECT 93.465 39.155 93.755 39.200 ;
        RECT 98.465 39.045 98.755 39.360 ;
        RECT 99.545 39.340 99.835 39.385 ;
        RECT 103.125 39.340 103.415 39.385 ;
        RECT 104.960 39.340 105.250 39.385 ;
        RECT 99.545 39.200 105.250 39.340 ;
        RECT 99.545 39.155 99.835 39.200 ;
        RECT 103.125 39.155 103.415 39.200 ;
        RECT 104.960 39.155 105.250 39.200 ;
        RECT 73.670 38.860 74.435 39.000 ;
        RECT 73.670 38.800 73.990 38.860 ;
        RECT 74.145 38.815 74.435 38.860 ;
        RECT 77.900 38.860 79.420 39.000 ;
        RECT 98.165 39.000 98.755 39.045 ;
        RECT 101.405 39.000 102.055 39.045 ;
        RECT 102.650 39.000 102.970 39.060 ;
        RECT 98.165 38.860 102.970 39.000 ;
        RECT 77.900 38.720 78.040 38.860 ;
        RECT 98.165 38.815 98.455 38.860 ;
        RECT 101.405 38.815 102.055 38.860 ;
        RECT 102.650 38.800 102.970 38.860 ;
        RECT 104.030 38.800 104.350 39.060 ;
        RECT 40.565 38.660 40.855 38.705 ;
        RECT 39.630 38.520 40.855 38.660 ;
        RECT 39.630 38.460 39.950 38.520 ;
        RECT 40.565 38.475 40.855 38.520 ;
        RECT 44.705 38.475 44.995 38.705 ;
        RECT 67.245 38.660 67.535 38.705 ;
        RECT 70.450 38.660 70.770 38.720 ;
        RECT 67.245 38.520 70.770 38.660 ;
        RECT 67.245 38.475 67.535 38.520 ;
        RECT 70.450 38.460 70.770 38.520 ;
        RECT 74.605 38.660 74.895 38.705 ;
        RECT 77.810 38.660 78.130 38.720 ;
        RECT 74.605 38.520 78.130 38.660 ;
        RECT 74.605 38.475 74.895 38.520 ;
        RECT 77.810 38.460 78.130 38.520 ;
        RECT 82.870 38.660 83.190 38.720 ;
        RECT 84.265 38.660 84.555 38.705 ;
        RECT 87.930 38.660 88.250 38.720 ;
        RECT 82.870 38.520 88.250 38.660 ;
        RECT 82.870 38.460 83.190 38.520 ;
        RECT 84.265 38.475 84.555 38.520 ;
        RECT 87.930 38.460 88.250 38.520 ;
        RECT 93.910 38.660 94.230 38.720 ;
        RECT 95.305 38.660 95.595 38.705 ;
        RECT 93.910 38.520 95.595 38.660 ;
        RECT 93.910 38.460 94.230 38.520 ;
        RECT 95.305 38.475 95.595 38.520 ;
        RECT 96.670 38.460 96.990 38.720 ;
        RECT 5.520 37.840 113.620 38.320 ;
        RECT 13.410 37.640 13.730 37.700 ;
        RECT 17.565 37.640 17.855 37.685 ;
        RECT 13.410 37.500 17.855 37.640 ;
        RECT 13.410 37.440 13.730 37.500 ;
        RECT 17.565 37.455 17.855 37.500 ;
        RECT 19.390 37.440 19.710 37.700 ;
        RECT 29.970 37.440 30.290 37.700 ;
        RECT 34.125 37.640 34.415 37.685 ;
        RECT 39.170 37.640 39.490 37.700 ;
        RECT 34.125 37.500 39.490 37.640 ;
        RECT 34.125 37.455 34.415 37.500 ;
        RECT 39.170 37.440 39.490 37.500 ;
        RECT 46.990 37.440 47.310 37.700 ;
        RECT 60.330 37.640 60.650 37.700 ;
        RECT 61.265 37.640 61.555 37.685 ;
        RECT 60.330 37.500 61.555 37.640 ;
        RECT 60.330 37.440 60.650 37.500 ;
        RECT 61.265 37.455 61.555 37.500 ;
        RECT 77.810 37.440 78.130 37.700 ;
        RECT 88.405 37.640 88.695 37.685 ;
        RECT 89.770 37.640 90.090 37.700 ;
        RECT 88.405 37.500 90.090 37.640 ;
        RECT 88.405 37.455 88.695 37.500 ;
        RECT 89.770 37.440 90.090 37.500 ;
        RECT 93.450 37.440 93.770 37.700 ;
        RECT 94.845 37.640 95.135 37.685 ;
        RECT 97.590 37.640 97.910 37.700 ;
        RECT 94.845 37.500 97.910 37.640 ;
        RECT 94.845 37.455 95.135 37.500 ;
        RECT 97.590 37.440 97.910 37.500 ;
        RECT 100.365 37.455 100.655 37.685 ;
        RECT 101.745 37.640 102.035 37.685 ;
        RECT 104.030 37.640 104.350 37.700 ;
        RECT 101.745 37.500 104.350 37.640 ;
        RECT 101.745 37.455 102.035 37.500 ;
        RECT 9.730 37.100 10.050 37.360 ;
        RECT 12.025 37.300 12.675 37.345 ;
        RECT 14.790 37.300 15.110 37.360 ;
        RECT 15.625 37.300 15.915 37.345 ;
        RECT 12.025 37.160 15.915 37.300 ;
        RECT 12.025 37.115 12.675 37.160 ;
        RECT 14.790 37.100 15.110 37.160 ;
        RECT 15.325 37.115 15.915 37.160 ;
        RECT 26.765 37.300 27.055 37.345 ;
        RECT 26.765 37.160 33.880 37.300 ;
        RECT 26.765 37.115 27.055 37.160 ;
        RECT 8.830 36.960 9.120 37.005 ;
        RECT 10.665 36.960 10.955 37.005 ;
        RECT 14.245 36.960 14.535 37.005 ;
        RECT 8.830 36.820 14.535 36.960 ;
        RECT 8.830 36.775 9.120 36.820 ;
        RECT 10.665 36.775 10.955 36.820 ;
        RECT 14.245 36.775 14.535 36.820 ;
        RECT 15.325 36.800 15.615 37.115 ;
        RECT 21.230 36.960 21.550 37.020 ;
        RECT 33.740 37.005 33.880 37.160 ;
        RECT 39.630 37.100 39.950 37.360 ;
        RECT 41.925 37.300 42.575 37.345 ;
        RECT 45.525 37.300 45.815 37.345 ;
        RECT 47.925 37.300 48.215 37.345 ;
        RECT 41.925 37.160 48.215 37.300 ;
        RECT 41.925 37.115 42.575 37.160 ;
        RECT 45.225 37.115 45.815 37.160 ;
        RECT 47.925 37.115 48.215 37.160 ;
        RECT 26.305 36.960 26.595 37.005 ;
        RECT 21.230 36.820 26.595 36.960 ;
        RECT 21.230 36.760 21.550 36.820 ;
        RECT 26.305 36.775 26.595 36.820 ;
        RECT 29.065 36.960 29.355 37.005 ;
        RECT 33.665 36.960 33.955 37.005 ;
        RECT 34.110 36.960 34.430 37.020 ;
        RECT 29.065 36.820 32.040 36.960 ;
        RECT 29.065 36.775 29.355 36.820 ;
        RECT 8.350 36.420 8.670 36.680 ;
        RECT 17.105 36.620 17.395 36.665 ;
        RECT 18.010 36.620 18.330 36.680 ;
        RECT 19.865 36.620 20.155 36.665 ;
        RECT 17.105 36.480 20.155 36.620 ;
        RECT 17.105 36.435 17.395 36.480 ;
        RECT 18.010 36.420 18.330 36.480 ;
        RECT 19.865 36.435 20.155 36.480 ;
        RECT 20.785 36.620 21.075 36.665 ;
        RECT 22.150 36.620 22.470 36.680 ;
        RECT 27.685 36.620 27.975 36.665 ;
        RECT 20.785 36.480 31.580 36.620 ;
        RECT 20.785 36.435 21.075 36.480 ;
        RECT 9.235 36.280 9.525 36.325 ;
        RECT 11.125 36.280 11.415 36.325 ;
        RECT 14.245 36.280 14.535 36.325 ;
        RECT 9.235 36.140 14.535 36.280 ;
        RECT 9.235 36.095 9.525 36.140 ;
        RECT 11.125 36.095 11.415 36.140 ;
        RECT 14.245 36.095 14.535 36.140 ;
        RECT 19.940 35.940 20.080 36.435 ;
        RECT 22.150 36.420 22.470 36.480 ;
        RECT 27.685 36.435 27.975 36.480 ;
        RECT 20.770 35.940 21.090 36.000 ;
        RECT 19.940 35.800 21.090 35.940 ;
        RECT 20.770 35.740 21.090 35.800 ;
        RECT 23.530 35.940 23.850 36.000 ;
        RECT 24.465 35.940 24.755 35.985 ;
        RECT 23.530 35.800 24.755 35.940 ;
        RECT 31.440 35.940 31.580 36.480 ;
        RECT 31.900 36.325 32.040 36.820 ;
        RECT 33.665 36.820 34.430 36.960 ;
        RECT 33.665 36.775 33.955 36.820 ;
        RECT 34.110 36.760 34.430 36.820 ;
        RECT 38.250 36.760 38.570 37.020 ;
        RECT 38.730 36.960 39.020 37.005 ;
        RECT 40.565 36.960 40.855 37.005 ;
        RECT 44.145 36.960 44.435 37.005 ;
        RECT 38.730 36.820 44.435 36.960 ;
        RECT 38.730 36.775 39.020 36.820 ;
        RECT 40.565 36.775 40.855 36.820 ;
        RECT 44.145 36.775 44.435 36.820 ;
        RECT 45.225 36.800 45.515 37.115 ;
        RECT 70.450 37.100 70.770 37.360 ;
        RECT 72.745 37.300 73.395 37.345 ;
        RECT 76.345 37.300 76.635 37.345 ;
        RECT 78.745 37.300 79.035 37.345 ;
        RECT 96.670 37.300 96.990 37.360 ;
        RECT 98.065 37.300 98.355 37.345 ;
        RECT 72.745 37.160 79.035 37.300 ;
        RECT 72.745 37.115 73.395 37.160 ;
        RECT 76.045 37.115 76.635 37.160 ;
        RECT 78.745 37.115 79.035 37.160 ;
        RECT 91.240 37.160 98.355 37.300 ;
        RECT 47.450 36.760 47.770 37.020 ;
        RECT 58.490 36.760 58.810 37.020 ;
        RECT 59.870 36.760 60.190 37.020 ;
        RECT 60.790 36.960 61.110 37.020 ;
        RECT 61.265 36.960 61.555 37.005 ;
        RECT 60.790 36.820 61.555 36.960 ;
        RECT 60.790 36.760 61.110 36.820 ;
        RECT 61.265 36.775 61.555 36.820 ;
        RECT 69.550 36.960 69.840 37.005 ;
        RECT 71.385 36.960 71.675 37.005 ;
        RECT 74.965 36.960 75.255 37.005 ;
        RECT 69.550 36.820 75.255 36.960 ;
        RECT 69.550 36.775 69.840 36.820 ;
        RECT 71.385 36.775 71.675 36.820 ;
        RECT 74.965 36.775 75.255 36.820 ;
        RECT 76.045 36.800 76.335 37.115 ;
        RECT 79.205 36.775 79.495 37.005 ;
        RECT 87.010 36.960 87.330 37.020 ;
        RECT 87.945 36.960 88.235 37.005 ;
        RECT 87.010 36.820 88.235 36.960 ;
        RECT 33.190 36.620 33.510 36.680 ;
        RECT 35.045 36.620 35.335 36.665 ;
        RECT 51.130 36.620 51.450 36.680 ;
        RECT 33.190 36.480 51.450 36.620 ;
        RECT 33.190 36.420 33.510 36.480 ;
        RECT 35.045 36.435 35.335 36.480 ;
        RECT 51.130 36.420 51.450 36.480 ;
        RECT 69.070 36.420 69.390 36.680 ;
        RECT 72.290 36.620 72.610 36.680 ;
        RECT 79.280 36.620 79.420 36.775 ;
        RECT 87.010 36.760 87.330 36.820 ;
        RECT 87.945 36.775 88.235 36.820 ;
        RECT 88.390 36.960 88.710 37.020 ;
        RECT 91.240 37.005 91.380 37.160 ;
        RECT 96.670 37.100 96.990 37.160 ;
        RECT 98.065 37.115 98.355 37.160 ;
        RECT 90.245 36.960 90.535 37.005 ;
        RECT 88.390 36.820 90.535 36.960 ;
        RECT 80.570 36.620 80.890 36.680 ;
        RECT 72.290 36.480 80.890 36.620 ;
        RECT 88.020 36.620 88.160 36.775 ;
        RECT 88.390 36.760 88.710 36.820 ;
        RECT 90.245 36.775 90.535 36.820 ;
        RECT 91.165 36.775 91.455 37.005 ;
        RECT 91.625 36.775 91.915 37.005 ;
        RECT 89.770 36.620 90.090 36.680 ;
        RECT 88.020 36.480 90.090 36.620 ;
        RECT 72.290 36.420 72.610 36.480 ;
        RECT 80.570 36.420 80.890 36.480 ;
        RECT 89.770 36.420 90.090 36.480 ;
        RECT 31.825 36.095 32.115 36.325 ;
        RECT 39.135 36.280 39.425 36.325 ;
        RECT 41.025 36.280 41.315 36.325 ;
        RECT 44.145 36.280 44.435 36.325 ;
        RECT 39.135 36.140 44.435 36.280 ;
        RECT 39.135 36.095 39.425 36.140 ;
        RECT 41.025 36.095 41.315 36.140 ;
        RECT 44.145 36.095 44.435 36.140 ;
        RECT 62.170 36.280 62.490 36.340 ;
        RECT 63.565 36.280 63.855 36.325 ;
        RECT 62.170 36.140 63.855 36.280 ;
        RECT 62.170 36.080 62.490 36.140 ;
        RECT 63.565 36.095 63.855 36.140 ;
        RECT 69.955 36.280 70.245 36.325 ;
        RECT 71.845 36.280 72.135 36.325 ;
        RECT 74.965 36.280 75.255 36.325 ;
        RECT 69.955 36.140 75.255 36.280 ;
        RECT 69.955 36.095 70.245 36.140 ;
        RECT 71.845 36.095 72.135 36.140 ;
        RECT 74.965 36.095 75.255 36.140 ;
        RECT 89.310 36.280 89.630 36.340 ;
        RECT 91.700 36.280 91.840 36.775 ;
        RECT 92.070 36.760 92.390 37.020 ;
        RECT 93.910 36.760 94.230 37.020 ;
        RECT 94.830 36.960 95.150 37.020 ;
        RECT 98.525 36.960 98.815 37.005 ;
        RECT 94.830 36.820 98.815 36.960 ;
        RECT 100.440 36.960 100.580 37.455 ;
        RECT 104.030 37.440 104.350 37.500 ;
        RECT 102.650 37.100 102.970 37.360 ;
        RECT 100.825 36.960 101.115 37.005 ;
        RECT 100.440 36.820 101.115 36.960 ;
        RECT 94.830 36.760 95.150 36.820 ;
        RECT 98.525 36.775 98.815 36.820 ;
        RECT 100.825 36.775 101.115 36.820 ;
        RECT 102.190 36.960 102.510 37.020 ;
        RECT 103.110 36.960 103.430 37.020 ;
        RECT 102.190 36.820 103.430 36.960 ;
        RECT 102.190 36.760 102.510 36.820 ;
        RECT 103.110 36.760 103.430 36.820 ;
        RECT 92.530 36.620 92.850 36.680 ;
        RECT 97.145 36.620 97.435 36.665 ;
        RECT 92.530 36.480 97.435 36.620 ;
        RECT 92.530 36.420 92.850 36.480 ;
        RECT 97.145 36.435 97.435 36.480 ;
        RECT 89.310 36.140 91.840 36.280 ;
        RECT 89.310 36.080 89.630 36.140 ;
        RECT 33.190 35.940 33.510 36.000 ;
        RECT 31.440 35.800 33.510 35.940 ;
        RECT 23.530 35.740 23.850 35.800 ;
        RECT 24.465 35.755 24.755 35.800 ;
        RECT 33.190 35.740 33.510 35.800 ;
        RECT 5.520 35.120 113.620 35.600 ;
        RECT 10.140 34.920 10.430 34.965 ;
        RECT 12.950 34.920 13.270 34.980 ;
        RECT 10.140 34.780 13.270 34.920 ;
        RECT 10.140 34.735 10.430 34.780 ;
        RECT 12.950 34.720 13.270 34.780 ;
        RECT 13.870 34.920 14.190 34.980 ;
        RECT 18.945 34.920 19.235 34.965 ;
        RECT 13.870 34.780 19.235 34.920 ;
        RECT 13.870 34.720 14.190 34.780 ;
        RECT 18.945 34.735 19.235 34.780 ;
        RECT 32.745 34.920 33.035 34.965 ;
        RECT 34.110 34.920 34.430 34.980 ;
        RECT 32.745 34.780 34.430 34.920 ;
        RECT 32.745 34.735 33.035 34.780 ;
        RECT 34.110 34.720 34.430 34.780 ;
        RECT 57.570 34.920 57.890 34.980 ;
        RECT 60.330 34.920 60.650 34.980 ;
        RECT 61.725 34.920 62.015 34.965 ;
        RECT 62.630 34.920 62.950 34.980 ;
        RECT 57.570 34.780 61.020 34.920 ;
        RECT 57.570 34.720 57.890 34.780 ;
        RECT 60.330 34.720 60.650 34.780 ;
        RECT 9.695 34.580 9.985 34.625 ;
        RECT 11.585 34.580 11.875 34.625 ;
        RECT 14.705 34.580 14.995 34.625 ;
        RECT 9.695 34.440 14.995 34.580 ;
        RECT 9.695 34.395 9.985 34.440 ;
        RECT 11.585 34.395 11.875 34.440 ;
        RECT 14.705 34.395 14.995 34.440 ;
        RECT 24.875 34.580 25.165 34.625 ;
        RECT 26.765 34.580 27.055 34.625 ;
        RECT 29.885 34.580 30.175 34.625 ;
        RECT 58.490 34.580 58.810 34.640 ;
        RECT 60.880 34.625 61.020 34.780 ;
        RECT 61.725 34.780 62.950 34.920 ;
        RECT 61.725 34.735 62.015 34.780 ;
        RECT 62.630 34.720 62.950 34.780 ;
        RECT 89.770 34.920 90.090 34.980 ;
        RECT 102.190 34.920 102.510 34.980 ;
        RECT 89.770 34.780 102.510 34.920 ;
        RECT 89.770 34.720 90.090 34.780 ;
        RECT 102.190 34.720 102.510 34.780 ;
        RECT 24.875 34.440 30.175 34.580 ;
        RECT 24.875 34.395 25.165 34.440 ;
        RECT 26.765 34.395 27.055 34.440 ;
        RECT 29.885 34.395 30.175 34.440 ;
        RECT 58.120 34.440 58.810 34.580 ;
        RECT 17.565 34.240 17.855 34.285 ;
        RECT 21.230 34.240 21.550 34.300 ;
        RECT 17.565 34.100 21.550 34.240 ;
        RECT 17.565 34.055 17.855 34.100 ;
        RECT 21.230 34.040 21.550 34.100 ;
        RECT 22.150 34.040 22.470 34.300 ;
        RECT 47.450 34.240 47.770 34.300 ;
        RECT 34.200 34.100 47.770 34.240 ;
        RECT 8.810 33.700 9.130 33.960 ;
        RECT 9.290 33.900 9.580 33.945 ;
        RECT 11.125 33.900 11.415 33.945 ;
        RECT 14.705 33.900 14.995 33.945 ;
        RECT 9.290 33.760 14.995 33.900 ;
        RECT 9.290 33.715 9.580 33.760 ;
        RECT 11.125 33.715 11.415 33.760 ;
        RECT 14.705 33.715 14.995 33.760 ;
        RECT 15.710 33.920 16.030 33.960 ;
        RECT 15.710 33.700 16.075 33.920 ;
        RECT 20.770 33.700 21.090 33.960 ;
        RECT 23.990 33.700 24.310 33.960 ;
        RECT 34.200 33.945 34.340 34.100 ;
        RECT 47.450 34.040 47.770 34.100 ;
        RECT 47.925 34.240 48.215 34.285 ;
        RECT 51.130 34.240 51.450 34.300 ;
        RECT 47.925 34.100 51.450 34.240 ;
        RECT 47.925 34.055 48.215 34.100 ;
        RECT 51.130 34.040 51.450 34.100 ;
        RECT 57.110 34.040 57.430 34.300 ;
        RECT 58.120 34.285 58.260 34.440 ;
        RECT 58.490 34.380 58.810 34.440 ;
        RECT 60.805 34.395 61.095 34.625 ;
        RECT 91.700 34.440 99.200 34.580 ;
        RECT 91.700 34.300 91.840 34.440 ;
        RECT 58.045 34.240 58.335 34.285 ;
        RECT 63.565 34.240 63.855 34.285 ;
        RECT 58.045 34.100 63.855 34.240 ;
        RECT 58.045 34.055 58.335 34.100 ;
        RECT 63.565 34.055 63.855 34.100 ;
        RECT 72.750 34.240 73.070 34.300 ;
        RECT 75.050 34.240 75.370 34.300 ;
        RECT 76.905 34.240 77.195 34.285 ;
        RECT 72.750 34.100 77.195 34.240 ;
        RECT 72.750 34.040 73.070 34.100 ;
        RECT 75.050 34.040 75.370 34.100 ;
        RECT 76.905 34.055 77.195 34.100 ;
        RECT 91.610 34.040 91.930 34.300 ;
        RECT 95.290 34.240 95.610 34.300 ;
        RECT 99.060 34.285 99.200 34.440 ;
        RECT 98.525 34.240 98.815 34.285 ;
        RECT 93.540 34.100 98.815 34.240 ;
        RECT 24.470 33.900 24.760 33.945 ;
        RECT 26.305 33.900 26.595 33.945 ;
        RECT 29.885 33.900 30.175 33.945 ;
        RECT 24.470 33.760 30.175 33.900 ;
        RECT 24.470 33.715 24.760 33.760 ;
        RECT 26.305 33.715 26.595 33.760 ;
        RECT 29.885 33.715 30.175 33.760 ;
        RECT 15.785 33.605 16.075 33.700 ;
        RECT 12.485 33.560 13.135 33.605 ;
        RECT 15.785 33.560 16.375 33.605 ;
        RECT 12.485 33.420 16.375 33.560 ;
        RECT 12.485 33.375 13.135 33.420 ;
        RECT 16.085 33.375 16.375 33.420 ;
        RECT 25.385 33.560 25.675 33.605 ;
        RECT 26.750 33.560 27.070 33.620 ;
        RECT 30.965 33.605 31.255 33.920 ;
        RECT 34.125 33.715 34.415 33.945 ;
        RECT 42.405 33.900 42.695 33.945 ;
        RECT 47.005 33.900 47.295 33.945 ;
        RECT 49.290 33.900 49.610 33.960 ;
        RECT 42.405 33.760 44.920 33.900 ;
        RECT 42.405 33.715 42.695 33.760 ;
        RECT 25.385 33.420 27.070 33.560 ;
        RECT 25.385 33.375 25.675 33.420 ;
        RECT 26.750 33.360 27.070 33.420 ;
        RECT 27.665 33.560 28.315 33.605 ;
        RECT 30.965 33.560 31.555 33.605 ;
        RECT 33.665 33.560 33.955 33.605 ;
        RECT 27.665 33.420 33.955 33.560 ;
        RECT 27.665 33.375 28.315 33.420 ;
        RECT 31.265 33.375 31.555 33.420 ;
        RECT 33.665 33.375 33.955 33.420 ;
        RECT 41.010 33.220 41.330 33.280 ;
        RECT 44.780 33.265 44.920 33.760 ;
        RECT 47.005 33.760 49.610 33.900 ;
        RECT 47.005 33.715 47.295 33.760 ;
        RECT 49.290 33.700 49.610 33.760 ;
        RECT 58.505 33.900 58.795 33.945 ;
        RECT 61.710 33.900 62.030 33.960 ;
        RECT 62.645 33.900 62.935 33.945 ;
        RECT 58.505 33.760 62.935 33.900 ;
        RECT 58.505 33.715 58.795 33.760 ;
        RECT 61.710 33.700 62.030 33.760 ;
        RECT 62.645 33.715 62.935 33.760 ;
        RECT 63.105 33.900 63.395 33.945 ;
        RECT 63.105 33.760 63.780 33.900 ;
        RECT 63.105 33.715 63.395 33.760 ;
        RECT 59.870 33.560 60.190 33.620 ;
        RECT 60.805 33.560 61.095 33.605 ;
        RECT 62.170 33.560 62.490 33.620 ;
        RECT 59.870 33.420 62.490 33.560 ;
        RECT 59.870 33.360 60.190 33.420 ;
        RECT 60.805 33.375 61.095 33.420 ;
        RECT 62.170 33.360 62.490 33.420 ;
        RECT 41.485 33.220 41.775 33.265 ;
        RECT 41.010 33.080 41.775 33.220 ;
        RECT 41.010 33.020 41.330 33.080 ;
        RECT 41.485 33.035 41.775 33.080 ;
        RECT 44.705 33.035 44.995 33.265 ;
        RECT 46.545 33.220 46.835 33.265 ;
        RECT 46.990 33.220 47.310 33.280 ;
        RECT 46.545 33.080 47.310 33.220 ;
        RECT 46.545 33.035 46.835 33.080 ;
        RECT 46.990 33.020 47.310 33.080 ;
        RECT 60.330 33.220 60.650 33.280 ;
        RECT 63.640 33.220 63.780 33.760 ;
        RECT 64.010 33.700 64.330 33.960 ;
        RECT 77.810 33.900 78.130 33.960 ;
        RECT 78.285 33.900 78.575 33.945 ;
        RECT 77.810 33.760 78.575 33.900 ;
        RECT 77.810 33.700 78.130 33.760 ;
        RECT 78.285 33.715 78.575 33.760 ;
        RECT 80.570 33.700 80.890 33.960 ;
        RECT 88.850 33.900 89.170 33.960 ;
        RECT 91.165 33.900 91.455 33.945 ;
        RECT 88.850 33.760 91.455 33.900 ;
        RECT 88.850 33.700 89.170 33.760 ;
        RECT 91.165 33.715 91.455 33.760 ;
        RECT 82.870 33.560 83.190 33.620 ;
        RECT 77.900 33.420 83.190 33.560 ;
        RECT 77.900 33.265 78.040 33.420 ;
        RECT 82.870 33.360 83.190 33.420 ;
        RECT 90.690 33.560 91.010 33.620 ;
        RECT 93.540 33.560 93.680 34.100 ;
        RECT 95.290 34.040 95.610 34.100 ;
        RECT 98.525 34.055 98.815 34.100 ;
        RECT 98.985 34.055 99.275 34.285 ;
        RECT 94.385 33.900 94.675 33.945 ;
        RECT 96.670 33.900 96.990 33.960 ;
        RECT 98.065 33.900 98.355 33.945 ;
        RECT 94.385 33.760 96.440 33.900 ;
        RECT 94.385 33.715 94.675 33.760 ;
        RECT 90.690 33.420 93.680 33.560 ;
        RECT 90.690 33.360 91.010 33.420 ;
        RECT 60.330 33.080 63.780 33.220 ;
        RECT 60.330 33.020 60.650 33.080 ;
        RECT 77.825 33.035 78.115 33.265 ;
        RECT 80.110 33.020 80.430 33.280 ;
        RECT 80.570 33.220 80.890 33.280 ;
        RECT 81.045 33.220 81.335 33.265 ;
        RECT 80.570 33.080 81.335 33.220 ;
        RECT 80.570 33.020 80.890 33.080 ;
        RECT 81.045 33.035 81.335 33.080 ;
        RECT 88.865 33.220 89.155 33.265 ;
        RECT 89.310 33.220 89.630 33.280 ;
        RECT 88.865 33.080 89.630 33.220 ;
        RECT 88.865 33.035 89.155 33.080 ;
        RECT 89.310 33.020 89.630 33.080 ;
        RECT 93.450 33.020 93.770 33.280 ;
        RECT 96.300 33.265 96.440 33.760 ;
        RECT 96.670 33.760 98.355 33.900 ;
        RECT 96.670 33.700 96.990 33.760 ;
        RECT 98.065 33.715 98.355 33.760 ;
        RECT 96.225 33.035 96.515 33.265 ;
        RECT 5.520 32.400 113.620 32.880 ;
        RECT 18.945 32.200 19.235 32.245 ;
        RECT 19.390 32.200 19.710 32.260 ;
        RECT 18.945 32.060 19.710 32.200 ;
        RECT 18.945 32.015 19.235 32.060 ;
        RECT 19.390 32.000 19.710 32.060 ;
        RECT 25.385 32.200 25.675 32.245 ;
        RECT 26.750 32.200 27.070 32.260 ;
        RECT 25.385 32.060 27.070 32.200 ;
        RECT 25.385 32.015 25.675 32.060 ;
        RECT 26.750 32.000 27.070 32.060 ;
        RECT 48.155 32.200 48.445 32.245 ;
        RECT 49.290 32.200 49.610 32.260 ;
        RECT 50.685 32.200 50.975 32.245 ;
        RECT 63.090 32.200 63.410 32.260 ;
        RECT 71.370 32.200 71.690 32.260 ;
        RECT 48.155 32.060 50.975 32.200 ;
        RECT 48.155 32.015 48.445 32.060 ;
        RECT 49.290 32.000 49.610 32.060 ;
        RECT 50.685 32.015 50.975 32.060 ;
        RECT 53.060 32.060 71.690 32.200 ;
        RECT 27.210 31.860 27.530 31.920 ;
        RECT 19.480 31.720 27.530 31.860 ;
        RECT 19.480 31.565 19.620 31.720 ;
        RECT 27.210 31.660 27.530 31.720 ;
        RECT 40.110 31.860 40.400 31.905 ;
        RECT 41.970 31.860 42.260 31.905 ;
        RECT 40.110 31.720 42.260 31.860 ;
        RECT 40.110 31.675 40.400 31.720 ;
        RECT 41.970 31.675 42.260 31.720 ;
        RECT 42.890 31.860 43.180 31.905 ;
        RECT 45.150 31.860 45.470 31.920 ;
        RECT 46.150 31.860 46.440 31.905 ;
        RECT 42.890 31.720 46.440 31.860 ;
        RECT 42.890 31.675 43.180 31.720 ;
        RECT 19.405 31.335 19.695 31.565 ;
        RECT 23.530 31.520 23.850 31.580 ;
        RECT 24.465 31.520 24.755 31.565 ;
        RECT 23.530 31.380 24.755 31.520 ;
        RECT 23.530 31.320 23.850 31.380 ;
        RECT 24.465 31.335 24.755 31.380 ;
        RECT 38.250 31.520 38.570 31.580 ;
        RECT 39.185 31.520 39.475 31.565 ;
        RECT 38.250 31.380 39.475 31.520 ;
        RECT 38.250 31.320 38.570 31.380 ;
        RECT 39.185 31.335 39.475 31.380 ;
        RECT 41.010 31.320 41.330 31.580 ;
        RECT 42.045 31.520 42.260 31.675 ;
        RECT 45.150 31.660 45.470 31.720 ;
        RECT 46.150 31.675 46.440 31.720 ;
        RECT 48.830 31.860 49.150 31.920 ;
        RECT 51.145 31.860 51.435 31.905 ;
        RECT 48.830 31.720 51.435 31.860 ;
        RECT 48.830 31.660 49.150 31.720 ;
        RECT 51.145 31.675 51.435 31.720 ;
        RECT 44.290 31.520 44.580 31.565 ;
        RECT 42.045 31.380 44.580 31.520 ;
        RECT 44.290 31.335 44.580 31.380 ;
        RECT 52.510 31.520 52.830 31.580 ;
        RECT 53.060 31.565 53.200 32.060 ;
        RECT 63.090 32.000 63.410 32.060 ;
        RECT 71.370 32.000 71.690 32.060 ;
        RECT 71.845 32.200 72.135 32.245 ;
        RECT 75.970 32.200 76.290 32.260 ;
        RECT 79.190 32.200 79.510 32.260 ;
        RECT 71.845 32.060 79.510 32.200 ;
        RECT 71.845 32.015 72.135 32.060 ;
        RECT 75.970 32.000 76.290 32.060 ;
        RECT 79.190 32.000 79.510 32.060 ;
        RECT 82.425 32.200 82.715 32.245 ;
        RECT 82.870 32.200 83.190 32.260 ;
        RECT 82.425 32.060 83.190 32.200 ;
        RECT 82.425 32.015 82.715 32.060 ;
        RECT 82.870 32.000 83.190 32.060 ;
        RECT 86.105 32.200 86.395 32.245 ;
        RECT 88.850 32.200 89.170 32.260 ;
        RECT 86.105 32.060 89.170 32.200 ;
        RECT 86.105 32.015 86.395 32.060 ;
        RECT 88.850 32.000 89.170 32.060 ;
        RECT 95.290 32.200 95.610 32.260 ;
        RECT 100.825 32.200 101.115 32.245 ;
        RECT 95.290 32.060 101.115 32.200 ;
        RECT 95.290 32.000 95.610 32.060 ;
        RECT 100.825 32.015 101.115 32.060 ;
        RECT 59.410 31.860 59.730 31.920 ;
        RECT 60.345 31.860 60.635 31.905 ;
        RECT 76.430 31.860 76.750 31.920 ;
        RECT 59.410 31.720 60.635 31.860 ;
        RECT 59.410 31.660 59.730 31.720 ;
        RECT 60.345 31.675 60.635 31.720 ;
        RECT 71.460 31.720 76.750 31.860 ;
        RECT 52.985 31.520 53.275 31.565 ;
        RECT 52.510 31.380 53.275 31.520 ;
        RECT 52.510 31.320 52.830 31.380 ;
        RECT 52.985 31.335 53.275 31.380 ;
        RECT 57.570 31.520 57.890 31.580 ;
        RECT 58.045 31.520 58.335 31.565 ;
        RECT 57.570 31.380 58.335 31.520 ;
        RECT 57.570 31.320 57.890 31.380 ;
        RECT 58.045 31.335 58.335 31.380 ;
        RECT 58.490 31.320 58.810 31.580 ;
        RECT 58.965 31.520 59.255 31.565 ;
        RECT 61.710 31.520 62.030 31.580 ;
        RECT 71.460 31.565 71.600 31.720 ;
        RECT 76.430 31.660 76.750 31.720 ;
        RECT 77.345 31.860 77.995 31.905 ;
        RECT 80.945 31.860 81.235 31.905 ;
        RECT 77.345 31.720 81.235 31.860 ;
        RECT 77.345 31.675 77.995 31.720 ;
        RECT 80.645 31.675 81.235 31.720 ;
        RECT 80.645 31.580 80.935 31.675 ;
        RECT 86.550 31.660 86.870 31.920 ;
        RECT 93.450 31.660 93.770 31.920 ;
        RECT 95.745 31.860 96.395 31.905 ;
        RECT 99.345 31.860 99.635 31.905 ;
        RECT 101.745 31.860 102.035 31.905 ;
        RECT 95.745 31.720 102.035 31.860 ;
        RECT 95.745 31.675 96.395 31.720 ;
        RECT 99.045 31.675 99.635 31.720 ;
        RECT 101.745 31.675 102.035 31.720 ;
        RECT 58.965 31.380 62.030 31.520 ;
        RECT 58.965 31.335 59.255 31.380 ;
        RECT 61.710 31.320 62.030 31.380 ;
        RECT 71.385 31.335 71.675 31.565 ;
        RECT 74.150 31.520 74.440 31.565 ;
        RECT 75.985 31.520 76.275 31.565 ;
        RECT 79.565 31.520 79.855 31.565 ;
        RECT 74.150 31.380 79.855 31.520 ;
        RECT 74.150 31.335 74.440 31.380 ;
        RECT 75.985 31.335 76.275 31.380 ;
        RECT 79.565 31.335 79.855 31.380 ;
        RECT 80.570 31.360 80.935 31.580 ;
        RECT 80.570 31.320 80.890 31.360 ;
        RECT 18.485 31.180 18.775 31.225 ;
        RECT 22.150 31.180 22.470 31.240 ;
        RECT 18.485 31.040 22.470 31.180 ;
        RECT 18.485 30.995 18.775 31.040 ;
        RECT 22.150 30.980 22.470 31.040 ;
        RECT 51.130 31.180 51.450 31.240 ;
        RECT 51.605 31.180 51.895 31.225 ;
        RECT 51.130 31.040 51.895 31.180 ;
        RECT 51.130 30.980 51.450 31.040 ;
        RECT 51.605 30.995 51.895 31.040 ;
        RECT 59.425 31.180 59.715 31.225 ;
        RECT 62.170 31.180 62.490 31.240 ;
        RECT 64.010 31.180 64.330 31.240 ;
        RECT 59.425 31.040 64.330 31.180 ;
        RECT 59.425 30.995 59.715 31.040 ;
        RECT 39.650 30.840 39.940 30.885 ;
        RECT 41.510 30.840 41.800 30.885 ;
        RECT 44.290 30.840 44.580 30.885 ;
        RECT 39.650 30.700 44.580 30.840 ;
        RECT 39.650 30.655 39.940 30.700 ;
        RECT 41.510 30.655 41.800 30.700 ;
        RECT 44.290 30.655 44.580 30.700 ;
        RECT 57.570 30.840 57.890 30.900 ;
        RECT 59.500 30.840 59.640 30.995 ;
        RECT 62.170 30.980 62.490 31.040 ;
        RECT 64.010 30.980 64.330 31.040 ;
        RECT 72.750 30.980 73.070 31.240 ;
        RECT 73.685 30.995 73.975 31.225 ;
        RECT 57.570 30.700 59.640 30.840 ;
        RECT 69.070 30.840 69.390 30.900 ;
        RECT 73.760 30.840 73.900 30.995 ;
        RECT 75.050 30.980 75.370 31.240 ;
        RECT 76.890 31.180 77.210 31.240 ;
        RECT 78.270 31.180 78.590 31.240 ;
        RECT 86.640 31.180 86.780 31.660 ;
        RECT 89.310 31.320 89.630 31.580 ;
        RECT 89.770 31.520 90.090 31.580 ;
        RECT 90.705 31.520 90.995 31.565 ;
        RECT 89.770 31.380 90.995 31.520 ;
        RECT 89.770 31.320 90.090 31.380 ;
        RECT 90.705 31.335 90.995 31.380 ;
        RECT 92.550 31.520 92.840 31.565 ;
        RECT 94.385 31.520 94.675 31.565 ;
        RECT 97.965 31.520 98.255 31.565 ;
        RECT 92.550 31.380 98.255 31.520 ;
        RECT 92.550 31.335 92.840 31.380 ;
        RECT 94.385 31.335 94.675 31.380 ;
        RECT 97.965 31.335 98.255 31.380 ;
        RECT 99.045 31.360 99.335 31.675 ;
        RECT 102.190 31.320 102.510 31.580 ;
        RECT 76.890 31.040 86.780 31.180 ;
        RECT 76.890 30.980 77.210 31.040 ;
        RECT 78.270 30.980 78.590 31.040 ;
        RECT 87.025 30.995 87.315 31.225 ;
        RECT 87.470 31.180 87.790 31.240 ;
        RECT 92.085 31.180 92.375 31.225 ;
        RECT 87.470 31.040 92.375 31.180 ;
        RECT 69.070 30.700 73.900 30.840 ;
        RECT 74.555 30.840 74.845 30.885 ;
        RECT 76.445 30.840 76.735 30.885 ;
        RECT 79.565 30.840 79.855 30.885 ;
        RECT 87.100 30.840 87.240 30.995 ;
        RECT 87.470 30.980 87.790 31.040 ;
        RECT 92.085 30.995 92.375 31.040 ;
        RECT 91.610 30.840 91.930 30.900 ;
        RECT 74.555 30.700 79.855 30.840 ;
        RECT 57.570 30.640 57.890 30.700 ;
        RECT 69.070 30.640 69.390 30.700 ;
        RECT 74.555 30.655 74.845 30.700 ;
        RECT 76.445 30.655 76.735 30.700 ;
        RECT 79.565 30.655 79.855 30.700 ;
        RECT 83.880 30.700 91.930 30.840 ;
        RECT 19.850 30.500 20.170 30.560 ;
        RECT 21.245 30.500 21.535 30.545 ;
        RECT 19.850 30.360 21.535 30.500 ;
        RECT 19.850 30.300 20.170 30.360 ;
        RECT 21.245 30.315 21.535 30.360 ;
        RECT 48.830 30.300 49.150 30.560 ;
        RECT 52.970 30.500 53.290 30.560 ;
        RECT 53.445 30.500 53.735 30.545 ;
        RECT 52.970 30.360 53.735 30.500 ;
        RECT 52.970 30.300 53.290 30.360 ;
        RECT 53.445 30.315 53.735 30.360 ;
        RECT 68.610 30.500 68.930 30.560 ;
        RECT 69.545 30.500 69.835 30.545 ;
        RECT 68.610 30.360 69.835 30.500 ;
        RECT 68.610 30.300 68.930 30.360 ;
        RECT 69.545 30.315 69.835 30.360 ;
        RECT 72.750 30.500 73.070 30.560 ;
        RECT 83.880 30.500 84.020 30.700 ;
        RECT 91.610 30.640 91.930 30.700 ;
        RECT 92.955 30.840 93.245 30.885 ;
        RECT 94.845 30.840 95.135 30.885 ;
        RECT 97.965 30.840 98.255 30.885 ;
        RECT 92.955 30.700 98.255 30.840 ;
        RECT 92.955 30.655 93.245 30.700 ;
        RECT 94.845 30.655 95.135 30.700 ;
        RECT 97.965 30.655 98.255 30.700 ;
        RECT 72.750 30.360 84.020 30.500 ;
        RECT 72.750 30.300 73.070 30.360 ;
        RECT 84.250 30.300 84.570 30.560 ;
        RECT 87.930 30.500 88.250 30.560 ;
        RECT 88.405 30.500 88.695 30.545 ;
        RECT 87.930 30.360 88.695 30.500 ;
        RECT 87.930 30.300 88.250 30.360 ;
        RECT 88.405 30.315 88.695 30.360 ;
        RECT 90.690 30.500 91.010 30.560 ;
        RECT 91.165 30.500 91.455 30.545 ;
        RECT 90.690 30.360 91.455 30.500 ;
        RECT 90.690 30.300 91.010 30.360 ;
        RECT 91.165 30.315 91.455 30.360 ;
        RECT 5.520 29.680 113.620 30.160 ;
        RECT 10.600 29.480 10.890 29.525 ;
        RECT 18.945 29.480 19.235 29.525 ;
        RECT 10.600 29.340 19.235 29.480 ;
        RECT 10.600 29.295 10.890 29.340 ;
        RECT 18.945 29.295 19.235 29.340 ;
        RECT 38.340 29.340 44.000 29.480 ;
        RECT 10.155 29.140 10.445 29.185 ;
        RECT 12.045 29.140 12.335 29.185 ;
        RECT 15.165 29.140 15.455 29.185 ;
        RECT 38.340 29.140 38.480 29.340 ;
        RECT 10.155 29.000 15.455 29.140 ;
        RECT 10.155 28.955 10.445 29.000 ;
        RECT 12.045 28.955 12.335 29.000 ;
        RECT 15.165 28.955 15.455 29.000 ;
        RECT 37.880 29.000 38.480 29.140 ;
        RECT 38.680 29.140 38.970 29.185 ;
        RECT 41.460 29.140 41.750 29.185 ;
        RECT 43.320 29.140 43.610 29.185 ;
        RECT 38.680 29.000 43.610 29.140 ;
        RECT 43.860 29.140 44.000 29.340 ;
        RECT 45.150 29.280 45.470 29.540 ;
        RECT 48.370 29.280 48.690 29.540 ;
        RECT 61.250 29.280 61.570 29.540 ;
        RECT 75.050 29.480 75.370 29.540 ;
        RECT 79.665 29.480 79.955 29.525 ;
        RECT 75.050 29.340 79.955 29.480 ;
        RECT 75.050 29.280 75.370 29.340 ;
        RECT 79.665 29.295 79.955 29.340 ;
        RECT 88.850 29.480 89.170 29.540 ;
        RECT 95.075 29.480 95.365 29.525 ;
        RECT 88.850 29.340 95.365 29.480 ;
        RECT 88.850 29.280 89.170 29.340 ;
        RECT 95.075 29.295 95.365 29.340 ;
        RECT 48.460 29.140 48.600 29.280 ;
        RECT 43.860 29.000 48.600 29.140 ;
        RECT 48.795 29.140 49.085 29.185 ;
        RECT 50.685 29.140 50.975 29.185 ;
        RECT 53.805 29.140 54.095 29.185 ;
        RECT 48.795 29.000 54.095 29.140 ;
        RECT 8.810 28.800 9.130 28.860 ;
        RECT 9.285 28.800 9.575 28.845 ;
        RECT 18.010 28.800 18.330 28.860 ;
        RECT 23.990 28.800 24.310 28.860 ;
        RECT 8.810 28.660 24.310 28.800 ;
        RECT 8.810 28.600 9.130 28.660 ;
        RECT 9.285 28.615 9.575 28.660 ;
        RECT 18.010 28.600 18.330 28.660 ;
        RECT 23.990 28.600 24.310 28.660 ;
        RECT 25.845 28.800 26.135 28.845 ;
        RECT 33.190 28.800 33.510 28.860 ;
        RECT 25.845 28.660 33.510 28.800 ;
        RECT 25.845 28.615 26.135 28.660 ;
        RECT 33.190 28.600 33.510 28.660 ;
        RECT 34.815 28.800 35.105 28.845 ;
        RECT 37.880 28.800 38.020 29.000 ;
        RECT 38.680 28.955 38.970 29.000 ;
        RECT 41.460 28.955 41.750 29.000 ;
        RECT 43.320 28.955 43.610 29.000 ;
        RECT 48.795 28.955 49.085 29.000 ;
        RECT 50.685 28.955 50.975 29.000 ;
        RECT 53.805 28.955 54.095 29.000 ;
        RECT 57.585 29.140 57.875 29.185 ;
        RECT 61.710 29.140 62.030 29.200 ;
        RECT 62.630 29.140 62.950 29.200 ;
        RECT 57.585 29.000 62.950 29.140 ;
        RECT 57.585 28.955 57.875 29.000 ;
        RECT 61.710 28.940 62.030 29.000 ;
        RECT 62.630 28.940 62.950 29.000 ;
        RECT 71.335 29.140 71.625 29.185 ;
        RECT 73.225 29.140 73.515 29.185 ;
        RECT 76.345 29.140 76.635 29.185 ;
        RECT 71.335 29.000 76.635 29.140 ;
        RECT 71.335 28.955 71.625 29.000 ;
        RECT 73.225 28.955 73.515 29.000 ;
        RECT 76.345 28.955 76.635 29.000 ;
        RECT 79.190 28.940 79.510 29.200 ;
        RECT 86.570 29.140 86.860 29.185 ;
        RECT 88.430 29.140 88.720 29.185 ;
        RECT 91.210 29.140 91.500 29.185 ;
        RECT 86.570 29.000 91.500 29.140 ;
        RECT 86.570 28.955 86.860 29.000 ;
        RECT 88.430 28.955 88.720 29.000 ;
        RECT 91.210 28.955 91.500 29.000 ;
        RECT 34.815 28.660 38.020 28.800 ;
        RECT 38.250 28.800 38.570 28.860 ;
        RECT 40.550 28.800 40.870 28.860 ;
        RECT 43.785 28.800 44.075 28.845 ;
        RECT 47.925 28.800 48.215 28.845 ;
        RECT 38.250 28.660 48.215 28.800 ;
        RECT 34.815 28.615 35.105 28.660 ;
        RECT 9.750 28.460 10.040 28.505 ;
        RECT 11.585 28.460 11.875 28.505 ;
        RECT 15.165 28.460 15.455 28.505 ;
        RECT 9.750 28.320 15.455 28.460 ;
        RECT 9.750 28.275 10.040 28.320 ;
        RECT 11.585 28.275 11.875 28.320 ;
        RECT 15.165 28.275 15.455 28.320 ;
        RECT 16.245 28.165 16.535 28.480 ;
        RECT 19.850 28.260 20.170 28.520 ;
        RECT 23.070 28.460 23.390 28.520 ;
        RECT 24.465 28.460 24.755 28.505 ;
        RECT 23.070 28.320 24.755 28.460 ;
        RECT 23.070 28.260 23.390 28.320 ;
        RECT 24.465 28.275 24.755 28.320 ;
        RECT 24.925 28.460 25.215 28.505 ;
        RECT 27.210 28.460 27.530 28.520 ;
        RECT 24.925 28.320 27.530 28.460 ;
        RECT 24.925 28.275 25.215 28.320 ;
        RECT 12.945 28.120 13.595 28.165 ;
        RECT 16.245 28.120 16.835 28.165 ;
        RECT 17.090 28.120 17.410 28.180 ;
        RECT 12.945 27.980 17.410 28.120 ;
        RECT 24.540 28.120 24.680 28.275 ;
        RECT 27.210 28.260 27.530 28.320 ;
        RECT 32.285 28.460 32.575 28.505 ;
        RECT 34.890 28.460 35.030 28.615 ;
        RECT 38.250 28.600 38.570 28.660 ;
        RECT 40.550 28.600 40.870 28.660 ;
        RECT 43.785 28.615 44.075 28.660 ;
        RECT 47.925 28.615 48.215 28.660 ;
        RECT 56.665 28.800 56.955 28.845 ;
        RECT 59.410 28.800 59.730 28.860 ;
        RECT 60.345 28.800 60.635 28.845 ;
        RECT 56.665 28.660 60.635 28.800 ;
        RECT 56.665 28.615 56.955 28.660 ;
        RECT 59.410 28.600 59.730 28.660 ;
        RECT 60.345 28.615 60.635 28.660 ;
        RECT 86.105 28.800 86.395 28.845 ;
        RECT 87.010 28.800 87.330 28.860 ;
        RECT 86.105 28.660 87.330 28.800 ;
        RECT 86.105 28.615 86.395 28.660 ;
        RECT 87.010 28.600 87.330 28.660 ;
        RECT 87.930 28.600 88.250 28.860 ;
        RECT 32.285 28.320 35.030 28.460 ;
        RECT 38.680 28.460 38.970 28.505 ;
        RECT 38.680 28.320 41.215 28.460 ;
        RECT 32.285 28.275 32.575 28.320 ;
        RECT 38.680 28.275 38.970 28.320 ;
        RECT 31.810 28.120 32.130 28.180 ;
        RECT 41.000 28.165 41.215 28.320 ;
        RECT 41.930 28.260 42.250 28.520 ;
        RECT 45.625 28.460 45.915 28.505 ;
        RECT 47.005 28.460 47.295 28.505 ;
        RECT 47.450 28.460 47.770 28.520 ;
        RECT 45.625 28.320 47.770 28.460 ;
        RECT 45.625 28.275 45.915 28.320 ;
        RECT 47.005 28.275 47.295 28.320 ;
        RECT 47.450 28.260 47.770 28.320 ;
        RECT 48.390 28.460 48.680 28.505 ;
        RECT 50.225 28.460 50.515 28.505 ;
        RECT 53.805 28.460 54.095 28.505 ;
        RECT 48.390 28.320 54.095 28.460 ;
        RECT 48.390 28.275 48.680 28.320 ;
        RECT 50.225 28.275 50.515 28.320 ;
        RECT 53.805 28.275 54.095 28.320 ;
        RECT 32.745 28.120 33.035 28.165 ;
        RECT 24.540 27.980 33.035 28.120 ;
        RECT 12.945 27.935 13.595 27.980 ;
        RECT 16.545 27.935 16.835 27.980 ;
        RECT 17.090 27.920 17.410 27.980 ;
        RECT 31.810 27.920 32.130 27.980 ;
        RECT 32.745 27.935 33.035 27.980 ;
        RECT 36.820 28.120 37.110 28.165 ;
        RECT 40.080 28.120 40.370 28.165 ;
        RECT 41.000 28.120 41.290 28.165 ;
        RECT 42.860 28.120 43.150 28.165 ;
        RECT 46.545 28.120 46.835 28.165 ;
        RECT 36.820 27.980 40.780 28.120 ;
        RECT 36.820 27.935 37.110 27.980 ;
        RECT 40.080 27.935 40.370 27.980 ;
        RECT 18.025 27.780 18.315 27.825 ;
        RECT 19.390 27.780 19.710 27.840 ;
        RECT 18.025 27.640 19.710 27.780 ;
        RECT 18.025 27.595 18.315 27.640 ;
        RECT 19.390 27.580 19.710 27.640 ;
        RECT 21.690 27.780 22.010 27.840 ;
        RECT 22.625 27.780 22.915 27.825 ;
        RECT 21.690 27.640 22.915 27.780 ;
        RECT 21.690 27.580 22.010 27.640 ;
        RECT 22.625 27.595 22.915 27.640 ;
        RECT 29.970 27.780 30.290 27.840 ;
        RECT 30.445 27.780 30.735 27.825 ;
        RECT 29.970 27.640 30.735 27.780 ;
        RECT 40.640 27.780 40.780 27.980 ;
        RECT 41.000 27.980 43.150 28.120 ;
        RECT 41.000 27.935 41.290 27.980 ;
        RECT 42.860 27.935 43.150 27.980 ;
        RECT 43.400 27.980 46.835 28.120 ;
        RECT 43.400 27.780 43.540 27.980 ;
        RECT 46.545 27.935 46.835 27.980 ;
        RECT 49.290 27.920 49.610 28.180 ;
        RECT 51.585 28.120 52.235 28.165 ;
        RECT 52.970 28.120 53.290 28.180 ;
        RECT 54.885 28.165 55.175 28.480 ;
        RECT 68.610 28.260 68.930 28.520 ;
        RECT 69.070 28.460 69.390 28.520 ;
        RECT 70.465 28.460 70.755 28.505 ;
        RECT 69.070 28.320 70.755 28.460 ;
        RECT 69.070 28.260 69.390 28.320 ;
        RECT 70.465 28.275 70.755 28.320 ;
        RECT 70.930 28.460 71.220 28.505 ;
        RECT 72.765 28.460 73.055 28.505 ;
        RECT 76.345 28.460 76.635 28.505 ;
        RECT 70.930 28.320 76.635 28.460 ;
        RECT 70.930 28.275 71.220 28.320 ;
        RECT 72.765 28.275 73.055 28.320 ;
        RECT 76.345 28.275 76.635 28.320 ;
        RECT 54.885 28.120 55.475 28.165 ;
        RECT 51.585 27.980 55.475 28.120 ;
        RECT 51.585 27.935 52.235 27.980 ;
        RECT 52.970 27.920 53.290 27.980 ;
        RECT 55.185 27.935 55.475 27.980 ;
        RECT 57.570 27.920 57.890 28.180 ;
        RECT 60.330 28.120 60.650 28.180 ;
        RECT 61.710 28.120 62.030 28.180 ;
        RECT 60.330 27.980 62.030 28.120 ;
        RECT 60.330 27.920 60.650 27.980 ;
        RECT 61.710 27.920 62.030 27.980 ;
        RECT 71.845 27.935 72.135 28.165 ;
        RECT 74.125 28.120 74.775 28.165 ;
        RECT 76.890 28.120 77.210 28.180 ;
        RECT 77.425 28.165 77.715 28.480 ;
        RECT 80.110 28.460 80.430 28.520 ;
        RECT 80.585 28.460 80.875 28.505 ;
        RECT 80.110 28.320 80.875 28.460 ;
        RECT 80.110 28.260 80.430 28.320 ;
        RECT 80.585 28.275 80.875 28.320 ;
        RECT 81.030 28.260 81.350 28.520 ;
        RECT 82.425 28.460 82.715 28.505 ;
        RECT 84.250 28.460 84.570 28.520 ;
        RECT 91.210 28.460 91.500 28.505 ;
        RECT 82.425 28.320 84.570 28.460 ;
        RECT 82.425 28.275 82.715 28.320 ;
        RECT 84.250 28.260 84.570 28.320 ;
        RECT 88.965 28.320 91.500 28.460 ;
        RECT 88.965 28.165 89.180 28.320 ;
        RECT 91.210 28.275 91.500 28.320 ;
        RECT 77.425 28.120 78.015 28.165 ;
        RECT 74.125 27.980 78.015 28.120 ;
        RECT 74.125 27.935 74.775 27.980 ;
        RECT 40.640 27.640 43.540 27.780 ;
        RECT 29.970 27.580 30.290 27.640 ;
        RECT 30.445 27.595 30.735 27.640 ;
        RECT 59.870 27.580 60.190 27.840 ;
        RECT 69.545 27.780 69.835 27.825 ;
        RECT 71.920 27.780 72.060 27.935 ;
        RECT 76.890 27.920 77.210 27.980 ;
        RECT 77.725 27.935 78.015 27.980 ;
        RECT 87.030 28.120 87.320 28.165 ;
        RECT 88.890 28.120 89.180 28.165 ;
        RECT 87.030 27.980 89.180 28.120 ;
        RECT 87.030 27.935 87.320 27.980 ;
        RECT 88.890 27.935 89.180 27.980 ;
        RECT 89.810 28.120 90.100 28.165 ;
        RECT 90.690 28.120 91.010 28.180 ;
        RECT 93.070 28.120 93.360 28.165 ;
        RECT 89.810 27.980 93.360 28.120 ;
        RECT 89.810 27.935 90.100 27.980 ;
        RECT 90.690 27.920 91.010 27.980 ;
        RECT 93.070 27.935 93.360 27.980 ;
        RECT 69.545 27.640 72.060 27.780 ;
        RECT 81.505 27.780 81.795 27.825 ;
        RECT 81.950 27.780 82.270 27.840 ;
        RECT 81.505 27.640 82.270 27.780 ;
        RECT 69.545 27.595 69.835 27.640 ;
        RECT 81.505 27.595 81.795 27.640 ;
        RECT 81.950 27.580 82.270 27.640 ;
        RECT 83.330 27.580 83.650 27.840 ;
        RECT 5.520 26.960 113.620 27.440 ;
        RECT 17.090 26.560 17.410 26.820 ;
        RECT 26.765 26.760 27.055 26.805 ;
        RECT 27.210 26.760 27.530 26.820 ;
        RECT 26.765 26.620 27.530 26.760 ;
        RECT 26.765 26.575 27.055 26.620 ;
        RECT 27.210 26.560 27.530 26.620 ;
        RECT 31.810 26.560 32.130 26.820 ;
        RECT 41.025 26.760 41.315 26.805 ;
        RECT 41.930 26.760 42.250 26.820 ;
        RECT 41.025 26.620 42.250 26.760 ;
        RECT 41.025 26.575 41.315 26.620 ;
        RECT 41.930 26.560 42.250 26.620 ;
        RECT 49.290 26.760 49.610 26.820 ;
        RECT 53.905 26.760 54.195 26.805 ;
        RECT 49.290 26.620 54.195 26.760 ;
        RECT 49.290 26.560 49.610 26.620 ;
        RECT 53.905 26.575 54.195 26.620 ;
        RECT 59.410 26.760 59.730 26.820 ;
        RECT 59.410 26.620 61.940 26.760 ;
        RECT 59.410 26.560 59.730 26.620 ;
        RECT 59.870 26.465 60.190 26.480 ;
        RECT 61.800 26.465 61.940 26.620 ;
        RECT 62.170 26.560 62.490 26.820 ;
        RECT 73.225 26.760 73.515 26.805 ;
        RECT 76.890 26.760 77.210 26.820 ;
        RECT 73.225 26.620 77.210 26.760 ;
        RECT 73.225 26.575 73.515 26.620 ;
        RECT 76.890 26.560 77.210 26.620 ;
        RECT 21.685 26.420 22.335 26.465 ;
        RECT 25.285 26.420 25.575 26.465 ;
        RECT 27.685 26.420 27.975 26.465 ;
        RECT 21.685 26.280 27.975 26.420 ;
        RECT 21.685 26.235 22.335 26.280 ;
        RECT 24.985 26.235 25.575 26.280 ;
        RECT 27.685 26.235 27.975 26.280 ;
        RECT 33.305 26.420 33.595 26.465 ;
        RECT 36.545 26.420 37.195 26.465 ;
        RECT 33.305 26.280 37.195 26.420 ;
        RECT 33.305 26.235 33.895 26.280 ;
        RECT 36.545 26.235 37.195 26.280 ;
        RECT 59.870 26.235 60.300 26.465 ;
        RECT 61.725 26.235 62.015 26.465 ;
        RECT 17.550 25.880 17.870 26.140 ;
        RECT 18.010 25.880 18.330 26.140 ;
        RECT 18.490 26.080 18.780 26.125 ;
        RECT 20.325 26.080 20.615 26.125 ;
        RECT 23.905 26.080 24.195 26.125 ;
        RECT 18.490 25.940 24.195 26.080 ;
        RECT 18.490 25.895 18.780 25.940 ;
        RECT 20.325 25.895 20.615 25.940 ;
        RECT 23.905 25.895 24.195 25.940 ;
        RECT 24.985 25.920 25.275 26.235 ;
        RECT 33.605 26.140 33.895 26.235 ;
        RECT 59.870 26.220 60.190 26.235 ;
        RECT 28.145 25.895 28.435 26.125 ;
        RECT 19.390 25.540 19.710 25.800 ;
        RECT 18.895 25.400 19.185 25.445 ;
        RECT 20.785 25.400 21.075 25.445 ;
        RECT 23.905 25.400 24.195 25.445 ;
        RECT 18.895 25.260 24.195 25.400 ;
        RECT 18.895 25.215 19.185 25.260 ;
        RECT 20.785 25.215 21.075 25.260 ;
        RECT 23.905 25.215 24.195 25.260 ;
        RECT 17.550 25.060 17.870 25.120 ;
        RECT 28.220 25.060 28.360 25.895 ;
        RECT 29.970 25.880 30.290 26.140 ;
        RECT 33.605 25.920 33.970 26.140 ;
        RECT 33.650 25.880 33.970 25.920 ;
        RECT 34.685 26.080 34.975 26.125 ;
        RECT 38.265 26.080 38.555 26.125 ;
        RECT 40.100 26.080 40.390 26.125 ;
        RECT 34.685 25.940 40.390 26.080 ;
        RECT 34.685 25.895 34.975 25.940 ;
        RECT 38.265 25.895 38.555 25.940 ;
        RECT 40.100 25.895 40.390 25.940 ;
        RECT 40.550 25.880 40.870 26.140 ;
        RECT 41.945 26.080 42.235 26.125 ;
        RECT 48.830 26.080 49.150 26.140 ;
        RECT 41.945 25.940 49.150 26.080 ;
        RECT 41.945 25.895 42.235 25.940 ;
        RECT 48.830 25.880 49.150 25.940 ;
        RECT 54.365 26.080 54.655 26.125 ;
        RECT 55.730 26.080 56.050 26.140 ;
        RECT 54.365 25.940 56.050 26.080 ;
        RECT 54.365 25.895 54.655 25.940 ;
        RECT 55.730 25.880 56.050 25.940 ;
        RECT 57.570 26.080 57.890 26.140 ;
        RECT 62.170 26.080 62.490 26.140 ;
        RECT 57.570 25.940 62.490 26.080 ;
        RECT 57.570 25.880 57.890 25.940 ;
        RECT 62.170 25.880 62.490 25.940 ;
        RECT 72.290 26.080 72.610 26.140 ;
        RECT 72.765 26.080 73.055 26.125 ;
        RECT 72.290 25.940 73.055 26.080 ;
        RECT 72.290 25.880 72.610 25.940 ;
        RECT 72.765 25.895 73.055 25.940 ;
        RECT 39.185 25.740 39.475 25.785 ;
        RECT 30.980 25.600 39.475 25.740 ;
        RECT 30.980 25.445 31.120 25.600 ;
        RECT 39.185 25.555 39.475 25.600 ;
        RECT 56.650 25.740 56.970 25.800 ;
        RECT 58.965 25.740 59.255 25.785 ;
        RECT 56.650 25.600 59.255 25.740 ;
        RECT 56.650 25.540 56.970 25.600 ;
        RECT 58.965 25.555 59.255 25.600 ;
        RECT 30.905 25.215 31.195 25.445 ;
        RECT 34.685 25.400 34.975 25.445 ;
        RECT 37.805 25.400 38.095 25.445 ;
        RECT 39.695 25.400 39.985 25.445 ;
        RECT 34.685 25.260 39.985 25.400 ;
        RECT 34.685 25.215 34.975 25.260 ;
        RECT 37.805 25.215 38.095 25.260 ;
        RECT 39.695 25.215 39.985 25.260 ;
        RECT 32.730 25.060 33.050 25.120 ;
        RECT 17.550 24.920 33.050 25.060 ;
        RECT 17.550 24.860 17.870 24.920 ;
        RECT 32.730 24.860 33.050 24.920 ;
        RECT 58.950 25.060 59.270 25.120 ;
        RECT 60.805 25.060 61.095 25.105 ;
        RECT 58.950 24.920 61.095 25.060 ;
        RECT 58.950 24.860 59.270 24.920 ;
        RECT 60.805 24.875 61.095 24.920 ;
        RECT 5.520 24.240 113.620 24.720 ;
        RECT 19.390 24.040 19.710 24.100 ;
        RECT 20.785 24.040 21.075 24.085 ;
        RECT 19.390 23.900 21.075 24.040 ;
        RECT 19.390 23.840 19.710 23.900 ;
        RECT 20.785 23.855 21.075 23.900 ;
        RECT 33.205 24.040 33.495 24.085 ;
        RECT 33.650 24.040 33.970 24.100 ;
        RECT 33.205 23.900 33.970 24.040 ;
        RECT 33.205 23.855 33.495 23.900 ;
        RECT 33.650 23.840 33.970 23.900 ;
        RECT 57.585 24.040 57.875 24.085 ;
        RECT 58.030 24.040 58.350 24.100 ;
        RECT 57.585 23.900 58.350 24.040 ;
        RECT 57.585 23.855 57.875 23.900 ;
        RECT 58.030 23.840 58.350 23.900 ;
        RECT 58.490 24.040 58.810 24.100 ;
        RECT 58.490 23.900 60.560 24.040 ;
        RECT 58.490 23.840 58.810 23.900 ;
        RECT 55.285 23.700 55.575 23.745 ;
        RECT 56.190 23.700 56.510 23.760 ;
        RECT 58.580 23.700 58.720 23.840 ;
        RECT 55.285 23.560 58.720 23.700 ;
        RECT 55.285 23.515 55.575 23.560 ;
        RECT 56.190 23.500 56.510 23.560 ;
        RECT 59.870 23.500 60.190 23.760 ;
        RECT 60.420 23.700 60.560 23.900 ;
        RECT 61.250 23.840 61.570 24.100 ;
        RECT 78.270 23.840 78.590 24.100 ;
        RECT 81.145 23.700 81.435 23.745 ;
        RECT 84.265 23.700 84.555 23.745 ;
        RECT 86.155 23.700 86.445 23.745 ;
        RECT 60.420 23.560 65.620 23.700 ;
        RECT 59.960 23.360 60.100 23.500 ;
        RECT 54.440 23.220 60.100 23.360 ;
        RECT 21.690 22.820 22.010 23.080 ;
        RECT 32.730 23.020 33.050 23.080 ;
        RECT 46.530 23.020 46.850 23.080 ;
        RECT 52.510 23.020 52.830 23.080 ;
        RECT 54.440 23.065 54.580 23.220 ;
        RECT 32.730 22.880 52.830 23.020 ;
        RECT 32.730 22.820 33.050 22.880 ;
        RECT 46.530 22.820 46.850 22.880 ;
        RECT 52.510 22.820 52.830 22.880 ;
        RECT 54.365 22.835 54.655 23.065 ;
        RECT 56.190 23.020 56.510 23.080 ;
        RECT 56.665 23.020 56.955 23.065 ;
        RECT 56.190 22.880 56.955 23.020 ;
        RECT 56.190 22.820 56.510 22.880 ;
        RECT 56.665 22.835 56.955 22.880 ;
        RECT 57.570 23.020 57.890 23.080 ;
        RECT 58.045 23.020 58.335 23.065 ;
        RECT 57.570 22.880 58.335 23.020 ;
        RECT 57.570 22.820 57.890 22.880 ;
        RECT 58.045 22.835 58.335 22.880 ;
        RECT 59.885 23.020 60.175 23.065 ;
        RECT 60.420 23.020 60.560 23.560 ;
        RECT 65.480 23.405 65.620 23.560 ;
        RECT 81.145 23.560 86.445 23.700 ;
        RECT 81.145 23.515 81.435 23.560 ;
        RECT 84.265 23.515 84.555 23.560 ;
        RECT 86.155 23.515 86.445 23.560 ;
        RECT 64.945 23.360 65.235 23.405 ;
        RECT 63.180 23.220 65.235 23.360 ;
        RECT 61.265 23.020 61.555 23.065 ;
        RECT 59.885 22.880 61.555 23.020 ;
        RECT 59.885 22.835 60.175 22.880 ;
        RECT 61.265 22.835 61.555 22.880 ;
        RECT 61.710 23.020 62.030 23.080 ;
        RECT 63.180 23.065 63.320 23.220 ;
        RECT 64.945 23.175 65.235 23.220 ;
        RECT 65.405 23.175 65.695 23.405 ;
        RECT 83.330 23.360 83.650 23.420 ;
        RECT 85.645 23.360 85.935 23.405 ;
        RECT 83.330 23.220 85.935 23.360 ;
        RECT 83.330 23.160 83.650 23.220 ;
        RECT 85.645 23.175 85.935 23.220 ;
        RECT 87.010 23.160 87.330 23.420 ;
        RECT 63.105 23.020 63.395 23.065 ;
        RECT 61.710 22.880 63.395 23.020 ;
        RECT 61.710 22.820 62.030 22.880 ;
        RECT 63.105 22.835 63.395 22.880 ;
        RECT 64.485 22.835 64.775 23.065 ;
        RECT 55.730 22.480 56.050 22.740 ;
        RECT 57.110 22.680 57.430 22.740 ;
        RECT 58.505 22.680 58.795 22.725 ;
        RECT 61.800 22.680 61.940 22.820 ;
        RECT 57.110 22.540 58.795 22.680 ;
        RECT 57.110 22.480 57.430 22.540 ;
        RECT 58.505 22.495 58.795 22.540 ;
        RECT 59.040 22.540 61.940 22.680 ;
        RECT 62.630 22.680 62.950 22.740 ;
        RECT 64.560 22.680 64.700 22.835 ;
        RECT 65.850 22.820 66.170 23.080 ;
        RECT 80.065 22.725 80.355 23.040 ;
        RECT 81.145 23.020 81.435 23.065 ;
        RECT 84.725 23.020 85.015 23.065 ;
        RECT 86.560 23.020 86.850 23.065 ;
        RECT 81.145 22.880 86.850 23.020 ;
        RECT 81.145 22.835 81.435 22.880 ;
        RECT 84.725 22.835 85.015 22.880 ;
        RECT 86.560 22.835 86.850 22.880 ;
        RECT 62.630 22.540 64.700 22.680 ;
        RECT 79.765 22.680 80.355 22.725 ;
        RECT 81.950 22.680 82.270 22.740 ;
        RECT 83.005 22.680 83.655 22.725 ;
        RECT 79.765 22.540 83.655 22.680 ;
        RECT 55.820 22.340 55.960 22.480 ;
        RECT 59.040 22.400 59.180 22.540 ;
        RECT 62.630 22.480 62.950 22.540 ;
        RECT 79.765 22.495 80.055 22.540 ;
        RECT 81.950 22.480 82.270 22.540 ;
        RECT 83.005 22.495 83.655 22.540 ;
        RECT 58.950 22.340 59.270 22.400 ;
        RECT 55.820 22.200 59.270 22.340 ;
        RECT 58.950 22.140 59.270 22.200 ;
        RECT 59.870 22.140 60.190 22.400 ;
        RECT 60.330 22.140 60.650 22.400 ;
        RECT 63.090 22.340 63.410 22.400 ;
        RECT 63.565 22.340 63.855 22.385 ;
        RECT 63.090 22.200 63.855 22.340 ;
        RECT 63.090 22.140 63.410 22.200 ;
        RECT 63.565 22.155 63.855 22.200 ;
        RECT 5.520 21.520 113.620 22.000 ;
        RECT 58.490 21.120 58.810 21.380 ;
        RECT 62.170 21.320 62.490 21.380 ;
        RECT 65.850 21.320 66.170 21.380 ;
        RECT 60.880 21.180 66.170 21.320 ;
        RECT 56.650 20.980 56.970 21.040 ;
        RECT 58.580 20.980 58.720 21.120 ;
        RECT 54.440 20.840 56.970 20.980 ;
        RECT 50.685 20.640 50.975 20.685 ;
        RECT 52.050 20.640 52.370 20.700 ;
        RECT 50.685 20.500 52.370 20.640 ;
        RECT 50.685 20.455 50.975 20.500 ;
        RECT 52.050 20.440 52.370 20.500 ;
        RECT 52.525 20.640 52.815 20.685 ;
        RECT 54.440 20.640 54.580 20.840 ;
        RECT 56.650 20.780 56.970 20.840 ;
        RECT 57.660 20.840 58.720 20.980 ;
        RECT 52.525 20.500 54.580 20.640 ;
        RECT 54.825 20.640 55.115 20.685 ;
        RECT 57.110 20.640 57.430 20.700 ;
        RECT 57.660 20.685 57.800 20.840 ;
        RECT 58.950 20.780 59.270 21.040 ;
        RECT 54.825 20.500 57.430 20.640 ;
        RECT 52.525 20.455 52.815 20.500 ;
        RECT 54.825 20.455 55.115 20.500 ;
        RECT 51.605 19.960 51.895 20.005 ;
        RECT 54.900 19.960 55.040 20.455 ;
        RECT 57.110 20.440 57.430 20.500 ;
        RECT 57.585 20.455 57.875 20.685 ;
        RECT 58.505 20.640 58.795 20.685 ;
        RECT 59.040 20.640 59.180 20.780 ;
        RECT 58.505 20.500 59.180 20.640 ;
        RECT 58.505 20.455 58.795 20.500 ;
        RECT 60.330 20.440 60.650 20.700 ;
        RECT 60.880 20.640 61.020 21.180 ;
        RECT 62.170 21.120 62.490 21.180 ;
        RECT 65.850 21.120 66.170 21.180 ;
        RECT 61.250 20.980 61.570 21.040 ;
        RECT 67.230 20.980 67.550 21.040 ;
        RECT 61.250 20.840 62.400 20.980 ;
        RECT 61.250 20.780 61.570 20.840 ;
        RECT 61.725 20.640 62.015 20.685 ;
        RECT 60.880 20.500 62.015 20.640 ;
        RECT 62.260 20.640 62.400 20.840 ;
        RECT 65.480 20.840 67.550 20.980 ;
        RECT 63.105 20.640 63.395 20.685 ;
        RECT 65.480 20.640 65.620 20.840 ;
        RECT 67.230 20.780 67.550 20.840 ;
        RECT 69.065 20.980 69.715 21.025 ;
        RECT 72.665 20.980 72.955 21.025 ;
        RECT 69.065 20.840 72.955 20.980 ;
        RECT 69.065 20.795 69.715 20.840 ;
        RECT 72.365 20.795 72.955 20.840 ;
        RECT 72.365 20.700 72.655 20.795 ;
        RECT 62.260 20.500 65.620 20.640 ;
        RECT 65.870 20.640 66.160 20.685 ;
        RECT 67.705 20.640 67.995 20.685 ;
        RECT 71.285 20.640 71.575 20.685 ;
        RECT 65.870 20.500 71.575 20.640 ;
        RECT 61.725 20.455 62.015 20.500 ;
        RECT 63.105 20.455 63.395 20.500 ;
        RECT 65.870 20.455 66.160 20.500 ;
        RECT 67.705 20.455 67.995 20.500 ;
        RECT 71.285 20.455 71.575 20.500 ;
        RECT 72.290 20.480 72.655 20.700 ;
        RECT 72.290 20.440 72.610 20.480 ;
        RECT 55.285 20.300 55.575 20.345 ;
        RECT 58.045 20.300 58.335 20.345 ;
        RECT 58.950 20.300 59.270 20.360 ;
        RECT 55.285 20.160 59.270 20.300 ;
        RECT 55.285 20.115 55.575 20.160 ;
        RECT 58.045 20.115 58.335 20.160 ;
        RECT 58.950 20.100 59.270 20.160 ;
        RECT 59.870 20.300 60.190 20.360 ;
        RECT 62.645 20.300 62.935 20.345 ;
        RECT 59.870 20.160 62.935 20.300 ;
        RECT 59.870 20.100 60.190 20.160 ;
        RECT 62.645 20.115 62.935 20.160 ;
        RECT 64.470 20.300 64.790 20.360 ;
        RECT 65.405 20.300 65.695 20.345 ;
        RECT 66.785 20.300 67.075 20.345 ;
        RECT 64.470 20.160 65.695 20.300 ;
        RECT 64.470 20.100 64.790 20.160 ;
        RECT 65.405 20.115 65.695 20.160 ;
        RECT 65.940 20.160 67.075 20.300 ;
        RECT 62.170 19.960 62.490 20.020 ;
        RECT 51.605 19.820 62.490 19.960 ;
        RECT 51.605 19.775 51.895 19.820 ;
        RECT 49.290 19.620 49.610 19.680 ;
        RECT 49.765 19.620 50.055 19.665 ;
        RECT 49.290 19.480 50.055 19.620 ;
        RECT 49.290 19.420 49.610 19.480 ;
        RECT 49.765 19.435 50.055 19.480 ;
        RECT 53.430 19.420 53.750 19.680 ;
        RECT 58.490 19.620 58.810 19.680 ;
        RECT 59.960 19.665 60.100 19.820 ;
        RECT 62.170 19.760 62.490 19.820 ;
        RECT 64.945 19.960 65.235 20.005 ;
        RECT 65.940 19.960 66.080 20.160 ;
        RECT 66.785 20.115 67.075 20.160 ;
        RECT 67.230 20.300 67.550 20.360 ;
        RECT 74.145 20.300 74.435 20.345 ;
        RECT 67.230 20.160 74.435 20.300 ;
        RECT 67.230 20.100 67.550 20.160 ;
        RECT 74.145 20.115 74.435 20.160 ;
        RECT 64.945 19.820 66.080 19.960 ;
        RECT 66.275 19.960 66.565 20.005 ;
        RECT 68.165 19.960 68.455 20.005 ;
        RECT 71.285 19.960 71.575 20.005 ;
        RECT 66.275 19.820 71.575 19.960 ;
        RECT 64.945 19.775 65.235 19.820 ;
        RECT 66.275 19.775 66.565 19.820 ;
        RECT 68.165 19.775 68.455 19.820 ;
        RECT 71.285 19.775 71.575 19.820 ;
        RECT 58.965 19.620 59.255 19.665 ;
        RECT 58.490 19.480 59.255 19.620 ;
        RECT 58.490 19.420 58.810 19.480 ;
        RECT 58.965 19.435 59.255 19.480 ;
        RECT 59.885 19.435 60.175 19.665 ;
        RECT 64.470 19.620 64.790 19.680 ;
        RECT 69.070 19.620 69.390 19.680 ;
        RECT 64.470 19.480 69.390 19.620 ;
        RECT 64.470 19.420 64.790 19.480 ;
        RECT 69.070 19.420 69.390 19.480 ;
        RECT 5.520 18.800 113.620 19.280 ;
        RECT 52.050 18.600 52.370 18.660 ;
        RECT 57.125 18.600 57.415 18.645 ;
        RECT 52.050 18.460 57.415 18.600 ;
        RECT 52.050 18.400 52.370 18.460 ;
        RECT 57.125 18.415 57.415 18.460 ;
        RECT 58.030 18.400 58.350 18.660 ;
        RECT 59.410 18.400 59.730 18.660 ;
        RECT 72.290 18.400 72.610 18.660 ;
        RECT 48.795 18.260 49.085 18.305 ;
        RECT 50.685 18.260 50.975 18.305 ;
        RECT 53.805 18.260 54.095 18.305 ;
        RECT 48.795 18.120 54.095 18.260 ;
        RECT 48.795 18.075 49.085 18.120 ;
        RECT 50.685 18.075 50.975 18.120 ;
        RECT 53.805 18.075 54.095 18.120 ;
        RECT 56.665 18.260 56.955 18.305 ;
        RECT 59.500 18.260 59.640 18.400 ;
        RECT 56.665 18.120 59.640 18.260 ;
        RECT 60.295 18.260 60.585 18.305 ;
        RECT 62.185 18.260 62.475 18.305 ;
        RECT 65.305 18.260 65.595 18.305 ;
        RECT 60.295 18.120 65.595 18.260 ;
        RECT 56.665 18.075 56.955 18.120 ;
        RECT 60.295 18.075 60.585 18.120 ;
        RECT 62.185 18.075 62.475 18.120 ;
        RECT 65.305 18.075 65.595 18.120 ;
        RECT 38.250 17.920 38.570 17.980 ;
        RECT 46.070 17.920 46.390 17.980 ;
        RECT 47.925 17.920 48.215 17.965 ;
        RECT 38.250 17.780 48.215 17.920 ;
        RECT 38.250 17.720 38.570 17.780 ;
        RECT 46.070 17.720 46.390 17.780 ;
        RECT 47.925 17.735 48.215 17.780 ;
        RECT 49.290 17.720 49.610 17.980 ;
        RECT 59.425 17.920 59.715 17.965 ;
        RECT 64.470 17.920 64.790 17.980 ;
        RECT 59.425 17.780 64.790 17.920 ;
        RECT 59.425 17.735 59.715 17.780 ;
        RECT 64.470 17.720 64.790 17.780 ;
        RECT 65.850 17.920 66.170 17.980 ;
        RECT 69.545 17.920 69.835 17.965 ;
        RECT 65.850 17.780 69.835 17.920 ;
        RECT 65.850 17.720 66.170 17.780 ;
        RECT 69.545 17.735 69.835 17.780 ;
        RECT 46.530 17.380 46.850 17.640 ;
        RECT 48.390 17.580 48.680 17.625 ;
        RECT 50.225 17.580 50.515 17.625 ;
        RECT 53.805 17.580 54.095 17.625 ;
        RECT 48.390 17.440 54.095 17.580 ;
        RECT 48.390 17.395 48.680 17.440 ;
        RECT 50.225 17.395 50.515 17.440 ;
        RECT 53.805 17.395 54.095 17.440 ;
        RECT 51.585 17.240 52.235 17.285 ;
        RECT 52.510 17.240 52.830 17.300 ;
        RECT 54.885 17.285 55.175 17.600 ;
        RECT 59.890 17.580 60.180 17.625 ;
        RECT 61.725 17.580 62.015 17.625 ;
        RECT 65.305 17.580 65.595 17.625 ;
        RECT 59.890 17.440 65.595 17.580 ;
        RECT 59.890 17.395 60.180 17.440 ;
        RECT 61.725 17.395 62.015 17.440 ;
        RECT 65.305 17.395 65.595 17.440 ;
        RECT 66.385 17.580 66.675 17.600 ;
        RECT 70.925 17.580 71.215 17.625 ;
        RECT 66.385 17.440 71.215 17.580 ;
        RECT 54.885 17.240 55.475 17.285 ;
        RECT 51.585 17.100 55.475 17.240 ;
        RECT 51.585 17.055 52.235 17.100 ;
        RECT 52.510 17.040 52.830 17.100 ;
        RECT 55.185 17.055 55.475 17.100 ;
        RECT 57.965 17.240 58.255 17.285 ;
        RECT 58.490 17.240 58.810 17.300 ;
        RECT 57.965 17.100 58.810 17.240 ;
        RECT 57.965 17.055 58.255 17.100 ;
        RECT 58.490 17.040 58.810 17.100 ;
        RECT 58.950 17.040 59.270 17.300 ;
        RECT 60.790 17.040 61.110 17.300 ;
        RECT 66.385 17.285 66.675 17.440 ;
        RECT 70.925 17.395 71.215 17.440 ;
        RECT 71.385 17.580 71.675 17.625 ;
        RECT 71.830 17.580 72.150 17.640 ;
        RECT 71.385 17.440 72.150 17.580 ;
        RECT 71.385 17.395 71.675 17.440 ;
        RECT 71.830 17.380 72.150 17.440 ;
        RECT 63.085 17.240 63.735 17.285 ;
        RECT 66.385 17.240 66.975 17.285 ;
        RECT 63.085 17.100 66.975 17.240 ;
        RECT 63.085 17.055 63.735 17.100 ;
        RECT 66.685 17.055 66.975 17.100 ;
        RECT 46.990 16.700 47.310 16.960 ;
        RECT 5.520 16.080 113.620 16.560 ;
        RECT 52.510 15.880 52.830 15.940 ;
        RECT 55.745 15.880 56.035 15.925 ;
        RECT 52.510 15.740 56.035 15.880 ;
        RECT 52.510 15.680 52.830 15.740 ;
        RECT 55.745 15.695 56.035 15.740 ;
        RECT 60.790 15.880 61.110 15.940 ;
        RECT 62.645 15.880 62.935 15.925 ;
        RECT 60.790 15.740 62.935 15.880 ;
        RECT 60.790 15.680 61.110 15.740 ;
        RECT 62.645 15.695 62.935 15.740 ;
        RECT 46.990 15.540 47.310 15.600 ;
        RECT 49.745 15.540 50.395 15.585 ;
        RECT 53.345 15.540 53.635 15.585 ;
        RECT 46.990 15.400 53.635 15.540 ;
        RECT 46.990 15.340 47.310 15.400 ;
        RECT 49.745 15.355 50.395 15.400 ;
        RECT 53.045 15.355 53.635 15.400 ;
        RECT 58.490 15.540 58.810 15.600 ;
        RECT 60.345 15.540 60.635 15.585 ;
        RECT 58.490 15.400 60.635 15.540 ;
        RECT 46.070 15.000 46.390 15.260 ;
        RECT 46.550 15.200 46.840 15.245 ;
        RECT 48.385 15.200 48.675 15.245 ;
        RECT 51.965 15.200 52.255 15.245 ;
        RECT 46.550 15.060 52.255 15.200 ;
        RECT 46.550 15.015 46.840 15.060 ;
        RECT 48.385 15.015 48.675 15.060 ;
        RECT 51.965 15.015 52.255 15.060 ;
        RECT 53.045 15.040 53.335 15.355 ;
        RECT 58.490 15.340 58.810 15.400 ;
        RECT 60.345 15.355 60.635 15.400 ;
        RECT 61.425 15.540 61.715 15.585 ;
        RECT 63.090 15.540 63.410 15.600 ;
        RECT 61.425 15.400 63.410 15.540 ;
        RECT 61.425 15.355 61.715 15.400 ;
        RECT 63.090 15.340 63.410 15.400 ;
        RECT 56.205 15.200 56.495 15.245 ;
        RECT 63.565 15.200 63.855 15.245 ;
        RECT 53.980 15.060 56.495 15.200 ;
        RECT 47.465 14.860 47.755 14.905 ;
        RECT 53.430 14.860 53.750 14.920 ;
        RECT 47.465 14.720 53.750 14.860 ;
        RECT 47.465 14.675 47.755 14.720 ;
        RECT 53.430 14.660 53.750 14.720 ;
        RECT 46.955 14.520 47.245 14.565 ;
        RECT 48.845 14.520 49.135 14.565 ;
        RECT 51.965 14.520 52.255 14.565 ;
        RECT 46.955 14.380 52.255 14.520 ;
        RECT 46.955 14.335 47.245 14.380 ;
        RECT 48.845 14.335 49.135 14.380 ;
        RECT 51.965 14.335 52.255 14.380 ;
        RECT 46.530 14.180 46.850 14.240 ;
        RECT 53.980 14.180 54.120 15.060 ;
        RECT 56.205 15.015 56.495 15.060 ;
        RECT 62.260 15.060 63.855 15.200 ;
        RECT 54.825 14.860 55.115 14.905 ;
        RECT 56.650 14.860 56.970 14.920 ;
        RECT 54.825 14.720 56.970 14.860 ;
        RECT 54.825 14.675 55.115 14.720 ;
        RECT 56.650 14.660 56.970 14.720 ;
        RECT 62.260 14.565 62.400 15.060 ;
        RECT 63.565 15.015 63.855 15.060 ;
        RECT 62.185 14.335 62.475 14.565 ;
        RECT 46.530 14.040 54.120 14.180 ;
        RECT 59.870 14.180 60.190 14.240 ;
        RECT 61.265 14.180 61.555 14.225 ;
        RECT 59.870 14.040 61.555 14.180 ;
        RECT 46.530 13.980 46.850 14.040 ;
        RECT 59.870 13.980 60.190 14.040 ;
        RECT 61.265 13.995 61.555 14.040 ;
        RECT 5.520 13.360 113.620 13.840 ;
        RECT 5.520 10.640 113.620 11.120 ;
      LAYER met2 ;
        RECT 39.010 128.790 39.400 128.930 ;
        RECT 104.790 128.790 106.100 128.930 ;
        RECT 1.940 115.270 2.200 115.590 ;
        RECT 2.000 113.405 2.140 115.270 ;
        RECT 1.930 113.035 2.210 113.405 ;
        RECT 2.920 110.490 3.060 128.280 ;
        RECT 2.860 110.170 3.120 110.490 ;
        RECT 8.900 108.450 9.040 128.280 ;
        RECT 9.580 116.775 11.460 117.145 ;
        RECT 14.880 113.970 15.020 128.280 ;
        RECT 14.420 113.890 15.020 113.970 ;
        RECT 14.360 113.830 15.020 113.890 ;
        RECT 14.360 113.570 14.620 113.830 ;
        RECT 18.040 113.230 18.300 113.550 ;
        RECT 20.860 113.290 21.000 128.280 ;
        RECT 24.580 114.055 26.460 114.425 ;
        RECT 26.840 113.890 26.980 128.280 ;
        RECT 32.820 116.610 32.960 128.280 ;
        RECT 32.760 116.290 33.020 116.610 ;
        RECT 35.520 115.610 35.780 115.930 ;
        RECT 33.680 115.270 33.940 115.590 ;
        RECT 26.780 113.570 27.040 113.890 ;
        RECT 17.580 112.550 17.840 112.870 ;
        RECT 9.580 111.335 11.460 111.705 ;
        RECT 13.440 110.170 13.700 110.490 ;
        RECT 8.840 108.130 9.100 108.450 ;
        RECT 7.000 107.110 7.260 107.430 ;
        RECT 8.380 107.110 8.640 107.430 ;
        RECT 7.060 99.610 7.200 107.110 ;
        RECT 8.440 105.730 8.580 107.110 ;
        RECT 9.580 105.895 11.460 106.265 ;
        RECT 8.380 105.410 8.640 105.730 ;
        RECT 13.500 101.990 13.640 110.170 ;
        RECT 14.360 109.490 14.620 109.810 ;
        RECT 15.740 109.490 16.000 109.810 ;
        RECT 14.420 105.390 14.560 109.490 ;
        RECT 15.280 107.450 15.540 107.770 ;
        RECT 14.360 105.070 14.620 105.390 ;
        RECT 15.340 104.710 15.480 107.450 ;
        RECT 15.800 105.730 15.940 109.490 ;
        RECT 17.640 107.090 17.780 112.550 ;
        RECT 18.100 108.450 18.240 113.230 ;
        RECT 20.860 113.150 21.460 113.290 ;
        RECT 29.540 113.230 29.800 113.550 ;
        RECT 20.800 112.550 21.060 112.870 ;
        RECT 20.860 110.490 21.000 112.550 ;
        RECT 20.800 110.170 21.060 110.490 ;
        RECT 20.800 109.380 21.060 109.470 ;
        RECT 21.320 109.380 21.460 113.150 ;
        RECT 22.640 112.550 22.900 112.870 ;
        RECT 20.800 109.240 21.460 109.380 ;
        RECT 20.800 109.150 21.060 109.240 ;
        RECT 22.700 108.450 22.840 112.550 ;
        RECT 29.600 110.490 29.740 113.230 ;
        RECT 33.740 110.490 33.880 115.270 ;
        RECT 29.540 110.170 29.800 110.490 ;
        RECT 33.680 110.170 33.940 110.490 ;
        RECT 32.760 109.830 33.020 110.150 ;
        RECT 33.220 109.830 33.480 110.150 ;
        RECT 26.780 109.490 27.040 109.810 ;
        RECT 27.240 109.490 27.500 109.810 ;
        RECT 24.580 108.615 26.460 108.985 ;
        RECT 26.840 108.450 26.980 109.490 ;
        RECT 18.040 108.130 18.300 108.450 ;
        RECT 22.640 108.130 22.900 108.450 ;
        RECT 26.780 108.130 27.040 108.450 ;
        RECT 23.560 107.450 23.820 107.770 ;
        RECT 21.720 107.110 21.980 107.430 ;
        RECT 17.580 106.770 17.840 107.090 ;
        RECT 15.740 105.410 16.000 105.730 ;
        RECT 15.280 104.390 15.540 104.710 ;
        RECT 18.040 104.050 18.300 104.370 ;
        RECT 13.440 101.670 13.700 101.990 ;
        RECT 17.580 101.670 17.840 101.990 ;
        RECT 9.580 100.455 11.460 100.825 ;
        RECT 13.500 99.610 13.640 101.670 ;
        RECT 7.000 99.290 7.260 99.610 ;
        RECT 13.440 99.290 13.700 99.610 ;
        RECT 14.820 99.290 15.080 99.610 ;
        RECT 9.760 98.950 10.020 99.270 ;
        RECT 9.820 97.570 9.960 98.950 ;
        RECT 12.520 98.610 12.780 98.930 ;
        RECT 12.580 97.570 12.720 98.610 ;
        RECT 9.760 97.250 10.020 97.570 ;
        RECT 12.520 97.250 12.780 97.570 ;
        RECT 13.500 96.550 13.640 99.290 ;
        RECT 14.360 96.910 14.620 97.230 ;
        RECT 13.440 96.230 13.700 96.550 ;
        RECT 9.580 95.015 11.460 95.385 ;
        RECT 9.760 92.830 10.020 93.150 ;
        RECT 12.520 92.830 12.780 93.150 ;
        RECT 9.820 91.450 9.960 92.830 ;
        RECT 12.580 91.790 12.720 92.830 ;
        RECT 12.520 91.470 12.780 91.790 ;
        RECT 9.760 91.130 10.020 91.450 ;
        RECT 8.840 90.790 9.100 91.110 ;
        RECT 8.900 88.730 9.040 90.790 ;
        RECT 9.580 89.575 11.460 89.945 ;
        RECT 13.500 88.730 13.640 96.230 ;
        RECT 14.420 94.850 14.560 96.910 ;
        RECT 14.880 96.890 15.020 99.290 ;
        RECT 16.660 98.950 16.920 99.270 ;
        RECT 14.820 96.570 15.080 96.890 ;
        RECT 14.360 94.530 14.620 94.850 ;
        RECT 14.880 93.830 15.020 96.570 ;
        RECT 16.720 93.830 16.860 98.950 ;
        RECT 17.640 97.570 17.780 101.670 ;
        RECT 17.580 97.250 17.840 97.570 ;
        RECT 14.820 93.510 15.080 93.830 ;
        RECT 16.660 93.510 16.920 93.830 ;
        RECT 8.840 88.410 9.100 88.730 ;
        RECT 13.440 88.410 13.700 88.730 ;
        RECT 7.920 79.230 8.180 79.550 ;
        RECT 7.980 74.790 8.120 79.230 ;
        RECT 8.900 77.850 9.040 88.410 ;
        RECT 10.680 88.070 10.940 88.390 ;
        RECT 10.740 86.350 10.880 88.070 ;
        RECT 14.360 87.730 14.620 88.050 ;
        RECT 14.420 86.350 14.560 87.730 ;
        RECT 10.680 86.030 10.940 86.350 ;
        RECT 14.360 86.030 14.620 86.350 ;
        RECT 14.880 86.010 15.020 93.510 ;
        RECT 16.720 88.050 16.860 93.510 ;
        RECT 17.580 90.110 17.840 90.430 ;
        RECT 16.660 87.730 16.920 88.050 ;
        RECT 17.640 86.010 17.780 90.110 ;
        RECT 14.820 85.690 15.080 86.010 ;
        RECT 17.580 85.690 17.840 86.010 ;
        RECT 9.580 84.135 11.460 84.505 ;
        RECT 14.880 83.970 15.020 85.690 ;
        RECT 14.820 83.650 15.080 83.970 ;
        RECT 11.600 79.230 11.860 79.550 ;
        RECT 9.580 78.695 11.460 79.065 ;
        RECT 11.660 77.850 11.800 79.230 ;
        RECT 8.840 77.530 9.100 77.850 ;
        RECT 11.600 77.530 11.860 77.850 ;
        RECT 13.440 77.530 13.700 77.850 ;
        RECT 8.380 75.040 8.640 75.130 ;
        RECT 8.900 75.040 9.040 77.530 ;
        RECT 12.520 75.150 12.780 75.470 ;
        RECT 8.380 74.900 9.040 75.040 ;
        RECT 8.380 74.810 8.640 74.900 ;
        RECT 7.920 74.470 8.180 74.790 ;
        RECT 9.580 73.255 11.460 73.625 ;
        RECT 12.580 73.090 12.720 75.150 ;
        RECT 12.520 72.770 12.780 73.090 ;
        RECT 13.500 72.070 13.640 77.530 ;
        RECT 13.440 71.750 13.700 72.070 ;
        RECT 11.600 68.350 11.860 68.670 ;
        RECT 9.580 67.815 11.460 68.185 ;
        RECT 11.660 66.630 11.800 68.350 ;
        RECT 13.500 66.630 13.640 71.750 ;
        RECT 11.600 66.310 11.860 66.630 ;
        RECT 13.440 66.310 13.700 66.630 ;
        RECT 8.840 65.630 9.100 65.950 ;
        RECT 11.600 65.630 11.860 65.950 ;
        RECT 12.980 65.630 13.240 65.950 ;
        RECT 8.900 64.250 9.040 65.630 ;
        RECT 8.840 63.930 9.100 64.250 ;
        RECT 7.920 63.590 8.180 63.910 ;
        RECT 7.980 61.190 8.120 63.590 ;
        RECT 9.580 62.375 11.460 62.745 ;
        RECT 11.660 61.530 11.800 65.630 ;
        RECT 13.040 64.590 13.180 65.630 ;
        RECT 12.980 64.270 13.240 64.590 ;
        RECT 13.500 64.250 13.640 66.310 ;
        RECT 13.440 63.930 13.700 64.250 ;
        RECT 11.600 61.210 11.860 61.530 ;
        RECT 7.920 60.870 8.180 61.190 ;
        RECT 7.980 53.030 8.120 60.870 ;
        RECT 9.580 56.935 11.460 57.305 ;
        RECT 13.500 56.090 13.640 63.930 ;
        RECT 14.880 62.170 15.020 83.650 ;
        RECT 16.660 80.590 16.920 80.910 ;
        RECT 16.720 75.810 16.860 80.590 ;
        RECT 16.660 75.490 16.920 75.810 ;
        RECT 15.280 74.810 15.540 75.130 ;
        RECT 15.340 69.350 15.480 74.810 ;
        RECT 16.660 70.050 16.920 70.370 ;
        RECT 15.280 69.030 15.540 69.350 ;
        RECT 15.340 64.930 15.480 69.030 ;
        RECT 16.720 66.970 16.860 70.050 ;
        RECT 17.580 69.710 17.840 70.030 ;
        RECT 17.640 66.970 17.780 69.710 ;
        RECT 18.100 69.350 18.240 104.050 ;
        RECT 18.500 98.270 18.760 98.590 ;
        RECT 18.560 96.890 18.700 98.270 ;
        RECT 18.500 96.570 18.760 96.890 ;
        RECT 20.330 96.715 20.610 97.085 ;
        RECT 20.340 96.570 20.600 96.715 ;
        RECT 18.960 93.170 19.220 93.490 ;
        RECT 19.020 89.410 19.160 93.170 ;
        RECT 20.800 92.830 21.060 93.150 ;
        RECT 19.420 91.130 19.680 91.450 ;
        RECT 18.960 89.090 19.220 89.410 ;
        RECT 19.480 89.070 19.620 91.130 ;
        RECT 20.860 90.770 21.000 92.830 ;
        RECT 20.800 90.450 21.060 90.770 ;
        RECT 19.420 88.750 19.680 89.070 ;
        RECT 19.480 86.350 19.620 88.750 ;
        RECT 20.860 88.390 21.000 90.450 ;
        RECT 20.800 88.070 21.060 88.390 ;
        RECT 19.420 86.030 19.680 86.350 ;
        RECT 20.860 85.670 21.000 88.070 ;
        RECT 21.260 86.370 21.520 86.690 ;
        RECT 21.320 86.010 21.460 86.370 ;
        RECT 21.260 85.690 21.520 86.010 ;
        RECT 20.800 85.350 21.060 85.670 ;
        RECT 21.260 84.670 21.520 84.990 ;
        RECT 18.960 80.250 19.220 80.570 ;
        RECT 19.020 75.810 19.160 80.250 ;
        RECT 19.880 79.910 20.140 80.230 ;
        RECT 19.940 79.550 20.080 79.910 ;
        RECT 19.880 79.230 20.140 79.550 ;
        RECT 18.960 75.490 19.220 75.810 ;
        RECT 19.940 74.790 20.080 79.230 ;
        RECT 19.880 74.470 20.140 74.790 ;
        RECT 19.940 70.030 20.080 74.470 ;
        RECT 19.880 69.710 20.140 70.030 ;
        RECT 18.040 69.030 18.300 69.350 ;
        RECT 19.880 69.030 20.140 69.350 ;
        RECT 20.800 69.030 21.060 69.350 ;
        RECT 16.660 66.650 16.920 66.970 ;
        RECT 17.580 66.650 17.840 66.970 ;
        RECT 15.280 64.610 15.540 64.930 ;
        RECT 16.720 62.210 16.860 66.650 ;
        RECT 17.120 62.910 17.380 63.230 ;
        RECT 14.880 62.030 15.480 62.170 ;
        RECT 15.340 59.150 15.480 62.030 ;
        RECT 16.660 61.890 16.920 62.210 ;
        RECT 17.180 60.850 17.320 62.910 ;
        RECT 17.120 60.530 17.380 60.850 ;
        RECT 17.580 60.530 17.840 60.850 ;
        RECT 15.280 58.830 15.540 59.150 ;
        RECT 16.200 58.490 16.460 58.810 ;
        RECT 13.440 55.770 13.700 56.090 ;
        RECT 16.260 55.750 16.400 58.490 ;
        RECT 12.980 55.430 13.240 55.750 ;
        RECT 16.200 55.430 16.460 55.750 ;
        RECT 11.140 54.750 11.400 55.070 ;
        RECT 11.200 53.710 11.340 54.750 ;
        RECT 11.140 53.390 11.400 53.710 ;
        RECT 7.920 52.710 8.180 53.030 ;
        RECT 9.580 51.495 11.460 51.865 ;
        RECT 13.040 50.990 13.180 55.430 ;
        RECT 13.900 55.090 14.160 55.410 ;
        RECT 13.960 51.330 14.100 55.090 ;
        RECT 17.120 53.390 17.380 53.710 ;
        RECT 13.900 51.010 14.160 51.330 ;
        RECT 12.980 50.670 13.240 50.990 ;
        RECT 8.380 49.650 8.640 49.970 ;
        RECT 11.140 49.650 11.400 49.970 ;
        RECT 8.440 48.125 8.580 49.650 ;
        RECT 11.200 48.610 11.340 49.650 ;
        RECT 11.140 48.290 11.400 48.610 ;
        RECT 8.370 47.755 8.650 48.125 ;
        RECT 15.740 47.270 16.000 47.590 ;
        RECT 9.580 46.055 11.460 46.425 ;
        RECT 15.800 45.550 15.940 47.270 ;
        RECT 15.740 45.230 16.000 45.550 ;
        RECT 17.180 45.210 17.320 53.390 ;
        RECT 17.640 49.970 17.780 60.530 ;
        RECT 19.420 55.090 19.680 55.410 ;
        RECT 18.040 54.750 18.300 55.070 ;
        RECT 18.100 53.710 18.240 54.750 ;
        RECT 18.040 53.390 18.300 53.710 ;
        RECT 19.480 53.030 19.620 55.090 ;
        RECT 19.420 52.710 19.680 53.030 ;
        RECT 17.580 49.650 17.840 49.970 ;
        RECT 17.580 47.950 17.840 48.270 ;
        RECT 17.640 45.890 17.780 47.950 ;
        RECT 18.960 46.590 19.220 46.910 ;
        RECT 19.020 45.890 19.160 46.590 ;
        RECT 17.580 45.570 17.840 45.890 ;
        RECT 18.960 45.570 19.220 45.890 ;
        RECT 17.120 44.890 17.380 45.210 ;
        RECT 18.040 42.170 18.300 42.490 ;
        RECT 9.580 40.615 11.460 40.985 ;
        RECT 13.440 39.110 13.700 39.430 ;
        RECT 13.900 39.110 14.160 39.430 ;
        RECT 17.580 39.110 17.840 39.430 ;
        RECT 9.760 38.430 10.020 38.750 ;
        RECT 12.980 38.430 13.240 38.750 ;
        RECT 9.820 37.390 9.960 38.430 ;
        RECT 9.760 37.070 10.020 37.390 ;
        RECT 8.380 36.390 8.640 36.710 ;
        RECT 8.440 34.570 8.580 36.390 ;
        RECT 9.580 35.175 11.460 35.545 ;
        RECT 13.040 35.010 13.180 38.430 ;
        RECT 13.500 37.730 13.640 39.110 ;
        RECT 13.440 37.410 13.700 37.730 ;
        RECT 13.960 35.010 14.100 39.110 ;
        RECT 14.820 38.430 15.080 38.750 ;
        RECT 15.740 38.430 16.000 38.750 ;
        RECT 14.880 37.390 15.020 38.430 ;
        RECT 14.820 37.070 15.080 37.390 ;
        RECT 12.980 34.690 13.240 35.010 ;
        RECT 13.900 34.690 14.160 35.010 ;
        RECT 8.440 34.430 9.040 34.570 ;
        RECT 8.900 33.990 9.040 34.430 ;
        RECT 15.800 33.990 15.940 38.430 ;
        RECT 8.840 33.670 9.100 33.990 ;
        RECT 15.740 33.670 16.000 33.990 ;
        RECT 8.900 28.890 9.040 33.670 ;
        RECT 9.580 29.735 11.460 30.105 ;
        RECT 8.840 28.570 9.100 28.890 ;
        RECT 17.120 27.890 17.380 28.210 ;
        RECT 17.180 26.850 17.320 27.890 ;
        RECT 17.120 26.530 17.380 26.850 ;
        RECT 17.640 26.170 17.780 39.110 ;
        RECT 18.100 36.710 18.240 42.170 ;
        RECT 19.420 41.830 19.680 42.150 ;
        RECT 19.480 37.730 19.620 41.830 ;
        RECT 19.940 40.110 20.080 69.030 ;
        RECT 20.860 64.930 21.000 69.030 ;
        RECT 21.320 68.670 21.460 84.670 ;
        RECT 21.780 78.190 21.920 107.110 ;
        RECT 23.100 102.350 23.360 102.670 ;
        RECT 22.640 100.990 22.900 101.310 ;
        RECT 22.700 98.930 22.840 100.990 ;
        RECT 23.160 100.290 23.300 102.350 ;
        RECT 23.100 99.970 23.360 100.290 ;
        RECT 23.100 98.950 23.360 99.270 ;
        RECT 22.640 98.610 22.900 98.930 ;
        RECT 22.180 95.550 22.440 95.870 ;
        RECT 22.240 93.830 22.380 95.550 ;
        RECT 22.180 93.510 22.440 93.830 ;
        RECT 22.240 83.290 22.380 93.510 ;
        RECT 22.700 91.450 22.840 98.610 ;
        RECT 23.160 96.890 23.300 98.950 ;
        RECT 23.100 96.570 23.360 96.890 ;
        RECT 23.100 93.850 23.360 94.170 ;
        RECT 22.640 91.130 22.900 91.450 ;
        RECT 23.160 91.110 23.300 93.850 ;
        RECT 23.100 90.790 23.360 91.110 ;
        RECT 23.160 88.730 23.300 90.790 ;
        RECT 23.100 88.410 23.360 88.730 ;
        RECT 22.640 87.390 22.900 87.710 ;
        RECT 22.180 82.970 22.440 83.290 ;
        RECT 22.700 78.530 22.840 87.390 ;
        RECT 23.100 82.630 23.360 82.950 ;
        RECT 23.160 81.250 23.300 82.630 ;
        RECT 23.100 80.930 23.360 81.250 ;
        RECT 23.100 79.910 23.360 80.230 ;
        RECT 22.640 78.210 22.900 78.530 ;
        RECT 21.720 77.870 21.980 78.190 ;
        RECT 22.640 77.530 22.900 77.850 ;
        RECT 22.180 76.850 22.440 77.170 ;
        RECT 22.240 73.090 22.380 76.850 ;
        RECT 22.180 72.770 22.440 73.090 ;
        RECT 21.720 72.430 21.980 72.750 ;
        RECT 21.780 70.030 21.920 72.430 ;
        RECT 22.180 71.070 22.440 71.390 ;
        RECT 21.720 69.710 21.980 70.030 ;
        RECT 22.240 69.690 22.380 71.070 ;
        RECT 22.180 69.370 22.440 69.690 ;
        RECT 21.260 68.350 21.520 68.670 ;
        RECT 22.180 66.650 22.440 66.970 ;
        RECT 21.720 66.310 21.980 66.630 ;
        RECT 21.260 65.970 21.520 66.290 ;
        RECT 20.800 64.610 21.060 64.930 ;
        RECT 20.800 55.430 21.060 55.750 ;
        RECT 21.320 55.490 21.460 65.970 ;
        RECT 21.780 64.930 21.920 66.310 ;
        RECT 21.720 64.610 21.980 64.930 ;
        RECT 21.780 61.190 21.920 64.610 ;
        RECT 22.240 63.230 22.380 66.650 ;
        RECT 22.180 62.910 22.440 63.230 ;
        RECT 21.720 60.870 21.980 61.190 ;
        RECT 22.240 60.510 22.380 62.910 ;
        RECT 22.180 60.190 22.440 60.510 ;
        RECT 22.180 58.150 22.440 58.470 ;
        RECT 22.240 56.090 22.380 58.150 ;
        RECT 22.180 55.770 22.440 56.090 ;
        RECT 20.340 52.090 20.600 52.350 ;
        RECT 20.860 52.090 21.000 55.430 ;
        RECT 21.320 55.410 21.920 55.490 ;
        RECT 21.320 55.350 21.980 55.410 ;
        RECT 21.320 54.050 21.460 55.350 ;
        RECT 21.720 55.090 21.980 55.350 ;
        RECT 21.260 53.730 21.520 54.050 ;
        RECT 20.340 52.030 21.000 52.090 ;
        RECT 20.400 51.950 21.000 52.030 ;
        RECT 20.860 49.630 21.000 51.950 ;
        RECT 21.320 50.310 21.460 53.730 ;
        RECT 21.720 50.670 21.980 50.990 ;
        RECT 21.260 49.990 21.520 50.310 ;
        RECT 20.800 49.310 21.060 49.630 ;
        RECT 21.260 49.310 21.520 49.630 ;
        RECT 20.860 47.590 21.000 49.310 ;
        RECT 21.320 48.270 21.460 49.310 ;
        RECT 21.260 47.950 21.520 48.270 ;
        RECT 20.800 47.270 21.060 47.590 ;
        RECT 21.780 47.500 21.920 50.670 ;
        RECT 22.240 50.650 22.380 55.770 ;
        RECT 22.180 50.330 22.440 50.650 ;
        RECT 21.320 47.360 21.920 47.500 ;
        RECT 21.320 44.870 21.460 47.360 ;
        RECT 21.260 44.550 21.520 44.870 ;
        RECT 22.700 43.170 22.840 77.530 ;
        RECT 23.160 76.830 23.300 79.910 ;
        RECT 23.620 78.530 23.760 107.450 ;
        RECT 27.300 107.090 27.440 109.490 ;
        RECT 27.240 106.770 27.500 107.090 ;
        RECT 29.540 106.430 29.800 106.750 ;
        RECT 24.580 103.175 26.460 103.545 ;
        RECT 26.780 102.010 27.040 102.330 ;
        RECT 26.840 100.290 26.980 102.010 ;
        RECT 26.780 99.970 27.040 100.290 ;
        RECT 27.240 98.950 27.500 99.270 ;
        RECT 24.020 98.270 24.280 98.590 ;
        RECT 24.080 94.170 24.220 98.270 ;
        RECT 24.580 97.735 26.460 98.105 ;
        RECT 24.020 93.850 24.280 94.170 ;
        RECT 24.580 92.295 26.460 92.665 ;
        RECT 27.300 92.130 27.440 98.950 ;
        RECT 27.240 91.810 27.500 92.130 ;
        RECT 27.240 91.130 27.500 91.450 ;
        RECT 26.780 90.110 27.040 90.430 ;
        RECT 24.020 88.070 24.280 88.390 ;
        RECT 24.080 86.690 24.220 88.070 ;
        RECT 24.580 86.855 26.460 87.225 ;
        RECT 24.020 86.370 24.280 86.690 ;
        RECT 24.080 86.010 24.220 86.370 ;
        RECT 24.020 85.690 24.280 86.010 ;
        RECT 24.580 81.415 26.460 81.785 ;
        RECT 26.840 78.530 26.980 90.110 ;
        RECT 27.300 88.390 27.440 91.130 ;
        RECT 27.240 88.070 27.500 88.390 ;
        RECT 28.620 87.390 28.880 87.710 ;
        RECT 28.160 84.670 28.420 84.990 ;
        RECT 27.700 81.950 27.960 82.270 ;
        RECT 27.760 81.250 27.900 81.950 ;
        RECT 27.700 80.930 27.960 81.250 ;
        RECT 23.560 78.210 23.820 78.530 ;
        RECT 26.780 78.210 27.040 78.530 ;
        RECT 24.020 77.530 24.280 77.850 ;
        RECT 23.560 77.190 23.820 77.510 ;
        RECT 23.100 76.510 23.360 76.830 ;
        RECT 23.160 75.130 23.300 76.510 ;
        RECT 23.100 74.810 23.360 75.130 ;
        RECT 23.100 74.130 23.360 74.450 ;
        RECT 23.160 72.070 23.300 74.130 ;
        RECT 23.100 71.750 23.360 72.070 ;
        RECT 23.620 67.650 23.760 77.190 ;
        RECT 23.560 67.330 23.820 67.650 ;
        RECT 23.100 66.540 23.360 66.630 ;
        RECT 23.100 66.400 23.760 66.540 ;
        RECT 23.100 66.310 23.360 66.400 ;
        RECT 23.100 63.930 23.360 64.250 ;
        RECT 23.160 50.990 23.300 63.930 ;
        RECT 23.620 63.570 23.760 66.400 ;
        RECT 23.560 63.250 23.820 63.570 ;
        RECT 23.620 61.530 23.760 63.250 ;
        RECT 23.560 61.210 23.820 61.530 ;
        RECT 23.100 50.670 23.360 50.990 ;
        RECT 23.160 49.970 23.300 50.670 ;
        RECT 23.100 49.650 23.360 49.970 ;
        RECT 24.080 48.010 24.220 77.530 ;
        RECT 27.700 77.190 27.960 77.510 ;
        RECT 26.780 76.850 27.040 77.170 ;
        RECT 24.580 75.975 26.460 76.345 ;
        RECT 26.840 75.810 26.980 76.850 ;
        RECT 26.780 75.490 27.040 75.810 ;
        RECT 24.940 75.150 25.200 75.470 ;
        RECT 24.480 74.130 24.740 74.450 ;
        RECT 24.540 72.070 24.680 74.130 ;
        RECT 25.000 72.750 25.140 75.150 ;
        RECT 26.320 74.810 26.580 75.130 ;
        RECT 25.400 73.790 25.660 74.110 ;
        RECT 24.940 72.430 25.200 72.750 ;
        RECT 25.460 72.070 25.600 73.790 ;
        RECT 26.380 72.070 26.520 74.810 ;
        RECT 24.480 71.925 24.740 72.070 ;
        RECT 24.470 71.555 24.750 71.925 ;
        RECT 25.400 71.750 25.660 72.070 ;
        RECT 26.320 71.750 26.580 72.070 ;
        RECT 26.770 71.555 27.050 71.925 ;
        RECT 24.580 70.535 26.460 70.905 ;
        RECT 26.840 70.370 26.980 71.555 ;
        RECT 27.240 71.070 27.500 71.390 ;
        RECT 26.780 70.050 27.040 70.370 ;
        RECT 26.320 69.370 26.580 69.690 ;
        RECT 26.380 69.010 26.520 69.370 ;
        RECT 26.320 68.690 26.580 69.010 ;
        RECT 26.380 65.950 26.520 68.690 ;
        RECT 26.780 66.650 27.040 66.970 ;
        RECT 26.320 65.630 26.580 65.950 ;
        RECT 24.580 65.095 26.460 65.465 ;
        RECT 24.480 64.610 24.740 64.930 ;
        RECT 24.540 64.250 24.680 64.610 ;
        RECT 26.840 64.330 26.980 66.650 ;
        RECT 24.480 63.930 24.740 64.250 ;
        RECT 25.860 64.160 26.120 64.250 ;
        RECT 26.380 64.190 26.980 64.330 ;
        RECT 26.380 64.160 26.520 64.190 ;
        RECT 25.860 64.020 26.520 64.160 ;
        RECT 25.860 63.930 26.120 64.020 ;
        RECT 25.920 63.570 26.060 63.930 ;
        RECT 26.780 63.590 27.040 63.910 ;
        RECT 25.860 63.250 26.120 63.570 ;
        RECT 24.580 59.655 26.460 60.025 ;
        RECT 26.840 59.490 26.980 63.590 ;
        RECT 27.300 62.210 27.440 71.070 ;
        RECT 27.760 64.930 27.900 77.190 ;
        RECT 28.220 73.090 28.360 84.670 ;
        RECT 28.160 72.770 28.420 73.090 ;
        RECT 28.160 72.090 28.420 72.410 ;
        RECT 28.220 69.690 28.360 72.090 ;
        RECT 28.160 69.370 28.420 69.690 ;
        RECT 28.680 68.670 28.820 87.390 ;
        RECT 29.080 82.290 29.340 82.610 ;
        RECT 29.140 81.250 29.280 82.290 ;
        RECT 29.080 80.930 29.340 81.250 ;
        RECT 29.600 73.090 29.740 106.430 ;
        RECT 30.460 104.730 30.720 105.050 ;
        RECT 30.000 100.990 30.260 101.310 ;
        RECT 30.060 99.270 30.200 100.990 ;
        RECT 30.000 98.950 30.260 99.270 ;
        RECT 30.000 95.550 30.260 95.870 ;
        RECT 30.060 93.490 30.200 95.550 ;
        RECT 30.520 93.570 30.660 104.730 ;
        RECT 30.920 99.290 31.180 99.610 ;
        RECT 30.980 96.550 31.120 99.290 ;
        RECT 31.380 98.950 31.640 99.270 ;
        RECT 31.440 97.570 31.580 98.950 ;
        RECT 31.380 97.250 31.640 97.570 ;
        RECT 30.920 96.230 31.180 96.550 ;
        RECT 30.000 93.170 30.260 93.490 ;
        RECT 30.520 93.430 31.120 93.570 ;
        RECT 30.460 92.830 30.720 93.150 ;
        RECT 30.520 92.130 30.660 92.830 ;
        RECT 30.460 91.810 30.720 92.130 ;
        RECT 30.000 85.350 30.260 85.670 ;
        RECT 30.060 83.970 30.200 85.350 ;
        RECT 30.000 83.650 30.260 83.970 ;
        RECT 30.060 80.570 30.200 83.650 ;
        RECT 30.000 80.250 30.260 80.570 ;
        RECT 29.540 72.770 29.800 73.090 ;
        RECT 29.080 71.750 29.340 72.070 ;
        RECT 28.620 68.350 28.880 68.670 ;
        RECT 28.620 66.310 28.880 66.630 ;
        RECT 27.700 64.610 27.960 64.930 ;
        RECT 27.240 61.890 27.500 62.210 ;
        RECT 26.780 59.170 27.040 59.490 ;
        RECT 26.840 55.490 26.980 59.170 ;
        RECT 28.160 57.470 28.420 57.790 ;
        RECT 27.240 55.770 27.500 56.090 ;
        RECT 26.380 55.350 26.980 55.490 ;
        RECT 26.380 55.070 26.520 55.350 ;
        RECT 26.320 54.750 26.580 55.070 ;
        RECT 24.580 54.215 26.460 54.585 ;
        RECT 26.840 54.050 26.980 55.350 ;
        RECT 27.300 54.050 27.440 55.770 ;
        RECT 26.780 53.730 27.040 54.050 ;
        RECT 27.240 53.730 27.500 54.050 ;
        RECT 28.220 53.370 28.360 57.470 ;
        RECT 28.160 53.050 28.420 53.370 ;
        RECT 28.680 50.310 28.820 66.310 ;
        RECT 28.620 49.990 28.880 50.310 ;
        RECT 28.160 49.650 28.420 49.970 ;
        RECT 24.580 48.775 26.460 49.145 ;
        RECT 28.220 48.805 28.360 49.650 ;
        RECT 28.150 48.435 28.430 48.805 ;
        RECT 23.160 47.870 24.220 48.010 ;
        RECT 22.640 42.850 22.900 43.170 ;
        RECT 20.800 42.170 21.060 42.490 ;
        RECT 20.860 41.470 21.000 42.170 ;
        RECT 20.800 41.150 21.060 41.470 ;
        RECT 22.640 41.150 22.900 41.470 ;
        RECT 19.880 39.790 20.140 40.110 ;
        RECT 22.700 39.430 22.840 41.150 ;
        RECT 23.160 40.450 23.300 47.870 ;
        RECT 23.560 47.270 23.820 47.590 ;
        RECT 23.620 45.210 23.760 47.270 ;
        RECT 23.560 45.120 23.820 45.210 ;
        RECT 23.560 44.980 24.220 45.120 ;
        RECT 23.560 44.890 23.820 44.980 ;
        RECT 23.560 41.830 23.820 42.150 ;
        RECT 23.100 40.130 23.360 40.450 ;
        RECT 22.640 39.110 22.900 39.430 ;
        RECT 21.260 38.770 21.520 39.090 ;
        RECT 19.420 37.410 19.680 37.730 ;
        RECT 18.040 36.390 18.300 36.710 ;
        RECT 19.480 32.290 19.620 37.410 ;
        RECT 21.320 37.050 21.460 38.770 ;
        RECT 21.260 36.730 21.520 37.050 ;
        RECT 20.800 35.710 21.060 36.030 ;
        RECT 20.860 33.990 21.000 35.710 ;
        RECT 21.320 34.330 21.460 36.730 ;
        RECT 22.180 36.390 22.440 36.710 ;
        RECT 23.620 36.450 23.760 41.830 ;
        RECT 22.240 34.330 22.380 36.390 ;
        RECT 23.160 36.310 23.760 36.450 ;
        RECT 21.260 34.010 21.520 34.330 ;
        RECT 22.180 34.010 22.440 34.330 ;
        RECT 20.800 33.670 21.060 33.990 ;
        RECT 19.420 31.970 19.680 32.290 ;
        RECT 18.040 28.570 18.300 28.890 ;
        RECT 18.100 26.170 18.240 28.570 ;
        RECT 19.480 27.870 19.620 31.970 ;
        RECT 22.240 31.270 22.380 34.010 ;
        RECT 22.180 30.950 22.440 31.270 ;
        RECT 19.880 30.270 20.140 30.590 ;
        RECT 19.940 28.550 20.080 30.270 ;
        RECT 23.160 28.550 23.300 36.310 ;
        RECT 23.560 35.710 23.820 36.030 ;
        RECT 23.620 31.610 23.760 35.710 ;
        RECT 24.080 33.990 24.220 44.980 ;
        RECT 24.580 43.335 26.460 43.705 ;
        RECT 29.140 43.170 29.280 71.750 ;
        RECT 30.980 70.370 31.120 93.430 ;
        RECT 31.840 90.110 32.100 90.430 ;
        RECT 31.380 73.790 31.640 74.110 ;
        RECT 31.440 72.070 31.580 73.790 ;
        RECT 31.900 73.090 32.040 90.110 ;
        RECT 32.300 85.690 32.560 86.010 ;
        RECT 32.360 81.250 32.500 85.690 ;
        RECT 32.820 85.580 32.960 109.830 ;
        RECT 33.280 108.110 33.420 109.830 ;
        RECT 35.580 109.470 35.720 115.610 ;
        RECT 35.980 109.490 36.240 109.810 ;
        RECT 35.520 109.150 35.780 109.470 ;
        RECT 36.040 108.450 36.180 109.490 ;
        RECT 39.260 109.470 39.400 128.790 ;
        RECT 39.580 116.775 41.460 117.145 ;
        RECT 41.960 115.270 42.220 115.590 ;
        RECT 42.020 112.190 42.160 115.270 ;
        RECT 44.780 113.970 44.920 128.280 ;
        RECT 44.320 113.890 44.920 113.970 ;
        RECT 44.260 113.830 44.920 113.890 ;
        RECT 44.260 113.570 44.520 113.830 ;
        RECT 44.720 113.230 44.980 113.550 ;
        RECT 42.420 112.550 42.680 112.870 ;
        RECT 41.960 111.870 42.220 112.190 ;
        RECT 39.580 111.335 41.460 111.705 ;
        RECT 42.020 110.490 42.160 111.870 ;
        RECT 41.960 110.170 42.220 110.490 ;
        RECT 41.040 109.490 41.300 109.810 ;
        RECT 39.200 109.150 39.460 109.470 ;
        RECT 41.100 108.450 41.240 109.490 ;
        RECT 35.980 108.130 36.240 108.450 ;
        RECT 41.040 108.130 41.300 108.450 ;
        RECT 33.220 107.790 33.480 108.110 ;
        RECT 39.580 105.895 41.460 106.265 ;
        RECT 35.520 103.710 35.780 104.030 ;
        RECT 35.580 102.670 35.720 103.710 ;
        RECT 35.520 102.350 35.780 102.670 ;
        RECT 42.020 101.990 42.160 110.170 ;
        RECT 42.480 108.450 42.620 112.550 ;
        RECT 44.780 108.450 44.920 113.230 ;
        RECT 47.020 112.550 47.280 112.870 ;
        RECT 49.320 112.550 49.580 112.870 ;
        RECT 47.080 110.490 47.220 112.550 ;
        RECT 47.020 110.170 47.280 110.490 ;
        RECT 45.180 109.830 45.440 110.150 ;
        RECT 42.420 108.130 42.680 108.450 ;
        RECT 44.720 108.130 44.980 108.450 ;
        RECT 42.880 104.390 43.140 104.710 ;
        RECT 42.940 102.330 43.080 104.390 ;
        RECT 42.880 102.010 43.140 102.330 ;
        RECT 41.960 101.670 42.220 101.990 ;
        RECT 33.680 100.990 33.940 101.310 ;
        RECT 39.200 100.990 39.460 101.310 ;
        RECT 33.740 97.230 33.880 100.990 ;
        RECT 39.260 98.930 39.400 100.990 ;
        RECT 39.580 100.455 41.460 100.825 ;
        RECT 42.020 99.610 42.160 101.670 ;
        RECT 41.960 99.290 42.220 99.610 ;
        RECT 42.420 98.950 42.680 99.270 ;
        RECT 39.200 98.610 39.460 98.930 ;
        RECT 41.500 98.610 41.760 98.930 ;
        RECT 41.560 97.570 41.700 98.610 ;
        RECT 41.500 97.250 41.760 97.570 ;
        RECT 33.680 96.910 33.940 97.230 ;
        RECT 38.740 96.910 39.000 97.230 ;
        RECT 33.740 91.450 33.880 96.910 ;
        RECT 37.820 96.570 38.080 96.890 ;
        RECT 37.880 91.790 38.020 96.570 ;
        RECT 38.800 94.850 38.940 96.910 ;
        RECT 41.960 96.230 42.220 96.550 ;
        RECT 39.580 95.015 41.460 95.385 ;
        RECT 38.740 94.530 39.000 94.850 ;
        RECT 41.040 92.830 41.300 93.150 ;
        RECT 41.100 91.790 41.240 92.830 ;
        RECT 37.820 91.470 38.080 91.790 ;
        RECT 41.040 91.470 41.300 91.790 ;
        RECT 33.220 91.130 33.480 91.450 ;
        RECT 33.680 91.130 33.940 91.450 ;
        RECT 33.280 88.730 33.420 91.130 ;
        RECT 42.020 91.110 42.160 96.230 ;
        RECT 42.480 94.850 42.620 98.950 ;
        RECT 42.420 94.530 42.680 94.850 ;
        RECT 42.940 93.830 43.080 102.010 ;
        RECT 44.720 98.270 44.980 98.590 ;
        RECT 44.780 96.890 44.920 98.270 ;
        RECT 44.720 96.570 44.980 96.890 ;
        RECT 42.880 93.510 43.140 93.830 ;
        RECT 41.960 90.790 42.220 91.110 ;
        RECT 39.580 89.575 41.460 89.945 ;
        RECT 33.220 88.410 33.480 88.730 ;
        RECT 38.740 87.390 39.000 87.710 ;
        RECT 38.800 86.010 38.940 87.390 ;
        RECT 42.420 86.030 42.680 86.350 ;
        RECT 37.360 85.690 37.620 86.010 ;
        RECT 38.740 85.690 39.000 86.010 ;
        RECT 32.820 85.440 33.420 85.580 ;
        RECT 32.760 84.670 33.020 84.990 ;
        RECT 32.820 83.290 32.960 84.670 ;
        RECT 32.760 82.970 33.020 83.290 ;
        RECT 32.300 80.930 32.560 81.250 ;
        RECT 33.280 73.090 33.420 85.440 ;
        RECT 36.900 85.350 37.160 85.670 ;
        RECT 35.520 84.670 35.780 84.990 ;
        RECT 34.600 83.650 34.860 83.970 ;
        RECT 34.140 81.950 34.400 82.270 ;
        RECT 34.200 80.570 34.340 81.950 ;
        RECT 34.660 81.250 34.800 83.650 ;
        RECT 35.580 82.610 35.720 84.670 ;
        RECT 36.960 83.290 37.100 85.350 ;
        RECT 36.900 82.970 37.160 83.290 ;
        RECT 35.520 82.290 35.780 82.610 ;
        RECT 34.600 80.930 34.860 81.250 ;
        RECT 34.140 80.250 34.400 80.570 ;
        RECT 34.200 75.130 34.340 80.250 ;
        RECT 33.680 74.810 33.940 75.130 ;
        RECT 34.140 74.810 34.400 75.130 ;
        RECT 35.060 74.810 35.320 75.130 ;
        RECT 31.840 72.770 32.100 73.090 ;
        RECT 33.220 72.770 33.480 73.090 ;
        RECT 33.740 72.750 33.880 74.810 ;
        RECT 34.600 74.470 34.860 74.790 ;
        RECT 33.680 72.430 33.940 72.750 ;
        RECT 34.660 72.410 34.800 74.470 ;
        RECT 32.300 72.090 32.560 72.410 ;
        RECT 34.600 72.090 34.860 72.410 ;
        RECT 31.380 71.750 31.640 72.070 ;
        RECT 30.920 70.050 31.180 70.370 ;
        RECT 29.540 69.030 29.800 69.350 ;
        RECT 29.600 43.170 29.740 69.030 ;
        RECT 30.000 66.310 30.260 66.630 ;
        RECT 30.060 64.250 30.200 66.310 ;
        RECT 30.000 63.930 30.260 64.250 ;
        RECT 30.000 55.090 30.260 55.410 ;
        RECT 30.060 54.050 30.200 55.090 ;
        RECT 30.000 53.730 30.260 54.050 ;
        RECT 31.840 53.050 32.100 53.370 ;
        RECT 30.920 50.670 31.180 50.990 ;
        RECT 30.980 50.310 31.120 50.670 ;
        RECT 30.920 49.990 31.180 50.310 ;
        RECT 30.980 45.890 31.120 49.990 ;
        RECT 30.920 45.570 31.180 45.890 ;
        RECT 31.900 44.870 32.040 53.050 ;
        RECT 31.840 44.550 32.100 44.870 ;
        RECT 32.360 43.170 32.500 72.090 ;
        RECT 33.680 71.750 33.940 72.070 ;
        RECT 35.120 71.925 35.260 74.810 ;
        RECT 36.960 74.790 37.100 82.970 ;
        RECT 37.420 82.950 37.560 85.690 ;
        RECT 39.580 84.135 41.460 84.505 ;
        RECT 42.480 82.950 42.620 86.030 ;
        RECT 44.720 84.670 44.980 84.990 ;
        RECT 37.360 82.630 37.620 82.950 ;
        RECT 42.420 82.630 42.680 82.950 ;
        RECT 41.960 82.290 42.220 82.610 ;
        RECT 39.200 79.230 39.460 79.550 ;
        RECT 39.260 75.130 39.400 79.230 ;
        RECT 39.580 78.695 41.460 79.065 ;
        RECT 42.020 77.510 42.160 82.290 ;
        RECT 44.780 81.250 44.920 84.670 ;
        RECT 44.720 80.930 44.980 81.250 ;
        RECT 45.240 80.650 45.380 109.830 ;
        RECT 49.380 108.450 49.520 112.550 ;
        RECT 50.760 110.490 50.900 128.280 ;
        RECT 51.160 115.270 51.420 115.590 ;
        RECT 50.700 110.170 50.960 110.490 ;
        RECT 49.320 108.130 49.580 108.450 ;
        RECT 51.220 108.110 51.360 115.270 ;
        RECT 51.620 114.590 51.880 114.910 ;
        RECT 53.000 114.590 53.260 114.910 ;
        RECT 51.680 109.810 51.820 114.590 ;
        RECT 53.060 113.550 53.200 114.590 ;
        RECT 54.580 114.055 56.460 114.425 ;
        RECT 56.740 113.890 56.880 128.280 ;
        RECT 57.140 114.930 57.400 115.250 ;
        RECT 56.680 113.570 56.940 113.890 ;
        RECT 53.000 113.230 53.260 113.550 ;
        RECT 57.200 110.150 57.340 114.930 ;
        RECT 62.200 111.870 62.460 112.190 ;
        RECT 62.260 110.490 62.400 111.870 ;
        RECT 62.720 110.490 62.860 128.280 ;
        RECT 68.700 113.890 68.840 128.280 ;
        RECT 69.580 116.775 71.460 117.145 ;
        RECT 74.680 113.890 74.820 128.280 ;
        RECT 68.640 113.570 68.900 113.890 ;
        RECT 74.620 113.570 74.880 113.890 ;
        RECT 76.000 113.230 76.260 113.550 ;
        RECT 69.100 112.890 69.360 113.210 ;
        RECT 63.580 112.550 63.840 112.870 ;
        RECT 63.640 111.170 63.780 112.550 ;
        RECT 69.160 111.170 69.300 112.890 ;
        RECT 72.780 112.550 73.040 112.870 ;
        RECT 69.580 111.335 71.460 111.705 ;
        RECT 72.840 111.170 72.980 112.550 ;
        RECT 73.240 111.870 73.500 112.190 ;
        RECT 63.580 110.850 63.840 111.170 ;
        RECT 69.100 110.850 69.360 111.170 ;
        RECT 72.780 110.850 73.040 111.170 ;
        RECT 73.300 110.490 73.440 111.870 ;
        RECT 73.700 110.850 73.960 111.170 ;
        RECT 62.200 110.170 62.460 110.490 ;
        RECT 62.660 110.170 62.920 110.490 ;
        RECT 73.240 110.170 73.500 110.490 ;
        RECT 57.140 109.830 57.400 110.150 ;
        RECT 65.880 109.830 66.140 110.150 ;
        RECT 69.100 109.830 69.360 110.150 ;
        RECT 69.560 109.830 69.820 110.150 ;
        RECT 51.620 109.490 51.880 109.810 ;
        RECT 61.740 109.150 62.000 109.470 ;
        RECT 62.200 109.150 62.460 109.470 ;
        RECT 54.580 108.615 56.460 108.985 ;
        RECT 51.160 107.790 51.420 108.110 ;
        RECT 61.800 107.850 61.940 109.150 ;
        RECT 62.260 108.450 62.400 109.150 ;
        RECT 65.940 108.450 66.080 109.830 ;
        RECT 62.200 108.130 62.460 108.450 ;
        RECT 65.880 108.130 66.140 108.450 ;
        RECT 69.160 108.110 69.300 109.830 ;
        RECT 53.000 107.450 53.260 107.770 ;
        RECT 61.800 107.710 62.400 107.850 ;
        RECT 68.180 107.790 68.440 108.110 ;
        RECT 69.100 107.790 69.360 108.110 ;
        RECT 48.860 106.430 49.120 106.750 ;
        RECT 47.940 104.730 48.200 105.050 ;
        RECT 46.560 103.710 46.820 104.030 ;
        RECT 47.480 103.710 47.740 104.030 ;
        RECT 45.640 101.670 45.900 101.990 ;
        RECT 45.700 100.290 45.840 101.670 ;
        RECT 45.640 99.970 45.900 100.290 ;
        RECT 46.100 99.290 46.360 99.610 ;
        RECT 46.160 97.230 46.300 99.290 ;
        RECT 46.620 99.270 46.760 103.710 ;
        RECT 47.540 99.270 47.680 103.710 ;
        RECT 46.560 98.950 46.820 99.270 ;
        RECT 47.480 98.950 47.740 99.270 ;
        RECT 46.560 98.270 46.820 98.590 ;
        RECT 46.100 96.910 46.360 97.230 ;
        RECT 46.620 94.170 46.760 98.270 ;
        RECT 47.010 96.715 47.290 97.085 ;
        RECT 47.020 96.570 47.280 96.715 ;
        RECT 46.560 93.850 46.820 94.170 ;
        RECT 47.540 91.110 47.680 98.950 ;
        RECT 48.000 96.550 48.140 104.730 ;
        RECT 47.940 96.230 48.200 96.550 ;
        RECT 48.000 94.170 48.140 96.230 ;
        RECT 47.940 93.850 48.200 94.170 ;
        RECT 47.480 90.790 47.740 91.110 ;
        RECT 48.920 89.410 49.060 106.430 ;
        RECT 51.620 104.050 51.880 104.370 ;
        RECT 49.320 102.350 49.580 102.670 ;
        RECT 49.380 94.850 49.520 102.350 ;
        RECT 51.680 101.310 51.820 104.050 ;
        RECT 51.620 100.990 51.880 101.310 ;
        RECT 49.320 94.530 49.580 94.850 ;
        RECT 51.680 94.170 51.820 100.990 ;
        RECT 52.540 98.610 52.800 98.930 ;
        RECT 52.600 97.570 52.740 98.610 ;
        RECT 52.540 97.250 52.800 97.570 ;
        RECT 51.160 93.850 51.420 94.170 ;
        RECT 51.620 93.850 51.880 94.170 ;
        RECT 51.220 92.130 51.360 93.850 ;
        RECT 51.160 91.810 51.420 92.130 ;
        RECT 51.680 91.360 51.820 93.850 ;
        RECT 52.540 92.830 52.800 93.150 ;
        RECT 52.080 91.360 52.340 91.450 ;
        RECT 51.680 91.220 52.340 91.360 ;
        RECT 52.080 91.130 52.340 91.220 ;
        RECT 50.700 90.110 50.960 90.430 ;
        RECT 51.620 90.110 51.880 90.430 ;
        RECT 48.860 89.090 49.120 89.410 ;
        RECT 49.780 88.410 50.040 88.730 ;
        RECT 46.560 88.070 46.820 88.390 ;
        RECT 49.320 88.070 49.580 88.390 ;
        RECT 46.620 86.690 46.760 88.070 ;
        RECT 47.020 87.730 47.280 88.050 ;
        RECT 46.560 86.370 46.820 86.690 ;
        RECT 47.080 83.970 47.220 87.730 ;
        RECT 47.940 85.690 48.200 86.010 ;
        RECT 47.480 85.350 47.740 85.670 ;
        RECT 47.020 83.650 47.280 83.970 ;
        RECT 47.020 82.970 47.280 83.290 ;
        RECT 45.240 80.510 45.840 80.650 ;
        RECT 45.180 79.910 45.440 80.230 ;
        RECT 41.960 77.190 42.220 77.510 ;
        RECT 44.720 77.190 44.980 77.510 ;
        RECT 41.500 76.510 41.760 76.830 ;
        RECT 41.560 75.470 41.700 76.510 ;
        RECT 41.500 75.150 41.760 75.470 ;
        RECT 39.200 74.810 39.460 75.130 ;
        RECT 36.900 74.470 37.160 74.790 ;
        RECT 39.580 73.255 41.460 73.625 ;
        RECT 43.340 72.090 43.600 72.410 ;
        RECT 33.220 69.370 33.480 69.690 ;
        RECT 33.280 67.650 33.420 69.370 ;
        RECT 33.220 67.330 33.480 67.650 ;
        RECT 33.220 66.650 33.480 66.970 ;
        RECT 32.760 66.310 33.020 66.630 ;
        RECT 32.820 56.090 32.960 66.310 ;
        RECT 33.280 64.330 33.420 66.650 ;
        RECT 33.740 64.930 33.880 71.750 ;
        RECT 35.050 71.555 35.330 71.925 ;
        RECT 41.500 71.410 41.760 71.730 ;
        RECT 42.880 71.410 43.140 71.730 ;
        RECT 41.560 70.030 41.700 71.410 ;
        RECT 42.940 70.370 43.080 71.410 ;
        RECT 43.400 70.370 43.540 72.090 ;
        RECT 44.260 71.070 44.520 71.390 ;
        RECT 42.880 70.050 43.140 70.370 ;
        RECT 43.340 70.050 43.600 70.370 ;
        RECT 41.500 69.710 41.760 70.030 ;
        RECT 44.320 69.690 44.460 71.070 ;
        RECT 44.780 69.690 44.920 77.190 ;
        RECT 45.240 74.790 45.380 79.910 ;
        RECT 45.700 75.810 45.840 80.510 ;
        RECT 47.080 77.850 47.220 82.970 ;
        RECT 47.540 80.230 47.680 85.350 ;
        RECT 48.000 83.630 48.140 85.690 ;
        RECT 47.940 83.310 48.200 83.630 ;
        RECT 47.480 79.910 47.740 80.230 ;
        RECT 47.020 77.530 47.280 77.850 ;
        RECT 45.640 75.490 45.900 75.810 ;
        RECT 45.180 74.470 45.440 74.790 ;
        RECT 45.240 72.070 45.380 74.470 ;
        RECT 47.540 74.020 47.680 79.910 ;
        RECT 47.940 74.810 48.200 75.130 ;
        RECT 48.000 74.530 48.140 74.810 ;
        RECT 48.000 74.390 48.600 74.530 ;
        RECT 47.540 73.880 48.140 74.020 ;
        RECT 48.000 72.410 48.140 73.880 ;
        RECT 48.460 72.410 48.600 74.390 ;
        RECT 47.940 72.090 48.200 72.410 ;
        RECT 48.400 72.090 48.660 72.410 ;
        RECT 45.180 71.750 45.440 72.070 ;
        RECT 44.260 69.370 44.520 69.690 ;
        RECT 44.720 69.370 44.980 69.690 ;
        RECT 48.000 69.350 48.140 72.090 ;
        RECT 47.940 69.030 48.200 69.350 ;
        RECT 42.880 68.690 43.140 69.010 ;
        RECT 35.520 68.350 35.780 68.670 ;
        RECT 35.580 66.970 35.720 68.350 ;
        RECT 39.580 67.815 41.460 68.185 ;
        RECT 42.940 67.650 43.080 68.690 ;
        RECT 42.880 67.330 43.140 67.650 ;
        RECT 35.520 66.650 35.780 66.970 ;
        RECT 35.980 66.650 36.240 66.970 ;
        RECT 36.040 65.950 36.180 66.650 ;
        RECT 39.200 65.970 39.460 66.290 ;
        RECT 48.860 65.970 49.120 66.290 ;
        RECT 35.980 65.630 36.240 65.950 ;
        RECT 33.680 64.610 33.940 64.930 ;
        RECT 33.280 64.250 33.880 64.330 ;
        RECT 36.040 64.250 36.180 65.630 ;
        RECT 39.260 64.930 39.400 65.970 ;
        RECT 39.200 64.610 39.460 64.930 ;
        RECT 33.280 64.190 33.940 64.250 ;
        RECT 33.680 63.930 33.940 64.190 ;
        RECT 34.140 63.930 34.400 64.250 ;
        RECT 35.980 63.930 36.240 64.250 ;
        RECT 43.800 63.930 44.060 64.250 ;
        RECT 33.740 63.230 33.880 63.930 ;
        RECT 33.680 62.910 33.940 63.230 ;
        RECT 34.200 59.490 34.340 63.930 ;
        RECT 39.580 62.375 41.460 62.745 ;
        RECT 43.340 60.530 43.600 60.850 ;
        RECT 43.400 59.490 43.540 60.530 ;
        RECT 34.140 59.170 34.400 59.490 ;
        RECT 43.340 59.170 43.600 59.490 ;
        RECT 34.200 56.770 34.340 59.170 ;
        RECT 43.860 58.810 44.000 63.930 ;
        RECT 44.720 60.870 44.980 61.190 ;
        RECT 44.260 60.190 44.520 60.510 ;
        RECT 44.320 59.490 44.460 60.190 ;
        RECT 44.260 59.170 44.520 59.490 ;
        RECT 43.800 58.490 44.060 58.810 ;
        RECT 36.900 58.150 37.160 58.470 ;
        RECT 35.520 57.470 35.780 57.790 ;
        RECT 34.140 56.450 34.400 56.770 ;
        RECT 32.760 55.770 33.020 56.090 ;
        RECT 32.820 47.930 32.960 55.770 ;
        RECT 34.600 55.430 34.860 55.750 ;
        RECT 34.660 54.050 34.800 55.430 ;
        RECT 34.600 53.730 34.860 54.050 ;
        RECT 35.580 53.370 35.720 57.470 ;
        RECT 36.960 56.770 37.100 58.150 ;
        RECT 39.580 56.935 41.460 57.305 ;
        RECT 36.900 56.450 37.160 56.770 ;
        RECT 37.360 55.090 37.620 55.410 ;
        RECT 37.420 54.050 37.560 55.090 ;
        RECT 37.360 53.730 37.620 54.050 ;
        RECT 43.860 53.370 44.000 58.490 ;
        RECT 35.520 53.050 35.780 53.370 ;
        RECT 43.800 53.050 44.060 53.370 ;
        RECT 39.580 51.495 41.460 51.865 ;
        RECT 41.960 49.650 42.220 49.970 ;
        RECT 34.600 49.310 34.860 49.630 ;
        RECT 32.760 47.610 33.020 47.930 ;
        RECT 34.660 47.590 34.800 49.310 ;
        RECT 35.980 47.950 36.240 48.270 ;
        RECT 34.600 47.270 34.860 47.590 ;
        RECT 33.680 46.590 33.940 46.910 ;
        RECT 33.220 45.230 33.480 45.550 ;
        RECT 29.080 42.850 29.340 43.170 ;
        RECT 29.540 42.850 29.800 43.170 ;
        RECT 32.300 42.850 32.560 43.170 ;
        RECT 33.280 42.490 33.420 45.230 ;
        RECT 33.740 42.490 33.880 46.590 ;
        RECT 36.040 44.870 36.180 47.950 ;
        RECT 42.020 47.590 42.160 49.650 ;
        RECT 43.860 47.930 44.000 53.050 ;
        RECT 44.780 53.030 44.920 60.870 ;
        RECT 48.920 60.510 49.060 65.970 ;
        RECT 48.860 60.190 49.120 60.510 ;
        RECT 48.920 59.490 49.060 60.190 ;
        RECT 49.380 59.490 49.520 88.070 ;
        RECT 49.840 83.630 49.980 88.410 ;
        RECT 50.240 85.690 50.500 86.010 ;
        RECT 49.780 83.310 50.040 83.630 ;
        RECT 50.300 82.950 50.440 85.690 ;
        RECT 50.240 82.630 50.500 82.950 ;
        RECT 49.780 75.490 50.040 75.810 ;
        RECT 49.840 74.450 49.980 75.490 ;
        RECT 49.780 74.130 50.040 74.450 ;
        RECT 49.840 71.980 49.980 74.130 ;
        RECT 50.300 72.750 50.440 82.630 ;
        RECT 50.240 72.430 50.500 72.750 ;
        RECT 50.240 71.980 50.500 72.070 ;
        RECT 49.840 71.840 50.500 71.980 ;
        RECT 49.840 63.765 49.980 71.840 ;
        RECT 50.240 71.750 50.500 71.840 ;
        RECT 50.240 71.070 50.500 71.390 ;
        RECT 50.300 70.030 50.440 71.070 ;
        RECT 50.240 69.710 50.500 70.030 ;
        RECT 50.760 68.670 50.900 90.110 ;
        RECT 51.680 89.410 51.820 90.110 ;
        RECT 51.620 89.090 51.880 89.410 ;
        RECT 51.160 88.925 51.420 89.070 ;
        RECT 51.150 88.555 51.430 88.925 ;
        RECT 52.600 88.640 52.740 92.830 ;
        RECT 51.680 88.500 52.740 88.640 ;
        RECT 51.160 88.070 51.420 88.390 ;
        RECT 51.220 77.850 51.360 88.070 ;
        RECT 51.160 77.530 51.420 77.850 ;
        RECT 51.150 76.995 51.430 77.365 ;
        RECT 51.220 74.790 51.360 76.995 ;
        RECT 51.680 74.790 51.820 88.500 ;
        RECT 53.060 88.130 53.200 107.450 ;
        RECT 57.140 106.770 57.400 107.090 ;
        RECT 54.580 103.175 56.460 103.545 ;
        RECT 53.920 102.010 54.180 102.330 ;
        RECT 53.460 99.290 53.720 99.610 ;
        RECT 53.520 97.230 53.660 99.290 ;
        RECT 53.460 96.910 53.720 97.230 ;
        RECT 53.520 96.210 53.660 96.910 ;
        RECT 53.460 95.890 53.720 96.210 ;
        RECT 53.520 88.390 53.660 95.890 ;
        RECT 53.980 94.850 54.120 102.010 ;
        RECT 54.380 100.990 54.640 101.310 ;
        RECT 54.440 99.270 54.580 100.990 ;
        RECT 54.380 98.950 54.640 99.270 ;
        RECT 54.580 97.735 56.460 98.105 ;
        RECT 53.920 94.530 54.180 94.850 ;
        RECT 53.920 93.510 54.180 93.830 ;
        RECT 53.980 91.450 54.120 93.510 ;
        RECT 54.580 92.295 56.460 92.665 ;
        RECT 53.920 91.130 54.180 91.450 ;
        RECT 53.920 90.110 54.180 90.430 ;
        RECT 52.600 87.990 53.200 88.130 ;
        RECT 53.460 88.070 53.720 88.390 ;
        RECT 52.070 85.835 52.350 86.205 ;
        RECT 52.080 85.690 52.340 85.835 ;
        RECT 52.140 82.610 52.280 85.690 ;
        RECT 52.080 82.290 52.340 82.610 ;
        RECT 52.140 75.810 52.280 82.290 ;
        RECT 52.080 75.490 52.340 75.810 ;
        RECT 51.160 74.470 51.420 74.790 ;
        RECT 51.620 74.470 51.880 74.790 ;
        RECT 52.080 74.470 52.340 74.790 ;
        RECT 51.220 72.070 51.360 74.470 ;
        RECT 51.620 73.790 51.880 74.110 ;
        RECT 51.680 72.605 51.820 73.790 ;
        RECT 51.610 72.235 51.890 72.605 ;
        RECT 51.160 71.750 51.420 72.070 ;
        RECT 51.620 71.410 51.880 71.730 ;
        RECT 51.680 70.370 51.820 71.410 ;
        RECT 51.620 70.050 51.880 70.370 ;
        RECT 51.620 69.370 51.880 69.690 ;
        RECT 51.160 69.030 51.420 69.350 ;
        RECT 50.700 68.350 50.960 68.670 ;
        RECT 50.700 66.990 50.960 67.310 ;
        RECT 50.240 66.310 50.500 66.630 ;
        RECT 50.300 64.590 50.440 66.310 ;
        RECT 50.240 64.270 50.500 64.590 ;
        RECT 50.760 64.250 50.900 66.990 ;
        RECT 50.700 63.930 50.960 64.250 ;
        RECT 49.770 63.395 50.050 63.765 ;
        RECT 50.760 61.190 50.900 63.930 ;
        RECT 50.700 60.870 50.960 61.190 ;
        RECT 48.860 59.170 49.120 59.490 ;
        RECT 49.320 59.170 49.580 59.490 ;
        RECT 47.020 58.490 47.280 58.810 ;
        RECT 47.080 56.770 47.220 58.490 ;
        RECT 47.020 56.450 47.280 56.770 ;
        RECT 48.920 55.750 49.060 59.170 ;
        RECT 50.760 59.150 50.900 60.870 ;
        RECT 50.700 58.830 50.960 59.150 ;
        RECT 49.780 58.150 50.040 58.470 ;
        RECT 49.840 56.090 49.980 58.150 ;
        RECT 49.780 55.770 50.040 56.090 ;
        RECT 48.860 55.430 49.120 55.750 ;
        RECT 47.020 54.750 47.280 55.070 ;
        RECT 47.080 53.370 47.220 54.750 ;
        RECT 47.020 53.050 47.280 53.370 ;
        RECT 44.720 52.710 44.980 53.030 ;
        RECT 44.780 50.310 44.920 52.710 ;
        RECT 44.720 49.990 44.980 50.310 ;
        RECT 43.340 47.610 43.600 47.930 ;
        RECT 43.800 47.610 44.060 47.930 ;
        RECT 41.960 47.270 42.220 47.590 ;
        RECT 42.420 46.930 42.680 47.250 ;
        RECT 39.580 46.055 41.460 46.425 ;
        RECT 35.980 44.550 36.240 44.870 ;
        RECT 38.280 44.550 38.540 44.870 ;
        RECT 38.340 42.830 38.480 44.550 ;
        RECT 42.480 43.170 42.620 46.930 ;
        RECT 43.400 44.530 43.540 47.610 ;
        RECT 44.780 44.870 44.920 49.990 ;
        RECT 49.320 49.650 49.580 49.970 ;
        RECT 49.380 48.270 49.520 49.650 ;
        RECT 47.010 47.755 47.290 48.125 ;
        RECT 49.320 47.950 49.580 48.270 ;
        RECT 44.720 44.550 44.980 44.870 ;
        RECT 43.340 44.210 43.600 44.530 ;
        RECT 42.420 42.850 42.680 43.170 ;
        RECT 38.280 42.510 38.540 42.830 ;
        RECT 26.320 42.170 26.580 42.490 ;
        RECT 28.160 42.170 28.420 42.490 ;
        RECT 33.220 42.170 33.480 42.490 ;
        RECT 33.680 42.170 33.940 42.490 ;
        RECT 34.140 42.170 34.400 42.490 ;
        RECT 26.380 41.470 26.520 42.170 ;
        RECT 26.320 41.150 26.580 41.470 ;
        RECT 27.700 39.340 27.960 39.430 ;
        RECT 28.220 39.340 28.360 42.170 ;
        RECT 29.080 41.830 29.340 42.150 ;
        RECT 29.140 39.770 29.280 41.830 ;
        RECT 29.540 41.490 29.800 41.810 ;
        RECT 29.080 39.450 29.340 39.770 ;
        RECT 29.600 39.430 29.740 41.490 ;
        RECT 27.700 39.200 28.360 39.340 ;
        RECT 27.700 39.110 27.960 39.200 ;
        RECT 29.540 39.110 29.800 39.430 ;
        RECT 27.240 38.770 27.500 39.090 ;
        RECT 30.000 38.770 30.260 39.090 ;
        RECT 24.580 37.895 26.460 38.265 ;
        RECT 24.020 33.670 24.280 33.990 ;
        RECT 23.560 31.290 23.820 31.610 ;
        RECT 24.080 28.890 24.220 33.670 ;
        RECT 26.780 33.330 27.040 33.650 ;
        RECT 24.580 32.455 26.460 32.825 ;
        RECT 26.840 32.290 26.980 33.330 ;
        RECT 26.780 31.970 27.040 32.290 ;
        RECT 27.300 31.950 27.440 38.770 ;
        RECT 30.060 37.730 30.200 38.770 ;
        RECT 30.000 37.410 30.260 37.730 ;
        RECT 34.200 37.050 34.340 42.170 ;
        RECT 35.520 41.490 35.780 41.810 ;
        RECT 35.580 39.090 35.720 41.490 ;
        RECT 38.340 39.770 38.480 42.510 ;
        RECT 43.400 42.490 43.540 44.210 ;
        RECT 47.080 42.830 47.220 47.755 ;
        RECT 51.220 45.890 51.360 69.030 ;
        RECT 51.680 64.930 51.820 69.370 ;
        RECT 51.620 64.610 51.880 64.930 ;
        RECT 51.620 63.590 51.880 63.910 ;
        RECT 51.680 61.530 51.820 63.590 ;
        RECT 51.620 61.210 51.880 61.530 ;
        RECT 51.680 58.810 51.820 61.210 ;
        RECT 51.620 58.490 51.880 58.810 ;
        RECT 51.160 45.570 51.420 45.890 ;
        RECT 48.860 44.550 49.120 44.870 ;
        RECT 49.320 44.550 49.580 44.870 ;
        RECT 47.480 44.210 47.740 44.530 ;
        RECT 48.400 44.210 48.660 44.530 ;
        RECT 47.020 42.685 47.280 42.830 ;
        RECT 43.340 42.170 43.600 42.490 ;
        RECT 47.010 42.315 47.290 42.685 ;
        RECT 47.020 41.830 47.280 42.150 ;
        RECT 39.580 40.615 41.460 40.985 ;
        RECT 47.080 39.770 47.220 41.830 ;
        RECT 38.280 39.450 38.540 39.770 ;
        RECT 47.020 39.450 47.280 39.770 ;
        RECT 35.520 38.770 35.780 39.090 ;
        RECT 38.340 37.050 38.480 39.450 ;
        RECT 39.200 38.430 39.460 38.750 ;
        RECT 39.660 38.430 39.920 38.750 ;
        RECT 39.260 37.730 39.400 38.430 ;
        RECT 39.200 37.410 39.460 37.730 ;
        RECT 39.720 37.390 39.860 38.430 ;
        RECT 47.080 37.730 47.220 39.450 ;
        RECT 47.020 37.410 47.280 37.730 ;
        RECT 39.660 37.070 39.920 37.390 ;
        RECT 34.140 36.730 34.400 37.050 ;
        RECT 38.280 36.730 38.540 37.050 ;
        RECT 33.220 36.390 33.480 36.710 ;
        RECT 33.280 36.030 33.420 36.390 ;
        RECT 33.220 35.710 33.480 36.030 ;
        RECT 27.240 31.630 27.500 31.950 ;
        RECT 24.020 28.570 24.280 28.890 ;
        RECT 27.300 28.550 27.440 31.630 ;
        RECT 33.280 28.890 33.420 35.710 ;
        RECT 34.200 35.010 34.340 36.730 ;
        RECT 34.140 34.690 34.400 35.010 ;
        RECT 38.340 31.610 38.480 36.730 ;
        RECT 39.580 35.175 41.460 35.545 ;
        RECT 47.080 33.310 47.220 37.410 ;
        RECT 47.540 37.050 47.680 44.210 ;
        RECT 48.460 42.490 48.600 44.210 ;
        RECT 48.400 42.170 48.660 42.490 ;
        RECT 48.460 41.470 48.600 42.170 ;
        RECT 48.400 41.150 48.660 41.470 ;
        RECT 48.460 39.430 48.600 41.150 ;
        RECT 48.400 39.110 48.660 39.430 ;
        RECT 47.480 36.730 47.740 37.050 ;
        RECT 47.540 34.330 47.680 36.730 ;
        RECT 47.480 34.010 47.740 34.330 ;
        RECT 41.040 32.990 41.300 33.310 ;
        RECT 47.020 32.990 47.280 33.310 ;
        RECT 41.100 31.610 41.240 32.990 ;
        RECT 45.180 31.630 45.440 31.950 ;
        RECT 38.280 31.290 38.540 31.610 ;
        RECT 41.040 31.290 41.300 31.610 ;
        RECT 38.340 28.890 38.480 31.290 ;
        RECT 39.580 29.735 41.460 30.105 ;
        RECT 45.240 29.570 45.380 31.630 ;
        RECT 45.180 29.250 45.440 29.570 ;
        RECT 33.220 28.570 33.480 28.890 ;
        RECT 38.280 28.570 38.540 28.890 ;
        RECT 40.580 28.570 40.840 28.890 ;
        RECT 19.880 28.230 20.140 28.550 ;
        RECT 23.100 28.230 23.360 28.550 ;
        RECT 27.240 28.230 27.500 28.550 ;
        RECT 19.420 27.550 19.680 27.870 ;
        RECT 21.720 27.550 21.980 27.870 ;
        RECT 17.580 25.850 17.840 26.170 ;
        RECT 18.040 25.850 18.300 26.170 ;
        RECT 17.640 25.150 17.780 25.850 ;
        RECT 19.420 25.510 19.680 25.830 ;
        RECT 17.580 24.830 17.840 25.150 ;
        RECT 9.580 24.295 11.460 24.665 ;
        RECT 19.480 24.130 19.620 25.510 ;
        RECT 19.420 23.810 19.680 24.130 ;
        RECT 21.780 23.110 21.920 27.550 ;
        RECT 24.580 27.015 26.460 27.385 ;
        RECT 27.300 26.850 27.440 28.230 ;
        RECT 31.840 27.890 32.100 28.210 ;
        RECT 30.000 27.550 30.260 27.870 ;
        RECT 27.240 26.530 27.500 26.850 ;
        RECT 30.060 26.170 30.200 27.550 ;
        RECT 31.900 26.850 32.040 27.890 ;
        RECT 31.840 26.530 32.100 26.850 ;
        RECT 30.000 25.850 30.260 26.170 ;
        RECT 33.680 25.850 33.940 26.170 ;
        RECT 32.760 24.830 33.020 25.150 ;
        RECT 32.820 23.110 32.960 24.830 ;
        RECT 33.740 24.130 33.880 25.850 ;
        RECT 33.680 23.810 33.940 24.130 ;
        RECT 21.720 22.790 21.980 23.110 ;
        RECT 32.760 22.790 33.020 23.110 ;
        RECT 24.580 21.575 26.460 21.945 ;
        RECT 9.580 18.855 11.460 19.225 ;
        RECT 38.340 18.010 38.480 28.570 ;
        RECT 40.640 26.170 40.780 28.570 ;
        RECT 47.540 28.550 47.680 34.010 ;
        RECT 48.920 31.950 49.060 44.550 ;
        RECT 49.380 43.250 49.520 44.550 ;
        RECT 49.380 43.110 49.980 43.250 ;
        RECT 52.140 43.170 52.280 74.470 ;
        RECT 52.600 70.370 52.740 87.990 ;
        RECT 53.000 85.690 53.260 86.010 ;
        RECT 53.460 85.690 53.720 86.010 ;
        RECT 53.060 82.270 53.200 85.690 ;
        RECT 53.000 81.950 53.260 82.270 ;
        RECT 53.060 78.045 53.200 81.950 ;
        RECT 52.990 77.675 53.270 78.045 ;
        RECT 53.000 77.190 53.260 77.510 ;
        RECT 53.060 75.810 53.200 77.190 ;
        RECT 53.000 75.490 53.260 75.810 ;
        RECT 53.000 74.810 53.260 75.130 ;
        RECT 52.540 70.050 52.800 70.370 ;
        RECT 52.540 66.990 52.800 67.310 ;
        RECT 52.600 66.630 52.740 66.990 ;
        RECT 52.540 66.310 52.800 66.630 ;
        RECT 52.540 65.630 52.800 65.950 ;
        RECT 52.600 64.250 52.740 65.630 ;
        RECT 52.540 63.930 52.800 64.250 ;
        RECT 52.540 63.250 52.800 63.570 ;
        RECT 52.600 56.770 52.740 63.250 ;
        RECT 53.060 62.210 53.200 74.810 ;
        RECT 53.520 67.650 53.660 85.690 ;
        RECT 53.980 84.990 54.120 90.110 ;
        RECT 56.680 88.070 56.940 88.390 ;
        RECT 54.580 86.855 56.460 87.225 ;
        RECT 56.740 86.690 56.880 88.070 ;
        RECT 56.680 86.370 56.940 86.690 ;
        RECT 55.300 85.350 55.560 85.670 ;
        RECT 53.920 84.670 54.180 84.990 ;
        RECT 55.360 83.970 55.500 85.350 ;
        RECT 57.200 85.330 57.340 106.770 ;
        RECT 60.360 100.990 60.620 101.310 ;
        RECT 61.740 100.990 62.000 101.310 ;
        RECT 58.520 98.950 58.780 99.270 ;
        RECT 58.580 97.570 58.720 98.950 ;
        RECT 60.420 98.930 60.560 100.990 ;
        RECT 60.360 98.610 60.620 98.930 ;
        RECT 58.520 97.250 58.780 97.570 ;
        RECT 61.800 96.890 61.940 100.990 ;
        RECT 57.600 96.570 57.860 96.890 ;
        RECT 61.740 96.570 62.000 96.890 ;
        RECT 57.660 94.170 57.800 96.570 ;
        RECT 57.600 93.850 57.860 94.170 ;
        RECT 57.140 85.010 57.400 85.330 ;
        RECT 57.660 84.730 57.800 93.850 ;
        RECT 62.260 91.450 62.400 107.710 ;
        RECT 64.500 107.110 64.760 107.430 ;
        RECT 64.560 104.710 64.700 107.110 ;
        RECT 64.500 104.390 64.760 104.710 ;
        RECT 64.560 102.330 64.700 104.390 ;
        RECT 64.500 102.010 64.760 102.330 ;
        RECT 62.660 101.670 62.920 101.990 ;
        RECT 62.720 98.590 62.860 101.670 ;
        RECT 62.660 98.270 62.920 98.590 ;
        RECT 60.820 91.130 61.080 91.450 ;
        RECT 62.200 91.130 62.460 91.450 ;
        RECT 60.880 88.390 61.020 91.130 ;
        RECT 60.820 88.070 61.080 88.390 ;
        RECT 57.200 84.590 57.800 84.730 ;
        RECT 55.300 83.650 55.560 83.970 ;
        RECT 54.580 81.415 56.460 81.785 ;
        RECT 56.680 76.850 56.940 77.170 ;
        RECT 54.580 75.975 56.460 76.345 ;
        RECT 56.740 75.810 56.880 76.850 ;
        RECT 56.680 75.490 56.940 75.810 ;
        RECT 53.920 72.090 54.180 72.410 ;
        RECT 53.980 70.370 54.120 72.090 ;
        RECT 54.580 70.535 56.460 70.905 ;
        RECT 53.920 70.050 54.180 70.370 ;
        RECT 54.840 69.710 55.100 70.030 ;
        RECT 57.200 69.940 57.340 84.590 ;
        RECT 57.600 83.650 57.860 83.970 ;
        RECT 56.280 69.800 57.340 69.940 ;
        RECT 54.900 67.650 55.040 69.710 ;
        RECT 53.460 67.330 53.720 67.650 ;
        RECT 54.840 67.330 55.100 67.650 ;
        RECT 53.920 66.650 54.180 66.970 ;
        RECT 53.980 64.840 54.120 66.650 ;
        RECT 56.280 65.860 56.420 69.800 ;
        RECT 56.680 66.540 56.940 66.630 ;
        RECT 56.680 66.400 57.340 66.540 ;
        RECT 56.680 66.310 56.940 66.400 ;
        RECT 56.280 65.720 56.880 65.860 ;
        RECT 54.580 65.095 56.460 65.465 ;
        RECT 53.980 64.700 54.580 64.840 ;
        RECT 53.460 63.930 53.720 64.250 ;
        RECT 53.920 63.930 54.180 64.250 ;
        RECT 53.000 61.890 53.260 62.210 ;
        RECT 53.520 61.610 53.660 63.930 ;
        RECT 53.980 61.870 54.120 63.930 ;
        RECT 54.440 63.910 54.580 64.700 ;
        RECT 54.380 63.590 54.640 63.910 ;
        RECT 55.750 63.395 56.030 63.765 ;
        RECT 55.820 63.230 55.960 63.395 ;
        RECT 55.300 62.910 55.560 63.230 ;
        RECT 55.760 62.910 56.020 63.230 ;
        RECT 55.360 62.210 55.500 62.910 ;
        RECT 55.300 61.890 55.560 62.210 ;
        RECT 53.060 61.470 53.660 61.610 ;
        RECT 53.920 61.550 54.180 61.870 ;
        RECT 53.060 58.890 53.200 61.470 ;
        RECT 53.060 58.750 53.660 58.890 ;
        RECT 53.980 58.810 54.120 61.550 ;
        RECT 54.580 59.655 56.460 60.025 ;
        RECT 54.380 59.170 54.640 59.490 ;
        RECT 52.540 56.450 52.800 56.770 ;
        RECT 53.000 55.770 53.260 56.090 ;
        RECT 52.540 54.750 52.800 55.070 ;
        RECT 52.600 51.330 52.740 54.750 ;
        RECT 53.060 53.710 53.200 55.770 ;
        RECT 53.520 55.070 53.660 58.750 ;
        RECT 53.920 58.490 54.180 58.810 ;
        RECT 54.440 55.750 54.580 59.170 ;
        RECT 54.380 55.660 54.640 55.750 ;
        RECT 53.980 55.520 54.640 55.660 ;
        RECT 53.460 54.750 53.720 55.070 ;
        RECT 53.000 53.390 53.260 53.710 ;
        RECT 52.540 51.010 52.800 51.330 ;
        RECT 53.520 49.630 53.660 54.750 ;
        RECT 53.980 54.050 54.120 55.520 ;
        RECT 54.380 55.430 54.640 55.520 ;
        RECT 54.580 54.215 56.460 54.585 ;
        RECT 53.920 53.730 54.180 54.050 ;
        RECT 56.740 53.030 56.880 65.720 ;
        RECT 57.200 64.250 57.340 66.400 ;
        RECT 57.140 63.930 57.400 64.250 ;
        RECT 56.680 52.710 56.940 53.030 ;
        RECT 53.460 49.310 53.720 49.630 ;
        RECT 54.580 48.775 56.460 49.145 ;
        RECT 54.380 47.950 54.640 48.270 ;
        RECT 53.460 47.270 53.720 47.590 ;
        RECT 49.840 42.490 49.980 43.110 ;
        RECT 52.080 42.850 52.340 43.170 ;
        RECT 50.700 42.510 50.960 42.830 ;
        RECT 49.320 42.170 49.580 42.490 ;
        RECT 49.780 42.170 50.040 42.490 ;
        RECT 49.380 33.990 49.520 42.170 ;
        RECT 49.840 41.810 49.980 42.170 ;
        RECT 49.780 41.490 50.040 41.810 ;
        RECT 49.840 39.340 49.980 41.490 ;
        RECT 50.760 39.430 50.900 42.510 ;
        RECT 53.520 42.490 53.660 47.270 ;
        RECT 54.440 45.210 54.580 47.950 ;
        RECT 56.680 46.590 56.940 46.910 ;
        RECT 56.740 45.550 56.880 46.590 ;
        RECT 56.680 45.405 56.940 45.550 ;
        RECT 54.380 44.890 54.640 45.210 ;
        RECT 56.670 45.035 56.950 45.405 ;
        RECT 53.920 44.550 54.180 44.870 ;
        RECT 53.980 42.490 54.120 44.550 ;
        RECT 56.680 43.870 56.940 44.190 ;
        RECT 54.580 43.335 56.460 43.705 ;
        RECT 52.080 42.170 52.340 42.490 ;
        RECT 53.460 42.170 53.720 42.490 ;
        RECT 53.920 42.170 54.180 42.490 ;
        RECT 52.140 41.470 52.280 42.170 ;
        RECT 56.740 42.150 56.880 43.870 ;
        RECT 56.680 41.830 56.940 42.150 ;
        RECT 52.080 41.150 52.340 41.470 ;
        RECT 52.070 40.275 52.350 40.645 ;
        RECT 52.080 40.130 52.340 40.275 ;
        RECT 51.160 39.450 51.420 39.770 ;
        RECT 50.240 39.340 50.500 39.430 ;
        RECT 49.840 39.200 50.500 39.340 ;
        RECT 50.240 39.110 50.500 39.200 ;
        RECT 50.700 39.110 50.960 39.430 ;
        RECT 51.220 36.710 51.360 39.450 ;
        RECT 54.580 37.895 56.460 38.265 ;
        RECT 51.160 36.390 51.420 36.710 ;
        RECT 51.220 34.330 51.360 36.390 ;
        RECT 57.200 34.330 57.340 63.930 ;
        RECT 57.660 43.170 57.800 83.650 ;
        RECT 60.880 82.610 61.020 88.070 ;
        RECT 59.900 82.290 60.160 82.610 ;
        RECT 60.820 82.290 61.080 82.610 ;
        RECT 58.060 77.870 58.320 78.190 ;
        RECT 58.120 75.130 58.260 77.870 ;
        RECT 59.440 77.530 59.700 77.850 ;
        RECT 58.060 74.810 58.320 75.130 ;
        RECT 58.060 72.090 58.320 72.410 ;
        RECT 58.970 72.235 59.250 72.605 ;
        RECT 58.120 67.650 58.260 72.090 ;
        RECT 58.520 71.750 58.780 72.070 ;
        RECT 58.580 68.670 58.720 71.750 ;
        RECT 58.520 68.350 58.780 68.670 ;
        RECT 58.060 67.330 58.320 67.650 ;
        RECT 58.580 67.050 58.720 68.350 ;
        RECT 58.120 66.910 58.720 67.050 ;
        RECT 58.120 63.910 58.260 66.910 ;
        RECT 58.520 66.310 58.780 66.630 ;
        RECT 58.580 64.250 58.720 66.310 ;
        RECT 58.520 63.930 58.780 64.250 ;
        RECT 58.060 63.590 58.320 63.910 ;
        RECT 58.060 60.530 58.320 60.850 ;
        RECT 58.120 59.490 58.260 60.530 ;
        RECT 58.060 59.170 58.320 59.490 ;
        RECT 58.060 54.750 58.320 55.070 ;
        RECT 58.120 50.650 58.260 54.750 ;
        RECT 58.580 52.350 58.720 63.930 ;
        RECT 59.040 63.570 59.180 72.235 ;
        RECT 59.500 72.070 59.640 77.530 ;
        RECT 59.960 74.530 60.100 82.290 ;
        RECT 61.740 77.870 62.000 78.190 ;
        RECT 61.800 76.830 61.940 77.870 ;
        RECT 60.820 76.510 61.080 76.830 ;
        RECT 61.740 76.510 62.000 76.830 ;
        RECT 60.880 75.130 61.020 76.510 ;
        RECT 60.820 74.810 61.080 75.130 ;
        RECT 59.960 74.390 61.020 74.530 ;
        RECT 61.280 74.470 61.540 74.790 ;
        RECT 59.900 72.430 60.160 72.750 ;
        RECT 59.440 71.750 59.700 72.070 ;
        RECT 59.960 70.280 60.100 72.430 ;
        RECT 60.350 72.235 60.630 72.605 ;
        RECT 60.420 72.070 60.560 72.235 ;
        RECT 60.360 71.750 60.620 72.070 ;
        RECT 59.960 70.140 60.560 70.280 ;
        RECT 59.900 69.370 60.160 69.690 ;
        RECT 59.960 67.310 60.100 69.370 ;
        RECT 60.420 69.010 60.560 70.140 ;
        RECT 60.880 69.770 61.020 74.390 ;
        RECT 61.340 70.370 61.480 74.470 ;
        RECT 61.280 70.050 61.540 70.370 ;
        RECT 60.880 69.630 61.480 69.770 ;
        RECT 60.360 68.690 60.620 69.010 ;
        RECT 59.430 66.795 59.710 67.165 ;
        RECT 59.900 66.990 60.160 67.310 ;
        RECT 60.820 66.990 61.080 67.310 ;
        RECT 59.500 66.630 59.640 66.795 ;
        RECT 59.440 66.310 59.700 66.630 ;
        RECT 59.960 64.250 60.100 66.990 ;
        RECT 60.360 66.650 60.620 66.970 ;
        RECT 59.900 63.930 60.160 64.250 ;
        RECT 58.980 63.250 59.240 63.570 ;
        RECT 59.960 62.170 60.100 63.930 ;
        RECT 59.040 62.030 60.100 62.170 ;
        RECT 59.040 55.070 59.180 62.030 ;
        RECT 59.440 60.870 59.700 61.190 ;
        RECT 59.500 58.810 59.640 60.870 ;
        RECT 59.440 58.490 59.700 58.810 ;
        RECT 58.980 54.750 59.240 55.070 ;
        RECT 58.980 53.390 59.240 53.710 ;
        RECT 58.520 52.030 58.780 52.350 ;
        RECT 59.040 51.330 59.180 53.390 ;
        RECT 58.980 51.010 59.240 51.330 ;
        RECT 58.060 50.330 58.320 50.650 ;
        RECT 58.520 50.330 58.780 50.650 ;
        RECT 58.120 47.930 58.260 50.330 ;
        RECT 58.060 47.610 58.320 47.930 ;
        RECT 58.120 44.190 58.260 47.610 ;
        RECT 58.060 43.870 58.320 44.190 ;
        RECT 57.600 42.850 57.860 43.170 ;
        RECT 58.060 42.850 58.320 43.170 ;
        RECT 57.600 39.450 57.860 39.770 ;
        RECT 57.660 35.010 57.800 39.450 ;
        RECT 58.120 39.430 58.260 42.850 ;
        RECT 58.580 42.490 58.720 50.330 ;
        RECT 58.980 50.220 59.240 50.310 ;
        RECT 59.500 50.220 59.640 58.490 ;
        RECT 59.900 55.430 60.160 55.750 ;
        RECT 59.960 50.310 60.100 55.430 ;
        RECT 60.420 50.650 60.560 66.650 ;
        RECT 60.880 62.210 61.020 66.990 ;
        RECT 60.820 61.890 61.080 62.210 ;
        RECT 61.340 61.610 61.480 69.630 ;
        RECT 61.800 69.090 61.940 76.510 ;
        RECT 62.260 71.130 62.400 91.130 ;
        RECT 62.720 87.450 62.860 98.270 ;
        RECT 64.560 91.450 64.700 102.010 ;
        RECT 67.720 101.670 67.980 101.990 ;
        RECT 67.780 100.290 67.920 101.670 ;
        RECT 67.720 99.970 67.980 100.290 ;
        RECT 67.260 96.230 67.520 96.550 ;
        RECT 65.420 95.550 65.680 95.870 ;
        RECT 64.500 91.130 64.760 91.450 ;
        RECT 63.120 90.110 63.380 90.430 ;
        RECT 63.180 88.050 63.320 90.110 ;
        RECT 63.120 87.730 63.380 88.050 ;
        RECT 62.720 87.310 63.320 87.450 ;
        RECT 63.580 87.390 63.840 87.710 ;
        RECT 62.660 86.370 62.920 86.690 ;
        RECT 62.720 77.510 62.860 86.370 ;
        RECT 63.180 86.350 63.320 87.310 ;
        RECT 63.640 86.690 63.780 87.390 ;
        RECT 63.580 86.370 63.840 86.690 ;
        RECT 63.120 86.030 63.380 86.350 ;
        RECT 64.040 86.030 64.300 86.350 ;
        RECT 62.660 77.190 62.920 77.510 ;
        RECT 63.180 72.070 63.320 86.030 ;
        RECT 63.580 85.350 63.840 85.670 ;
        RECT 63.640 83.290 63.780 85.350 ;
        RECT 63.580 82.970 63.840 83.290 ;
        RECT 63.640 75.810 63.780 82.970 ;
        RECT 64.100 77.850 64.240 86.030 ;
        RECT 64.040 77.530 64.300 77.850 ;
        RECT 63.580 75.490 63.840 75.810 ;
        RECT 64.100 74.790 64.240 77.530 ;
        RECT 64.560 76.830 64.700 91.130 ;
        RECT 65.480 91.110 65.620 95.550 ;
        RECT 67.320 94.850 67.460 96.230 ;
        RECT 67.260 94.530 67.520 94.850 ;
        RECT 65.420 90.790 65.680 91.110 ;
        RECT 65.480 89.410 65.620 90.790 ;
        RECT 65.420 89.090 65.680 89.410 ;
        RECT 65.880 87.390 66.140 87.710 ;
        RECT 65.940 86.010 66.080 87.390 ;
        RECT 65.880 85.690 66.140 86.010 ;
        RECT 67.260 82.630 67.520 82.950 ;
        RECT 64.960 77.190 65.220 77.510 ;
        RECT 66.340 77.190 66.600 77.510 ;
        RECT 64.500 76.510 64.760 76.830 ;
        RECT 64.040 74.470 64.300 74.790 ;
        RECT 64.100 73.090 64.240 74.470 ;
        RECT 64.040 72.770 64.300 73.090 ;
        RECT 63.580 72.430 63.840 72.750 ;
        RECT 62.660 71.925 62.920 72.070 ;
        RECT 62.650 71.555 62.930 71.925 ;
        RECT 63.120 71.750 63.380 72.070 ;
        RECT 62.260 70.990 63.320 71.130 ;
        RECT 62.200 70.050 62.460 70.370 ;
        RECT 62.260 69.690 62.400 70.050 ;
        RECT 62.200 69.370 62.460 69.690 ;
        RECT 62.660 69.600 62.920 69.690 ;
        RECT 63.180 69.600 63.320 70.990 ;
        RECT 63.640 70.370 63.780 72.430 ;
        RECT 64.030 72.235 64.310 72.605 ;
        RECT 64.100 72.070 64.240 72.235 ;
        RECT 65.020 72.070 65.160 77.190 ;
        RECT 66.400 72.410 66.540 77.190 ;
        RECT 66.800 74.130 67.060 74.450 ;
        RECT 66.340 72.090 66.600 72.410 ;
        RECT 66.860 72.070 67.000 74.130 ;
        RECT 64.040 71.750 64.300 72.070 ;
        RECT 64.960 71.925 65.220 72.070 ;
        RECT 64.950 71.555 65.230 71.925 ;
        RECT 66.800 71.750 67.060 72.070 ;
        RECT 64.500 71.070 64.760 71.390 ;
        RECT 63.580 70.050 63.840 70.370 ;
        RECT 62.660 69.460 63.320 69.600 ;
        RECT 62.660 69.370 62.920 69.460 ;
        RECT 61.800 68.950 62.860 69.090 ;
        RECT 62.200 63.250 62.460 63.570 ;
        RECT 60.880 61.470 61.480 61.610 ;
        RECT 60.360 50.330 60.620 50.650 ;
        RECT 58.980 50.080 59.640 50.220 ;
        RECT 58.980 49.990 59.240 50.080 ;
        RECT 59.900 49.990 60.160 50.310 ;
        RECT 58.520 42.170 58.780 42.490 ;
        RECT 58.060 39.110 58.320 39.430 ;
        RECT 58.520 39.110 58.780 39.430 ;
        RECT 58.580 37.050 58.720 39.110 ;
        RECT 58.520 36.730 58.780 37.050 ;
        RECT 57.600 34.690 57.860 35.010 ;
        RECT 51.160 34.010 51.420 34.330 ;
        RECT 57.140 34.010 57.400 34.330 ;
        RECT 49.320 33.670 49.580 33.990 ;
        RECT 49.380 32.290 49.520 33.670 ;
        RECT 49.320 31.970 49.580 32.290 ;
        RECT 48.860 31.630 49.120 31.950 ;
        RECT 48.920 31.010 49.060 31.630 ;
        RECT 51.220 31.270 51.360 34.010 ;
        RECT 54.580 32.455 56.460 32.825 ;
        RECT 57.660 31.610 57.800 34.690 ;
        RECT 58.580 34.670 58.720 36.730 ;
        RECT 58.520 34.350 58.780 34.670 ;
        RECT 58.580 31.610 58.720 34.350 ;
        RECT 52.540 31.290 52.800 31.610 ;
        RECT 57.600 31.290 57.860 31.610 ;
        RECT 58.520 31.290 58.780 31.610 ;
        RECT 48.460 30.870 49.060 31.010 ;
        RECT 51.160 30.950 51.420 31.270 ;
        RECT 48.460 29.570 48.600 30.870 ;
        RECT 48.860 30.270 49.120 30.590 ;
        RECT 48.400 29.250 48.660 29.570 ;
        RECT 41.960 28.230 42.220 28.550 ;
        RECT 47.480 28.230 47.740 28.550 ;
        RECT 42.020 26.850 42.160 28.230 ;
        RECT 41.960 26.530 42.220 26.850 ;
        RECT 48.920 26.170 49.060 30.270 ;
        RECT 49.320 27.890 49.580 28.210 ;
        RECT 49.380 26.850 49.520 27.890 ;
        RECT 49.320 26.530 49.580 26.850 ;
        RECT 40.580 25.850 40.840 26.170 ;
        RECT 48.860 25.850 49.120 26.170 ;
        RECT 39.580 24.295 41.460 24.665 ;
        RECT 52.600 23.110 52.740 31.290 ;
        RECT 57.600 30.610 57.860 30.930 ;
        RECT 53.000 30.270 53.260 30.590 ;
        RECT 53.060 28.210 53.200 30.270 ;
        RECT 57.660 28.210 57.800 30.610 ;
        RECT 53.000 27.890 53.260 28.210 ;
        RECT 57.600 27.890 57.860 28.210 ;
        RECT 54.580 27.015 56.460 27.385 ;
        RECT 57.660 26.170 57.800 27.890 ;
        RECT 55.760 25.850 56.020 26.170 ;
        RECT 57.600 25.850 57.860 26.170 ;
        RECT 46.560 22.790 46.820 23.110 ;
        RECT 52.540 22.790 52.800 23.110 ;
        RECT 39.580 18.855 41.460 19.225 ;
        RECT 38.280 17.690 38.540 18.010 ;
        RECT 46.100 17.690 46.360 18.010 ;
        RECT 24.580 16.135 26.460 16.505 ;
        RECT 46.160 15.290 46.300 17.690 ;
        RECT 46.620 17.670 46.760 22.790 ;
        RECT 55.820 22.770 55.960 25.850 ;
        RECT 56.680 25.510 56.940 25.830 ;
        RECT 56.220 23.470 56.480 23.790 ;
        RECT 56.280 23.110 56.420 23.470 ;
        RECT 56.220 22.790 56.480 23.110 ;
        RECT 55.760 22.450 56.020 22.770 ;
        RECT 54.580 21.575 56.460 21.945 ;
        RECT 56.740 21.070 56.880 25.510 ;
        RECT 57.660 23.110 57.800 25.850 ;
        RECT 58.580 24.130 58.720 31.290 ;
        RECT 59.040 25.150 59.180 49.990 ;
        RECT 59.440 44.550 59.700 44.870 ;
        RECT 59.500 42.490 59.640 44.550 ;
        RECT 59.440 42.170 59.700 42.490 ;
        RECT 59.500 31.950 59.640 42.170 ;
        RECT 59.960 40.450 60.100 49.990 ;
        RECT 60.880 47.160 61.020 61.470 ;
        RECT 61.740 60.870 62.000 61.190 ;
        RECT 61.800 55.750 61.940 60.870 ;
        RECT 62.260 59.150 62.400 63.250 ;
        RECT 62.200 58.830 62.460 59.150 ;
        RECT 61.740 55.430 62.000 55.750 ;
        RECT 61.740 52.030 62.000 52.350 ;
        RECT 60.420 47.020 61.020 47.160 ;
        RECT 59.900 40.130 60.160 40.450 ;
        RECT 59.900 39.110 60.160 39.430 ;
        RECT 59.960 37.050 60.100 39.110 ;
        RECT 60.420 37.730 60.560 47.020 ;
        RECT 61.280 45.570 61.540 45.890 ;
        RECT 60.820 43.870 61.080 44.190 ;
        RECT 60.880 41.470 61.020 43.870 ;
        RECT 61.340 43.170 61.480 45.570 ;
        RECT 61.280 42.850 61.540 43.170 ;
        RECT 61.280 41.830 61.540 42.150 ;
        RECT 60.820 41.150 61.080 41.470 ;
        RECT 61.340 40.450 61.480 41.830 ;
        RECT 61.280 40.130 61.540 40.450 ;
        RECT 60.880 39.770 61.480 39.850 ;
        RECT 60.880 39.710 61.540 39.770 ;
        RECT 60.360 37.410 60.620 37.730 ;
        RECT 60.880 37.050 61.020 39.710 ;
        RECT 61.280 39.450 61.540 39.710 ;
        RECT 61.800 39.170 61.940 52.030 ;
        RECT 62.720 50.990 62.860 68.950 ;
        RECT 63.180 66.970 63.320 69.460 ;
        RECT 63.120 66.650 63.380 66.970 ;
        RECT 64.040 65.630 64.300 65.950 ;
        RECT 64.100 56.770 64.240 65.630 ;
        RECT 64.560 63.230 64.700 71.070 ;
        RECT 64.500 62.910 64.760 63.230 ;
        RECT 64.500 61.210 64.760 61.530 ;
        RECT 64.560 58.470 64.700 61.210 ;
        RECT 64.500 58.150 64.760 58.470 ;
        RECT 64.040 56.450 64.300 56.770 ;
        RECT 64.560 53.710 64.700 58.150 ;
        RECT 64.500 53.390 64.760 53.710 ;
        RECT 63.580 53.050 63.840 53.370 ;
        RECT 62.660 50.670 62.920 50.990 ;
        RECT 62.720 48.270 62.860 50.670 ;
        RECT 63.640 50.310 63.780 53.050 ;
        RECT 63.580 49.990 63.840 50.310 ;
        RECT 65.020 48.610 65.160 71.555 ;
        RECT 66.860 69.690 67.000 71.750 ;
        RECT 66.800 69.370 67.060 69.690 ;
        RECT 67.320 66.630 67.460 82.630 ;
        RECT 67.720 77.190 67.980 77.510 ;
        RECT 67.780 72.070 67.920 77.190 ;
        RECT 67.720 71.750 67.980 72.070 ;
        RECT 67.720 69.030 67.980 69.350 ;
        RECT 68.240 69.260 68.380 107.790 ;
        RECT 69.620 107.770 69.760 109.830 ;
        RECT 69.560 107.450 69.820 107.770 ;
        RECT 69.580 105.895 71.460 106.265 ;
        RECT 69.560 104.730 69.820 105.050 ;
        RECT 69.100 103.710 69.360 104.030 ;
        RECT 69.160 99.270 69.300 103.710 ;
        RECT 69.620 101.310 69.760 104.730 ;
        RECT 72.320 103.710 72.580 104.030 ;
        RECT 69.560 100.990 69.820 101.310 ;
        RECT 71.860 100.990 72.120 101.310 ;
        RECT 69.580 100.455 71.460 100.825 ;
        RECT 69.100 98.950 69.360 99.270 ;
        RECT 69.100 96.910 69.360 97.230 ;
        RECT 69.160 92.130 69.300 96.910 ;
        RECT 69.580 95.015 71.460 95.385 ;
        RECT 70.480 93.510 70.740 93.830 ;
        RECT 70.540 92.130 70.680 93.510 ;
        RECT 69.100 91.810 69.360 92.130 ;
        RECT 70.480 91.810 70.740 92.130 ;
        RECT 69.100 91.130 69.360 91.450 ;
        RECT 69.160 82.950 69.300 91.130 ;
        RECT 71.920 91.110 72.060 100.990 ;
        RECT 72.380 96.550 72.520 103.710 ;
        RECT 73.300 101.990 73.440 110.170 ;
        RECT 73.760 107.770 73.900 110.850 ;
        RECT 76.060 108.450 76.200 113.230 ;
        RECT 80.660 110.490 80.800 128.280 ;
        RECT 81.520 115.270 81.780 115.590 ;
        RECT 81.580 113.210 81.720 115.270 ;
        RECT 84.580 114.055 86.460 114.425 ;
        RECT 86.640 113.890 86.780 128.280 ;
        RECT 87.040 114.590 87.300 114.910 ;
        RECT 90.720 114.590 90.980 114.910 ;
        RECT 86.580 113.570 86.840 113.890 ;
        RECT 87.100 113.550 87.240 114.590 ;
        RECT 87.040 113.230 87.300 113.550 ;
        RECT 81.520 112.890 81.780 113.210 ;
        RECT 81.060 111.870 81.320 112.190 ;
        RECT 80.600 110.170 80.860 110.490 ;
        RECT 81.120 110.150 81.260 111.870 ;
        RECT 81.580 111.170 81.720 112.890 ;
        RECT 84.740 112.550 85.000 112.870 ;
        RECT 84.800 111.170 84.940 112.550 ;
        RECT 81.520 110.850 81.780 111.170 ;
        RECT 84.740 110.850 85.000 111.170 ;
        RECT 81.060 109.830 81.320 110.150 ;
        RECT 83.360 109.830 83.620 110.150 ;
        RECT 76.920 109.490 77.180 109.810 ;
        RECT 76.980 108.450 77.120 109.490 ;
        RECT 77.380 109.150 77.640 109.470 ;
        RECT 76.000 108.130 76.260 108.450 ;
        RECT 76.920 108.130 77.180 108.450 ;
        RECT 76.460 107.790 76.720 108.110 ;
        RECT 73.700 107.450 73.960 107.770 ;
        RECT 75.540 104.390 75.800 104.710 ;
        RECT 73.700 103.710 73.960 104.030 ;
        RECT 75.080 103.710 75.340 104.030 ;
        RECT 73.760 103.010 73.900 103.710 ;
        RECT 73.700 102.690 73.960 103.010 ;
        RECT 73.240 101.670 73.500 101.990 ;
        RECT 73.300 99.270 73.440 101.670 ;
        RECT 73.760 101.310 73.900 102.690 ;
        RECT 75.140 102.670 75.280 103.710 ;
        RECT 75.080 102.350 75.340 102.670 ;
        RECT 75.600 102.330 75.740 104.390 ;
        RECT 75.540 102.010 75.800 102.330 ;
        RECT 73.700 100.990 73.960 101.310 ;
        RECT 73.240 98.950 73.500 99.270 ;
        RECT 73.300 97.570 73.440 98.950 ;
        RECT 73.240 97.250 73.500 97.570 ;
        RECT 72.320 96.230 72.580 96.550 ;
        RECT 72.380 92.130 72.520 96.230 ;
        RECT 72.770 96.035 73.050 96.405 ;
        RECT 72.840 93.830 72.980 96.035 ;
        RECT 72.780 93.510 73.040 93.830 ;
        RECT 72.320 91.810 72.580 92.130 ;
        RECT 72.320 91.130 72.580 91.450 ;
        RECT 71.860 90.790 72.120 91.110 ;
        RECT 69.580 89.575 71.460 89.945 ;
        RECT 72.380 88.050 72.520 91.130 ;
        RECT 73.760 91.110 73.900 100.990 ;
        RECT 75.080 96.800 75.340 96.890 ;
        RECT 74.680 96.660 75.340 96.800 ;
        RECT 74.680 91.450 74.820 96.660 ;
        RECT 75.080 96.570 75.340 96.660 ;
        RECT 76.000 95.890 76.260 96.210 ;
        RECT 74.620 91.130 74.880 91.450 ;
        RECT 73.240 90.790 73.500 91.110 ;
        RECT 73.700 90.790 73.960 91.110 ;
        RECT 72.320 87.730 72.580 88.050 ;
        RECT 72.380 86.350 72.520 87.730 ;
        RECT 71.860 86.030 72.120 86.350 ;
        RECT 72.320 86.030 72.580 86.350 ;
        RECT 69.580 84.135 71.460 84.505 ;
        RECT 71.920 83.970 72.060 86.030 ;
        RECT 73.300 85.670 73.440 90.790 ;
        RECT 74.680 88.390 74.820 91.130 ;
        RECT 76.060 90.770 76.200 95.890 ;
        RECT 76.000 90.450 76.260 90.770 ;
        RECT 73.700 88.070 73.960 88.390 ;
        RECT 74.620 88.070 74.880 88.390 ;
        RECT 75.540 88.300 75.800 88.390 ;
        RECT 76.060 88.300 76.200 90.450 ;
        RECT 75.540 88.160 76.200 88.300 ;
        RECT 75.540 88.070 75.800 88.160 ;
        RECT 73.760 86.690 73.900 88.070 ;
        RECT 73.700 86.370 73.960 86.690 ;
        RECT 73.240 85.350 73.500 85.670 ;
        RECT 72.780 84.670 73.040 84.990 ;
        RECT 71.860 83.650 72.120 83.970 ;
        RECT 72.840 83.630 72.980 84.670 ;
        RECT 72.780 83.310 73.040 83.630 ;
        RECT 69.100 82.630 69.360 82.950 ;
        RECT 71.400 82.630 71.660 82.950 ;
        RECT 72.320 82.630 72.580 82.950 ;
        RECT 71.460 80.910 71.600 82.630 ;
        RECT 72.380 81.250 72.520 82.630 ;
        RECT 72.320 80.930 72.580 81.250 ;
        RECT 71.400 80.590 71.660 80.910 ;
        RECT 69.580 78.695 71.460 79.065 ;
        RECT 69.100 76.510 69.360 76.830 ;
        RECT 69.160 75.470 69.300 76.510 ;
        RECT 69.100 75.150 69.360 75.470 ;
        RECT 71.400 74.810 71.660 75.130 ;
        RECT 73.700 74.810 73.960 75.130 ;
        RECT 71.460 74.450 71.600 74.810 ;
        RECT 71.400 74.130 71.660 74.450 ;
        RECT 72.320 74.130 72.580 74.450 ;
        RECT 71.860 73.790 72.120 74.110 ;
        RECT 69.580 73.255 71.460 73.625 ;
        RECT 71.920 72.070 72.060 73.790 ;
        RECT 72.380 73.090 72.520 74.130 ;
        RECT 72.320 72.770 72.580 73.090 ;
        RECT 72.780 72.770 73.040 73.090 ;
        RECT 71.860 71.750 72.120 72.070 ;
        RECT 72.320 71.980 72.580 72.070 ;
        RECT 72.840 71.980 72.980 72.770 ;
        RECT 73.760 72.070 73.900 74.810 ;
        RECT 74.160 73.790 74.420 74.110 ;
        RECT 74.220 72.070 74.360 73.790 ;
        RECT 74.680 73.090 74.820 88.070 ;
        RECT 75.600 86.690 75.740 88.070 ;
        RECT 75.540 86.370 75.800 86.690 ;
        RECT 75.600 86.205 75.740 86.370 ;
        RECT 75.530 85.835 75.810 86.205 ;
        RECT 76.520 78.530 76.660 107.790 ;
        RECT 76.920 98.950 77.180 99.270 ;
        RECT 76.980 97.570 77.120 98.950 ;
        RECT 76.920 97.250 77.180 97.570 ;
        RECT 76.980 93.150 77.120 97.250 ;
        RECT 76.920 92.830 77.180 93.150 ;
        RECT 76.980 83.290 77.120 92.830 ;
        RECT 77.440 87.710 77.580 109.150 ;
        RECT 79.220 107.450 79.480 107.770 ;
        RECT 77.840 96.970 78.100 97.230 ;
        RECT 77.840 96.910 78.500 96.970 ;
        RECT 78.760 96.910 79.020 97.230 ;
        RECT 77.900 96.830 78.500 96.910 ;
        RECT 77.840 91.130 78.100 91.450 ;
        RECT 77.900 89.410 78.040 91.130 ;
        RECT 78.360 91.110 78.500 96.830 ;
        RECT 78.300 90.790 78.560 91.110 ;
        RECT 77.840 89.090 78.100 89.410 ;
        RECT 78.360 88.730 78.500 90.790 ;
        RECT 78.820 89.490 78.960 96.910 ;
        RECT 79.280 92.130 79.420 107.450 ;
        RECT 79.680 102.010 79.940 102.330 ;
        RECT 79.740 97.570 79.880 102.010 ;
        RECT 80.600 100.990 80.860 101.310 ;
        RECT 80.660 99.610 80.800 100.990 ;
        RECT 80.600 99.290 80.860 99.610 ;
        RECT 79.680 97.250 79.940 97.570 ;
        RECT 82.900 96.910 83.160 97.230 ;
        RECT 80.600 96.570 80.860 96.890 ;
        RECT 79.220 91.810 79.480 92.130 ;
        RECT 80.140 90.790 80.400 91.110 ;
        RECT 80.200 90.285 80.340 90.790 ;
        RECT 80.130 89.915 80.410 90.285 ;
        RECT 78.820 89.350 79.420 89.490 ;
        RECT 80.660 89.410 80.800 96.570 ;
        RECT 82.960 93.830 83.100 96.910 ;
        RECT 82.900 93.510 83.160 93.830 ;
        RECT 81.060 92.830 81.320 93.150 ;
        RECT 82.900 92.830 83.160 93.150 ;
        RECT 81.120 90.430 81.260 92.830 ;
        RECT 81.980 91.130 82.240 91.450 ;
        RECT 81.060 90.110 81.320 90.430 ;
        RECT 82.040 90.285 82.180 91.130 ;
        RECT 81.970 89.915 82.250 90.285 ;
        RECT 78.300 88.410 78.560 88.730 ;
        RECT 78.760 88.410 79.020 88.730 ;
        RECT 77.840 87.730 78.100 88.050 ;
        RECT 77.380 87.390 77.640 87.710 ;
        RECT 77.900 86.690 78.040 87.730 ;
        RECT 78.360 86.690 78.500 88.410 ;
        RECT 77.840 86.370 78.100 86.690 ;
        RECT 78.300 86.370 78.560 86.690 ;
        RECT 77.380 85.690 77.640 86.010 ;
        RECT 77.440 83.970 77.580 85.690 ;
        RECT 77.840 85.350 78.100 85.670 ;
        RECT 77.380 83.650 77.640 83.970 ;
        RECT 76.920 82.970 77.180 83.290 ;
        RECT 76.460 78.210 76.720 78.530 ;
        RECT 76.000 74.470 76.260 74.790 ;
        RECT 74.620 72.770 74.880 73.090 ;
        RECT 76.060 72.750 76.200 74.470 ;
        RECT 76.000 72.430 76.260 72.750 ;
        RECT 76.980 72.410 77.120 82.970 ;
        RECT 77.440 81.250 77.580 83.650 ;
        RECT 77.380 80.930 77.640 81.250 ;
        RECT 77.380 80.250 77.640 80.570 ;
        RECT 77.440 75.470 77.580 80.250 ;
        RECT 77.900 80.230 78.040 85.350 ;
        RECT 77.840 79.910 78.100 80.230 ;
        RECT 77.840 76.510 78.100 76.830 ;
        RECT 77.380 75.150 77.640 75.470 ;
        RECT 77.900 72.410 78.040 76.510 ;
        RECT 78.360 75.130 78.500 86.370 ;
        RECT 78.820 83.485 78.960 88.410 ;
        RECT 79.280 88.050 79.420 89.350 ;
        RECT 80.600 89.090 80.860 89.410 ;
        RECT 82.960 89.070 83.100 92.830 ;
        RECT 83.420 89.410 83.560 109.830 ;
        RECT 90.780 109.810 90.920 114.590 ;
        RECT 86.580 109.490 86.840 109.810 ;
        RECT 87.040 109.490 87.300 109.810 ;
        RECT 90.720 109.490 90.980 109.810 ;
        RECT 84.580 108.615 86.460 108.985 ;
        RECT 84.580 103.175 86.460 103.545 ;
        RECT 86.640 102.330 86.780 109.490 ;
        RECT 87.100 108.450 87.240 109.490 ;
        RECT 92.100 109.380 92.360 109.470 ;
        RECT 92.620 109.380 92.760 128.280 ;
        RECT 97.620 115.270 97.880 115.590 ;
        RECT 97.160 114.590 97.420 114.910 ;
        RECT 97.220 113.550 97.360 114.590 ;
        RECT 97.160 113.230 97.420 113.550 ;
        RECT 93.940 112.550 94.200 112.870 ;
        RECT 94.000 111.170 94.140 112.550 ;
        RECT 97.680 112.190 97.820 115.270 ;
        RECT 98.600 112.610 98.740 128.280 ;
        RECT 99.580 116.775 101.460 117.145 ;
        RECT 104.520 115.610 104.780 115.930 ;
        RECT 100.840 114.930 101.100 115.250 ;
        RECT 100.900 113.890 101.040 114.930 ;
        RECT 100.840 113.570 101.100 113.890 ;
        RECT 104.580 113.210 104.720 115.610 ;
        RECT 102.680 112.890 102.940 113.210 ;
        RECT 104.520 112.890 104.780 113.210 ;
        RECT 98.600 112.530 99.200 112.610 ;
        RECT 98.600 112.470 99.260 112.530 ;
        RECT 99.000 112.210 99.260 112.470 ;
        RECT 97.620 111.870 97.880 112.190 ;
        RECT 93.940 110.850 94.200 111.170 ;
        RECT 97.680 110.490 97.820 111.870 ;
        RECT 99.580 111.335 101.460 111.705 ;
        RECT 102.740 111.170 102.880 112.890 ;
        RECT 104.060 111.870 104.320 112.190 ;
        RECT 99.460 110.850 99.720 111.170 ;
        RECT 102.680 110.850 102.940 111.170 ;
        RECT 97.620 110.170 97.880 110.490 ;
        RECT 92.100 109.240 92.760 109.380 ;
        RECT 92.100 109.150 92.360 109.240 ;
        RECT 87.040 108.130 87.300 108.450 ;
        RECT 97.680 107.770 97.820 110.170 ;
        RECT 99.000 109.490 99.260 109.810 ;
        RECT 98.080 109.150 98.340 109.470 ;
        RECT 87.960 107.450 88.220 107.770 ;
        RECT 95.780 107.450 96.040 107.770 ;
        RECT 97.620 107.450 97.880 107.770 ;
        RECT 83.820 102.010 84.080 102.330 ;
        RECT 86.580 102.010 86.840 102.330 ;
        RECT 83.880 97.570 84.020 102.010 ;
        RECT 84.580 97.735 86.460 98.105 ;
        RECT 83.820 97.250 84.080 97.570 ;
        RECT 86.640 97.230 86.780 102.010 ;
        RECT 87.500 100.990 87.760 101.310 ;
        RECT 87.040 99.290 87.300 99.610 ;
        RECT 86.580 96.910 86.840 97.230 ;
        RECT 85.660 96.290 85.920 96.550 ;
        RECT 87.100 96.290 87.240 99.290 ;
        RECT 87.560 98.930 87.700 100.990 ;
        RECT 87.500 98.610 87.760 98.930 ;
        RECT 85.660 96.230 87.240 96.290 ;
        RECT 85.720 96.150 87.240 96.230 ;
        RECT 85.720 94.170 85.860 96.150 ;
        RECT 85.660 93.850 85.920 94.170 ;
        RECT 87.040 93.510 87.300 93.830 ;
        RECT 86.580 92.830 86.840 93.150 ;
        RECT 84.580 92.295 86.460 92.665 ;
        RECT 83.820 90.790 84.080 91.110 ;
        RECT 83.360 89.090 83.620 89.410 ;
        RECT 82.900 88.750 83.160 89.070 ;
        RECT 81.520 88.410 81.780 88.730 ;
        RECT 80.140 88.070 80.400 88.390 ;
        RECT 79.220 87.730 79.480 88.050 ;
        RECT 79.220 86.370 79.480 86.690 ;
        RECT 79.280 86.010 79.420 86.370 ;
        RECT 79.220 85.690 79.480 86.010 ;
        RECT 78.750 83.115 79.030 83.485 ;
        RECT 79.680 82.290 79.940 82.610 ;
        RECT 79.740 81.250 79.880 82.290 ;
        RECT 79.680 80.930 79.940 81.250 ;
        RECT 79.220 77.530 79.480 77.850 ;
        RECT 78.760 77.190 79.020 77.510 ;
        RECT 78.820 75.810 78.960 77.190 ;
        RECT 78.760 75.490 79.020 75.810 ;
        RECT 78.300 74.810 78.560 75.130 ;
        RECT 76.920 72.090 77.180 72.410 ;
        RECT 77.840 72.090 78.100 72.410 ;
        RECT 72.320 71.840 72.980 71.980 ;
        RECT 72.320 71.750 72.580 71.840 ;
        RECT 73.700 71.750 73.960 72.070 ;
        RECT 74.160 71.750 74.420 72.070 ;
        RECT 70.480 71.070 70.740 71.390 ;
        RECT 70.540 70.030 70.680 71.070 ;
        RECT 72.380 70.370 72.520 71.750 ;
        RECT 73.760 70.370 73.900 71.750 ;
        RECT 77.380 71.640 77.640 71.730 ;
        RECT 78.360 71.640 78.500 74.810 ;
        RECT 79.280 71.810 79.420 77.530 ;
        RECT 79.680 77.190 79.940 77.510 ;
        RECT 77.380 71.500 78.500 71.640 ;
        RECT 77.380 71.410 77.640 71.500 ;
        RECT 72.320 70.050 72.580 70.370 ;
        RECT 73.700 70.050 73.960 70.370 ;
        RECT 70.480 69.710 70.740 70.030 ;
        RECT 72.780 69.710 73.040 70.030 ;
        RECT 69.100 69.260 69.360 69.350 ;
        RECT 68.240 69.120 69.360 69.260 ;
        RECT 69.100 69.030 69.360 69.120 ;
        RECT 67.260 66.310 67.520 66.630 ;
        RECT 66.340 63.930 66.600 64.250 ;
        RECT 66.400 62.210 66.540 63.930 ;
        RECT 66.340 61.890 66.600 62.210 ;
        RECT 65.420 58.830 65.680 59.150 ;
        RECT 65.480 56.770 65.620 58.830 ;
        RECT 65.420 56.450 65.680 56.770 ;
        RECT 67.320 56.090 67.460 66.310 ;
        RECT 67.780 57.790 67.920 69.030 ;
        RECT 69.580 67.815 71.460 68.185 ;
        RECT 72.840 67.650 72.980 69.710 ;
        RECT 77.840 69.370 78.100 69.690 ;
        RECT 72.780 67.330 73.040 67.650 ;
        RECT 68.170 66.795 68.450 67.165 ;
        RECT 68.180 66.650 68.440 66.795 ;
        RECT 77.900 64.930 78.040 69.370 ;
        RECT 77.840 64.610 78.100 64.930 ;
        RECT 68.640 64.270 68.900 64.590 ;
        RECT 77.380 64.270 77.640 64.590 ;
        RECT 68.700 59.490 68.840 64.270 ;
        RECT 71.400 64.160 71.660 64.250 ;
        RECT 71.400 64.020 72.060 64.160 ;
        RECT 71.400 63.930 71.660 64.020 ;
        RECT 69.580 62.375 71.460 62.745 ;
        RECT 71.920 62.170 72.060 64.020 ;
        RECT 72.320 63.930 72.580 64.250 ;
        RECT 71.460 62.030 72.060 62.170 ;
        RECT 69.560 60.870 69.820 61.190 ;
        RECT 69.100 60.190 69.360 60.510 ;
        RECT 68.640 59.170 68.900 59.490 ;
        RECT 69.160 57.790 69.300 60.190 ;
        RECT 69.620 59.490 69.760 60.870 ;
        RECT 71.460 60.850 71.600 62.030 ;
        RECT 72.380 61.530 72.520 63.930 ;
        RECT 76.000 63.590 76.260 63.910 ;
        RECT 76.060 61.870 76.200 63.590 ;
        RECT 76.000 61.550 76.260 61.870 ;
        RECT 72.320 61.210 72.580 61.530 ;
        RECT 76.060 61.190 76.200 61.550 ;
        RECT 77.440 61.190 77.580 64.270 ;
        RECT 78.360 63.230 78.500 71.500 ;
        RECT 78.820 71.670 79.420 71.810 ;
        RECT 78.300 62.910 78.560 63.230 ;
        RECT 76.000 60.870 76.260 61.190 ;
        RECT 76.920 60.870 77.180 61.190 ;
        RECT 77.380 60.870 77.640 61.190 ;
        RECT 71.400 60.530 71.660 60.850 ;
        RECT 71.460 59.490 71.600 60.530 ;
        RECT 71.860 60.190 72.120 60.510 ;
        RECT 69.560 59.170 69.820 59.490 ;
        RECT 71.400 59.170 71.660 59.490 ;
        RECT 67.720 57.470 67.980 57.790 ;
        RECT 68.640 57.470 68.900 57.790 ;
        RECT 69.100 57.470 69.360 57.790 ;
        RECT 68.700 56.090 68.840 57.470 ;
        RECT 69.580 56.935 71.460 57.305 ;
        RECT 67.260 55.770 67.520 56.090 ;
        RECT 68.640 55.770 68.900 56.090 ;
        RECT 65.880 55.430 66.140 55.750 ;
        RECT 66.340 55.430 66.600 55.750 ;
        RECT 65.940 53.030 66.080 55.430 ;
        RECT 66.400 53.710 66.540 55.430 ;
        RECT 71.920 55.410 72.060 60.190 ;
        RECT 73.700 58.830 73.960 59.150 ;
        RECT 72.380 56.090 72.980 56.170 ;
        RECT 72.320 56.030 72.980 56.090 ;
        RECT 72.320 55.770 72.580 56.030 ;
        RECT 71.860 55.090 72.120 55.410 ;
        RECT 66.340 53.390 66.600 53.710 ;
        RECT 68.180 53.050 68.440 53.370 ;
        RECT 65.880 52.710 66.140 53.030 ;
        RECT 68.240 50.310 68.380 53.050 ;
        RECT 72.840 52.350 72.980 56.030 ;
        RECT 73.760 55.070 73.900 58.830 ;
        RECT 76.980 58.810 77.120 60.870 ;
        RECT 76.920 58.490 77.180 58.810 ;
        RECT 74.620 58.150 74.880 58.470 ;
        RECT 74.680 56.090 74.820 58.150 ;
        RECT 74.620 55.770 74.880 56.090 ;
        RECT 74.620 55.090 74.880 55.410 ;
        RECT 73.700 54.750 73.960 55.070 ;
        RECT 73.760 53.030 73.900 54.750 ;
        RECT 74.680 54.050 74.820 55.090 ;
        RECT 74.620 53.730 74.880 54.050 ;
        RECT 77.380 53.390 77.640 53.710 ;
        RECT 73.700 52.710 73.960 53.030 ;
        RECT 72.320 52.030 72.580 52.350 ;
        RECT 72.780 52.030 73.040 52.350 ;
        RECT 69.580 51.495 71.460 51.865 ;
        RECT 68.180 49.990 68.440 50.310 ;
        RECT 68.640 49.650 68.900 49.970 ;
        RECT 68.700 48.610 68.840 49.650 ;
        RECT 64.960 48.290 65.220 48.610 ;
        RECT 68.640 48.290 68.900 48.610 ;
        RECT 62.660 47.950 62.920 48.270 ;
        RECT 64.500 47.950 64.760 48.270 ;
        RECT 63.120 47.270 63.380 47.590 ;
        RECT 63.180 45.890 63.320 47.270 ;
        RECT 63.120 45.570 63.380 45.890 ;
        RECT 62.660 44.890 62.920 45.210 ;
        RECT 62.720 41.810 62.860 44.890 ;
        RECT 62.660 41.490 62.920 41.810 ;
        RECT 61.340 39.030 61.940 39.170 ;
        RECT 62.200 39.110 62.460 39.430 ;
        RECT 59.900 36.730 60.160 37.050 ;
        RECT 60.820 36.730 61.080 37.050 ;
        RECT 59.960 33.650 60.100 36.730 ;
        RECT 60.360 34.690 60.620 35.010 ;
        RECT 59.900 33.330 60.160 33.650 ;
        RECT 60.420 33.310 60.560 34.690 ;
        RECT 60.360 32.990 60.620 33.310 ;
        RECT 59.440 31.630 59.700 31.950 ;
        RECT 59.440 28.570 59.700 28.890 ;
        RECT 59.500 26.850 59.640 28.570 ;
        RECT 60.420 28.210 60.560 32.990 ;
        RECT 60.880 28.970 61.020 36.730 ;
        RECT 61.340 29.570 61.480 39.030 ;
        RECT 62.260 36.370 62.400 39.110 ;
        RECT 62.200 36.050 62.460 36.370 ;
        RECT 62.260 34.410 62.400 36.050 ;
        RECT 62.720 35.010 62.860 41.490 ;
        RECT 64.560 39.430 64.700 47.950 ;
        RECT 69.100 47.610 69.360 47.930 ;
        RECT 69.160 44.190 69.300 47.610 ;
        RECT 69.580 46.055 71.460 46.425 ;
        RECT 64.960 43.870 65.220 44.190 ;
        RECT 69.100 43.870 69.360 44.190 ;
        RECT 65.020 43.170 65.160 43.870 ;
        RECT 64.960 42.850 65.220 43.170 ;
        RECT 66.340 42.510 66.600 42.830 ;
        RECT 66.400 40.450 66.540 42.510 ;
        RECT 69.160 42.150 69.300 43.870 ;
        RECT 71.860 42.170 72.120 42.490 ;
        RECT 69.100 41.830 69.360 42.150 ;
        RECT 66.340 40.130 66.600 40.450 ;
        RECT 64.500 39.110 64.760 39.430 ;
        RECT 63.120 38.770 63.380 39.090 ;
        RECT 62.660 34.690 62.920 35.010 ;
        RECT 61.800 34.270 62.400 34.410 ;
        RECT 61.800 33.990 61.940 34.270 ;
        RECT 61.740 33.670 62.000 33.990 ;
        RECT 61.800 31.610 61.940 33.670 ;
        RECT 62.200 33.330 62.460 33.650 ;
        RECT 61.740 31.290 62.000 31.610 ;
        RECT 61.280 29.250 61.540 29.570 ;
        RECT 61.800 29.230 61.940 31.290 ;
        RECT 62.260 31.270 62.400 33.330 ;
        RECT 63.180 32.290 63.320 38.770 ;
        RECT 69.160 36.710 69.300 41.830 ;
        RECT 69.580 40.615 71.460 40.985 ;
        RECT 71.920 40.450 72.060 42.170 ;
        RECT 71.860 40.130 72.120 40.450 ;
        RECT 72.380 39.430 72.520 52.030 ;
        RECT 72.840 47.930 72.980 52.030 ;
        RECT 77.440 51.330 77.580 53.390 ;
        RECT 77.380 51.010 77.640 51.330 ;
        RECT 78.820 48.270 78.960 71.670 ;
        RECT 79.220 71.070 79.480 71.390 ;
        RECT 79.280 70.030 79.420 71.070 ;
        RECT 79.220 69.710 79.480 70.030 ;
        RECT 79.740 62.210 79.880 77.190 ;
        RECT 79.680 61.890 79.940 62.210 ;
        RECT 80.200 61.530 80.340 88.070 ;
        RECT 80.600 86.030 80.860 86.350 ;
        RECT 80.660 75.040 80.800 86.030 ;
        RECT 81.580 83.485 81.720 88.410 ;
        RECT 83.360 88.070 83.620 88.390 ;
        RECT 82.900 87.390 83.160 87.710 ;
        RECT 82.440 85.690 82.700 86.010 ;
        RECT 81.510 83.115 81.790 83.485 ;
        RECT 81.060 76.850 81.320 77.170 ;
        RECT 81.120 75.810 81.260 76.850 ;
        RECT 81.060 75.490 81.320 75.810 ;
        RECT 82.500 75.130 82.640 85.690 ;
        RECT 81.060 75.040 81.320 75.130 ;
        RECT 80.660 74.900 81.320 75.040 ;
        RECT 80.660 74.110 80.800 74.900 ;
        RECT 81.060 74.810 81.320 74.900 ;
        RECT 81.520 74.810 81.780 75.130 ;
        RECT 82.440 74.810 82.700 75.130 ;
        RECT 80.600 73.790 80.860 74.110 ;
        RECT 81.580 73.090 81.720 74.810 ;
        RECT 81.060 72.770 81.320 73.090 ;
        RECT 81.520 72.770 81.780 73.090 ;
        RECT 81.120 72.490 81.260 72.770 ;
        RECT 82.500 72.490 82.640 74.810 ;
        RECT 81.120 72.350 82.640 72.490 ;
        RECT 81.980 69.030 82.240 69.350 ;
        RECT 81.060 63.930 81.320 64.250 ;
        RECT 80.140 61.210 80.400 61.530 ;
        RECT 81.120 61.190 81.260 63.930 ;
        RECT 81.060 60.870 81.320 61.190 ;
        RECT 81.120 59.150 81.260 60.870 ;
        RECT 81.060 58.830 81.320 59.150 ;
        RECT 79.220 58.490 79.480 58.810 ;
        RECT 79.280 56.770 79.420 58.490 ;
        RECT 80.600 57.470 80.860 57.790 ;
        RECT 79.220 56.450 79.480 56.770 ;
        RECT 80.660 55.750 80.800 57.470 ;
        RECT 80.600 55.430 80.860 55.750 ;
        RECT 79.680 54.750 79.940 55.070 ;
        RECT 79.740 53.710 79.880 54.750 ;
        RECT 79.680 53.390 79.940 53.710 ;
        RECT 78.760 47.950 79.020 48.270 ;
        RECT 72.780 47.610 73.040 47.930 ;
        RECT 75.540 47.610 75.800 47.930 ;
        RECT 76.000 47.610 76.260 47.930 ;
        RECT 77.380 47.610 77.640 47.930 ;
        RECT 75.600 45.210 75.740 47.610 ;
        RECT 75.540 44.890 75.800 45.210 ;
        RECT 72.780 44.725 73.040 44.870 ;
        RECT 72.770 44.355 73.050 44.725 ;
        RECT 72.840 42.685 72.980 44.355 ;
        RECT 72.770 42.315 73.050 42.685 ;
        RECT 76.060 42.490 76.200 47.610 ;
        RECT 77.440 45.550 77.580 47.610 ;
        RECT 81.060 47.270 81.320 47.590 ;
        RECT 77.380 45.230 77.640 45.550 ;
        RECT 77.440 44.870 77.580 45.230 ;
        RECT 77.380 44.550 77.640 44.870 ;
        RECT 77.440 42.830 77.580 44.550 ;
        RECT 81.120 44.530 81.260 47.270 ;
        RECT 82.040 45.890 82.180 69.030 ;
        RECT 82.960 68.670 83.100 87.390 ;
        RECT 82.900 68.350 83.160 68.670 ;
        RECT 82.900 66.310 83.160 66.630 ;
        RECT 82.960 61.870 83.100 66.310 ;
        RECT 83.420 64.930 83.560 88.070 ;
        RECT 83.880 78.530 84.020 90.790 ;
        RECT 85.200 90.450 85.460 90.770 ;
        RECT 85.260 88.390 85.400 90.450 ;
        RECT 86.640 89.410 86.780 92.830 ;
        RECT 87.100 91.450 87.240 93.510 ;
        RECT 87.040 91.130 87.300 91.450 ;
        RECT 86.580 89.090 86.840 89.410 ;
        RECT 87.100 88.390 87.240 91.130 ;
        RECT 88.020 89.410 88.160 107.450 ;
        RECT 89.800 100.990 90.060 101.310 ;
        RECT 89.340 98.270 89.600 98.590 ;
        RECT 89.400 97.570 89.540 98.270 ;
        RECT 89.340 97.250 89.600 97.570 ;
        RECT 88.420 96.910 88.680 97.230 ;
        RECT 88.480 91.450 88.620 96.910 ;
        RECT 88.880 96.800 89.140 96.890 ;
        RECT 89.400 96.800 89.540 97.250 ;
        RECT 89.860 96.890 90.000 100.990 ;
        RECT 95.320 99.630 95.580 99.950 ;
        RECT 93.480 98.270 93.740 98.590 ;
        RECT 93.540 96.890 93.680 98.270 ;
        RECT 88.880 96.660 89.540 96.800 ;
        RECT 88.880 96.570 89.140 96.660 ;
        RECT 89.800 96.570 90.060 96.890 ;
        RECT 93.480 96.570 93.740 96.890 ;
        RECT 89.860 94.170 90.000 96.570 ;
        RECT 95.380 96.550 95.520 99.630 ;
        RECT 94.400 96.230 94.660 96.550 ;
        RECT 95.320 96.230 95.580 96.550 ;
        RECT 89.800 93.850 90.060 94.170 ;
        RECT 88.420 91.130 88.680 91.450 ;
        RECT 87.960 89.090 88.220 89.410 ;
        RECT 89.860 89.070 90.000 93.850 ;
        RECT 91.180 93.510 91.440 93.830 ;
        RECT 90.260 92.830 90.520 93.150 ;
        RECT 90.320 91.450 90.460 92.830 ;
        RECT 90.260 91.130 90.520 91.450 ;
        RECT 91.240 89.410 91.380 93.510 ;
        RECT 94.460 91.110 94.600 96.230 ;
        RECT 95.380 94.510 95.520 96.230 ;
        RECT 95.320 94.190 95.580 94.510 ;
        RECT 95.320 91.470 95.580 91.790 ;
        RECT 94.400 90.790 94.660 91.110 ;
        RECT 91.180 89.090 91.440 89.410 ;
        RECT 89.800 88.750 90.060 89.070 ;
        RECT 94.460 88.730 94.600 90.790 ;
        RECT 95.380 89.410 95.520 91.470 ;
        RECT 95.320 89.090 95.580 89.410 ;
        RECT 88.420 88.640 88.680 88.730 ;
        RECT 88.420 88.500 89.080 88.640 ;
        RECT 88.420 88.410 88.680 88.500 ;
        RECT 85.200 88.070 85.460 88.390 ;
        RECT 86.580 88.070 86.840 88.390 ;
        RECT 87.040 88.070 87.300 88.390 ;
        RECT 84.580 86.855 86.460 87.225 ;
        RECT 84.580 81.415 86.460 81.785 ;
        RECT 84.280 80.250 84.540 80.570 ;
        RECT 83.820 78.210 84.080 78.530 ;
        RECT 84.340 76.740 84.480 80.250 ;
        RECT 83.880 76.600 84.480 76.740 ;
        RECT 83.880 75.130 84.020 76.600 ;
        RECT 84.580 75.975 86.460 76.345 ;
        RECT 83.820 74.810 84.080 75.130 ;
        RECT 86.120 74.810 86.380 75.130 ;
        RECT 83.820 73.790 84.080 74.110 ;
        RECT 83.880 71.730 84.020 73.790 ;
        RECT 83.820 71.410 84.080 71.730 ;
        RECT 86.180 71.390 86.320 74.810 ;
        RECT 86.120 71.070 86.380 71.390 ;
        RECT 84.580 70.535 86.460 70.905 ;
        RECT 86.120 69.710 86.380 70.030 ;
        RECT 86.180 66.630 86.320 69.710 ;
        RECT 86.640 67.650 86.780 88.070 ;
        RECT 87.960 76.510 88.220 76.830 ;
        RECT 87.500 74.810 87.760 75.130 ;
        RECT 87.040 74.470 87.300 74.790 ;
        RECT 86.580 67.330 86.840 67.650 ;
        RECT 86.120 66.540 86.380 66.630 ;
        RECT 85.720 66.400 86.380 66.540 ;
        RECT 83.820 65.970 84.080 66.290 ;
        RECT 83.360 64.610 83.620 64.930 ;
        RECT 83.880 62.210 84.020 65.970 ;
        RECT 85.720 65.950 85.860 66.400 ;
        RECT 86.120 66.310 86.380 66.400 ;
        RECT 85.660 65.630 85.920 65.950 ;
        RECT 84.580 65.095 86.460 65.465 ;
        RECT 85.660 63.930 85.920 64.250 ;
        RECT 86.580 63.930 86.840 64.250 ;
        RECT 83.820 61.890 84.080 62.210 ;
        RECT 82.900 61.550 83.160 61.870 ;
        RECT 83.350 61.355 83.630 61.725 ;
        RECT 83.360 61.210 83.620 61.355 ;
        RECT 82.440 60.870 82.700 61.190 ;
        RECT 83.820 60.870 84.080 61.190 ;
        RECT 82.500 55.750 82.640 60.870 ;
        RECT 83.360 60.530 83.620 60.850 ;
        RECT 82.900 58.490 83.160 58.810 ;
        RECT 82.440 55.430 82.700 55.750 ;
        RECT 82.960 47.250 83.100 58.490 ;
        RECT 83.420 58.380 83.560 60.530 ;
        RECT 83.880 59.150 84.020 60.870 ;
        RECT 85.720 60.510 85.860 63.930 ;
        RECT 86.640 61.870 86.780 63.930 ;
        RECT 86.580 61.550 86.840 61.870 ;
        RECT 86.120 61.100 86.380 61.190 ;
        RECT 86.120 60.960 86.780 61.100 ;
        RECT 86.120 60.870 86.380 60.960 ;
        RECT 85.660 60.190 85.920 60.510 ;
        RECT 84.580 59.655 86.460 60.025 ;
        RECT 83.820 58.830 84.080 59.150 ;
        RECT 84.740 58.720 85.000 58.810 ;
        RECT 84.340 58.580 85.000 58.720 ;
        RECT 84.340 58.380 84.480 58.580 ;
        RECT 84.740 58.490 85.000 58.580 ;
        RECT 83.420 58.240 84.480 58.380 ;
        RECT 86.640 55.750 86.780 60.960 ;
        RECT 87.100 59.490 87.240 74.470 ;
        RECT 87.040 59.170 87.300 59.490 ;
        RECT 86.580 55.430 86.840 55.750 ;
        RECT 86.580 54.750 86.840 55.070 ;
        RECT 84.580 54.215 86.460 54.585 ;
        RECT 86.640 53.030 86.780 54.750 ;
        RECT 83.360 52.710 83.620 53.030 ;
        RECT 86.580 52.710 86.840 53.030 ;
        RECT 83.420 47.590 83.560 52.710 ;
        RECT 87.560 51.330 87.700 74.810 ;
        RECT 88.020 74.110 88.160 76.510 ;
        RECT 87.960 73.790 88.220 74.110 ;
        RECT 87.960 54.750 88.220 55.070 ;
        RECT 87.500 51.010 87.760 51.330 ;
        RECT 87.040 50.670 87.300 50.990 ;
        RECT 86.580 49.990 86.840 50.310 ;
        RECT 83.820 49.650 84.080 49.970 ;
        RECT 83.360 47.270 83.620 47.590 ;
        RECT 82.900 46.930 83.160 47.250 ;
        RECT 81.980 45.570 82.240 45.890 ;
        RECT 81.520 44.890 81.780 45.210 ;
        RECT 81.060 44.210 81.320 44.530 ;
        RECT 81.120 42.830 81.260 44.210 ;
        RECT 77.380 42.510 77.640 42.830 ;
        RECT 81.060 42.510 81.320 42.830 ;
        RECT 76.000 42.170 76.260 42.490 ;
        RECT 79.680 42.400 79.940 42.490 ;
        RECT 79.680 42.260 80.340 42.400 ;
        RECT 79.680 42.170 79.940 42.260 ;
        RECT 73.700 41.830 73.960 42.150 ;
        RECT 73.240 41.150 73.500 41.470 ;
        RECT 73.300 40.110 73.440 41.150 ;
        RECT 73.240 39.790 73.500 40.110 ;
        RECT 72.320 39.110 72.580 39.430 ;
        RECT 70.480 38.430 70.740 38.750 ;
        RECT 70.540 37.390 70.680 38.430 ;
        RECT 70.480 37.070 70.740 37.390 ;
        RECT 72.380 36.710 72.520 39.110 ;
        RECT 73.760 39.090 73.900 41.830 ;
        RECT 74.160 41.150 74.420 41.470 ;
        RECT 74.220 39.770 74.360 41.150 ;
        RECT 74.160 39.450 74.420 39.770 ;
        RECT 75.080 39.450 75.340 39.770 ;
        RECT 73.700 38.770 73.960 39.090 ;
        RECT 69.100 36.390 69.360 36.710 ;
        RECT 72.320 36.390 72.580 36.710 ;
        RECT 64.040 33.670 64.300 33.990 ;
        RECT 63.120 31.970 63.380 32.290 ;
        RECT 64.100 31.270 64.240 33.670 ;
        RECT 62.200 30.950 62.460 31.270 ;
        RECT 64.040 30.950 64.300 31.270 ;
        RECT 69.160 30.930 69.300 36.390 ;
        RECT 69.580 35.175 71.460 35.545 ;
        RECT 71.400 31.970 71.660 32.290 ;
        RECT 71.460 31.010 71.600 31.970 ;
        RECT 69.100 30.610 69.360 30.930 ;
        RECT 71.460 30.870 72.060 31.010 ;
        RECT 68.640 30.270 68.900 30.590 ;
        RECT 60.880 28.830 61.480 28.970 ;
        RECT 61.740 28.910 62.000 29.230 ;
        RECT 62.660 28.910 62.920 29.230 ;
        RECT 60.360 27.890 60.620 28.210 ;
        RECT 59.900 27.550 60.160 27.870 ;
        RECT 59.440 26.530 59.700 26.850 ;
        RECT 59.960 26.510 60.100 27.550 ;
        RECT 59.900 26.190 60.160 26.510 ;
        RECT 58.980 24.830 59.240 25.150 ;
        RECT 58.060 23.810 58.320 24.130 ;
        RECT 58.520 23.810 58.780 24.130 ;
        RECT 57.600 22.790 57.860 23.110 ;
        RECT 57.140 22.450 57.400 22.770 ;
        RECT 56.680 20.750 56.940 21.070 ;
        RECT 52.080 20.410 52.340 20.730 ;
        RECT 49.320 19.390 49.580 19.710 ;
        RECT 49.380 18.010 49.520 19.390 ;
        RECT 52.140 18.690 52.280 20.410 ;
        RECT 53.460 19.390 53.720 19.710 ;
        RECT 52.080 18.370 52.340 18.690 ;
        RECT 49.320 17.690 49.580 18.010 ;
        RECT 46.560 17.350 46.820 17.670 ;
        RECT 46.100 14.970 46.360 15.290 ;
        RECT 46.620 14.270 46.760 17.350 ;
        RECT 52.540 17.010 52.800 17.330 ;
        RECT 47.020 16.670 47.280 16.990 ;
        RECT 47.080 15.630 47.220 16.670 ;
        RECT 52.600 15.970 52.740 17.010 ;
        RECT 52.540 15.650 52.800 15.970 ;
        RECT 47.020 15.310 47.280 15.630 ;
        RECT 53.520 14.950 53.660 19.390 ;
        RECT 54.580 16.135 56.460 16.505 ;
        RECT 56.740 14.950 56.880 20.750 ;
        RECT 57.200 20.730 57.340 22.450 ;
        RECT 57.140 20.410 57.400 20.730 ;
        RECT 58.120 18.690 58.260 23.810 ;
        RECT 58.580 21.410 58.720 23.810 ;
        RECT 59.960 23.790 60.100 26.190 ;
        RECT 61.340 24.130 61.480 28.830 ;
        RECT 61.740 27.890 62.000 28.210 ;
        RECT 61.800 26.930 61.940 27.890 ;
        RECT 61.800 26.850 62.400 26.930 ;
        RECT 61.800 26.790 62.460 26.850 ;
        RECT 61.280 23.810 61.540 24.130 ;
        RECT 59.900 23.470 60.160 23.790 ;
        RECT 59.960 22.850 60.100 23.470 ;
        RECT 59.500 22.710 60.100 22.850 ;
        RECT 58.980 22.110 59.240 22.430 ;
        RECT 58.520 21.090 58.780 21.410 ;
        RECT 59.040 21.070 59.180 22.110 ;
        RECT 58.980 20.750 59.240 21.070 ;
        RECT 58.980 20.070 59.240 20.390 ;
        RECT 58.520 19.390 58.780 19.710 ;
        RECT 58.060 18.370 58.320 18.690 ;
        RECT 58.580 17.330 58.720 19.390 ;
        RECT 59.040 17.330 59.180 20.070 ;
        RECT 59.500 18.690 59.640 22.710 ;
        RECT 59.900 22.110 60.160 22.430 ;
        RECT 60.360 22.110 60.620 22.430 ;
        RECT 59.960 20.390 60.100 22.110 ;
        RECT 60.420 20.730 60.560 22.110 ;
        RECT 61.340 21.070 61.480 23.810 ;
        RECT 61.800 23.110 61.940 26.790 ;
        RECT 62.200 26.530 62.460 26.790 ;
        RECT 62.200 25.850 62.460 26.170 ;
        RECT 61.740 22.790 62.000 23.110 ;
        RECT 62.260 21.410 62.400 25.850 ;
        RECT 62.720 22.770 62.860 28.910 ;
        RECT 68.700 28.550 68.840 30.270 ;
        RECT 69.160 28.550 69.300 30.610 ;
        RECT 69.580 29.735 71.460 30.105 ;
        RECT 68.640 28.230 68.900 28.550 ;
        RECT 69.100 28.230 69.360 28.550 ;
        RECT 65.880 22.790 66.140 23.110 ;
        RECT 62.660 22.450 62.920 22.770 ;
        RECT 62.200 21.090 62.460 21.410 ;
        RECT 61.280 20.750 61.540 21.070 ;
        RECT 62.720 20.810 62.860 22.450 ;
        RECT 63.120 22.110 63.380 22.430 ;
        RECT 60.360 20.410 60.620 20.730 ;
        RECT 62.260 20.670 62.860 20.810 ;
        RECT 59.900 20.070 60.160 20.390 ;
        RECT 59.440 18.370 59.700 18.690 ;
        RECT 58.520 17.010 58.780 17.330 ;
        RECT 58.980 17.010 59.240 17.330 ;
        RECT 58.580 15.630 58.720 17.010 ;
        RECT 58.520 15.310 58.780 15.630 ;
        RECT 53.460 14.630 53.720 14.950 ;
        RECT 56.680 14.630 56.940 14.950 ;
        RECT 59.960 14.270 60.100 20.070 ;
        RECT 62.260 20.050 62.400 20.670 ;
        RECT 62.200 19.730 62.460 20.050 ;
        RECT 60.820 17.010 61.080 17.330 ;
        RECT 60.880 15.970 61.020 17.010 ;
        RECT 60.820 15.650 61.080 15.970 ;
        RECT 63.180 15.630 63.320 22.110 ;
        RECT 65.940 21.410 66.080 22.790 ;
        RECT 65.880 21.090 66.140 21.410 ;
        RECT 64.500 20.070 64.760 20.390 ;
        RECT 64.560 19.710 64.700 20.070 ;
        RECT 64.500 19.390 64.760 19.710 ;
        RECT 64.560 18.010 64.700 19.390 ;
        RECT 65.940 18.010 66.080 21.090 ;
        RECT 67.260 20.750 67.520 21.070 ;
        RECT 67.320 20.390 67.460 20.750 ;
        RECT 67.260 20.070 67.520 20.390 ;
        RECT 69.160 19.710 69.300 28.230 ;
        RECT 69.580 24.295 71.460 24.665 ;
        RECT 69.100 19.390 69.360 19.710 ;
        RECT 69.580 18.855 71.460 19.225 ;
        RECT 64.500 17.690 64.760 18.010 ;
        RECT 65.880 17.690 66.140 18.010 ;
        RECT 71.920 17.670 72.060 30.870 ;
        RECT 72.380 26.170 72.520 36.390 ;
        RECT 75.140 34.330 75.280 39.450 ;
        RECT 72.780 34.010 73.040 34.330 ;
        RECT 75.080 34.010 75.340 34.330 ;
        RECT 72.840 31.270 72.980 34.010 ;
        RECT 76.060 32.290 76.200 42.170 ;
        RECT 78.290 41.635 78.570 42.005 ;
        RECT 78.360 41.470 78.500 41.635 ;
        RECT 78.760 41.490 79.020 41.810 ;
        RECT 78.300 41.150 78.560 41.470 ;
        RECT 78.820 39.430 78.960 41.490 ;
        RECT 80.200 39.430 80.340 42.260 ;
        RECT 81.120 39.770 81.260 42.510 ;
        RECT 81.580 42.490 81.720 44.890 ;
        RECT 81.520 42.170 81.780 42.490 ;
        RECT 82.960 41.470 83.100 46.930 ;
        RECT 83.360 45.570 83.620 45.890 ;
        RECT 83.420 44.870 83.560 45.570 ;
        RECT 83.880 44.870 84.020 49.650 ;
        RECT 84.580 48.775 86.460 49.145 ;
        RECT 86.120 47.270 86.380 47.590 ;
        RECT 86.180 46.910 86.320 47.270 ;
        RECT 86.120 46.590 86.380 46.910 ;
        RECT 85.200 45.570 85.460 45.890 ;
        RECT 85.650 45.715 85.930 46.085 ;
        RECT 85.660 45.570 85.920 45.715 ;
        RECT 83.360 44.550 83.620 44.870 ;
        RECT 83.820 44.550 84.080 44.870 ;
        RECT 85.260 44.780 85.400 45.570 ;
        RECT 86.640 45.210 86.780 49.990 ;
        RECT 86.580 44.890 86.840 45.210 ;
        RECT 85.660 44.780 85.920 44.870 ;
        RECT 85.260 44.640 85.920 44.780 ;
        RECT 85.660 44.550 85.920 44.640 ;
        RECT 86.580 44.210 86.840 44.530 ;
        RECT 83.360 43.870 83.620 44.190 ;
        RECT 83.420 42.490 83.560 43.870 ;
        RECT 84.580 43.335 86.460 43.705 ;
        RECT 83.360 42.170 83.620 42.490 ;
        RECT 84.740 41.830 85.000 42.150 ;
        RECT 82.900 41.150 83.160 41.470 ;
        RECT 81.510 40.275 81.790 40.645 ;
        RECT 84.800 40.450 84.940 41.830 ;
        RECT 81.520 40.130 81.780 40.275 ;
        RECT 84.740 40.130 85.000 40.450 ;
        RECT 86.120 39.790 86.380 40.110 ;
        RECT 81.060 39.450 81.320 39.770 ;
        RECT 86.180 39.430 86.320 39.790 ;
        RECT 78.760 39.110 79.020 39.430 ;
        RECT 80.140 39.110 80.400 39.430 ;
        RECT 86.120 39.110 86.380 39.430 ;
        RECT 77.840 38.430 78.100 38.750 ;
        RECT 82.900 38.430 83.160 38.750 ;
        RECT 77.900 37.730 78.040 38.430 ;
        RECT 77.840 37.410 78.100 37.730 ;
        RECT 77.900 33.990 78.040 37.410 ;
        RECT 80.600 36.390 80.860 36.710 ;
        RECT 80.660 33.990 80.800 36.390 ;
        RECT 77.840 33.670 78.100 33.990 ;
        RECT 80.600 33.900 80.860 33.990 ;
        RECT 80.600 33.760 81.260 33.900 ;
        RECT 80.600 33.670 80.860 33.760 ;
        RECT 80.140 32.990 80.400 33.310 ;
        RECT 80.600 32.990 80.860 33.310 ;
        RECT 76.000 31.970 76.260 32.290 ;
        RECT 79.220 31.970 79.480 32.290 ;
        RECT 76.460 31.860 76.720 31.950 ;
        RECT 76.460 31.720 77.120 31.860 ;
        RECT 76.460 31.630 76.720 31.720 ;
        RECT 76.980 31.270 77.120 31.720 ;
        RECT 72.780 30.950 73.040 31.270 ;
        RECT 75.080 30.950 75.340 31.270 ;
        RECT 76.920 30.950 77.180 31.270 ;
        RECT 78.300 30.950 78.560 31.270 ;
        RECT 72.840 30.590 72.980 30.950 ;
        RECT 72.780 30.270 73.040 30.590 ;
        RECT 75.140 29.570 75.280 30.950 ;
        RECT 75.080 29.250 75.340 29.570 ;
        RECT 76.920 27.890 77.180 28.210 ;
        RECT 76.980 26.850 77.120 27.890 ;
        RECT 76.920 26.530 77.180 26.850 ;
        RECT 72.320 25.850 72.580 26.170 ;
        RECT 78.360 24.130 78.500 30.950 ;
        RECT 79.280 29.230 79.420 31.970 ;
        RECT 79.220 28.910 79.480 29.230 ;
        RECT 80.200 28.550 80.340 32.990 ;
        RECT 80.660 31.610 80.800 32.990 ;
        RECT 80.600 31.290 80.860 31.610 ;
        RECT 81.120 28.550 81.260 33.760 ;
        RECT 82.960 33.650 83.100 38.430 ;
        RECT 84.580 37.895 86.460 38.265 ;
        RECT 82.900 33.330 83.160 33.650 ;
        RECT 82.960 32.290 83.100 33.330 ;
        RECT 84.580 32.455 86.460 32.825 ;
        RECT 82.900 31.970 83.160 32.290 ;
        RECT 86.640 31.950 86.780 44.210 ;
        RECT 87.100 37.050 87.240 50.670 ;
        RECT 88.020 48.270 88.160 54.750 ;
        RECT 87.960 47.950 88.220 48.270 ;
        RECT 87.500 46.590 87.760 46.910 ;
        RECT 87.560 42.150 87.700 46.590 ;
        RECT 88.940 45.890 89.080 88.500 ;
        RECT 94.400 88.410 94.660 88.730 ;
        RECT 90.260 84.670 90.520 84.990 ;
        RECT 93.940 84.670 94.200 84.990 ;
        RECT 89.800 80.250 90.060 80.570 ;
        RECT 89.860 78.530 90.000 80.250 ;
        RECT 89.800 78.210 90.060 78.530 ;
        RECT 90.320 77.510 90.460 84.670 ;
        RECT 94.000 82.950 94.140 84.670 ;
        RECT 94.860 82.970 95.120 83.290 ;
        RECT 93.940 82.630 94.200 82.950 ;
        RECT 93.020 80.930 93.280 81.250 ;
        RECT 90.260 77.190 90.520 77.510 ;
        RECT 90.320 72.070 90.460 77.190 ;
        RECT 91.640 76.510 91.900 76.830 ;
        RECT 91.700 74.110 91.840 76.510 ;
        RECT 93.080 75.810 93.220 80.930 ;
        RECT 93.940 77.870 94.200 78.190 ;
        RECT 93.020 75.490 93.280 75.810 ;
        RECT 94.000 75.470 94.140 77.870 ;
        RECT 93.940 75.150 94.200 75.470 ;
        RECT 93.480 74.810 93.740 75.130 ;
        RECT 92.100 74.470 92.360 74.790 ;
        RECT 91.640 73.790 91.900 74.110 ;
        RECT 90.260 71.750 90.520 72.070 ;
        RECT 90.720 69.370 90.980 69.690 ;
        RECT 91.640 69.370 91.900 69.690 ;
        RECT 90.780 68.670 90.920 69.370 ;
        RECT 90.720 68.350 90.980 68.670 ;
        RECT 90.780 66.630 90.920 68.350 ;
        RECT 91.700 67.310 91.840 69.370 ;
        RECT 91.640 67.220 91.900 67.310 ;
        RECT 91.240 67.080 91.900 67.220 ;
        RECT 90.720 66.310 90.980 66.630 ;
        RECT 91.240 66.290 91.380 67.080 ;
        RECT 91.640 66.990 91.900 67.080 ;
        RECT 91.640 66.310 91.900 66.630 ;
        RECT 91.180 65.970 91.440 66.290 ;
        RECT 91.700 65.950 91.840 66.310 ;
        RECT 91.640 65.630 91.900 65.950 ;
        RECT 89.800 63.140 90.060 63.230 ;
        RECT 89.800 63.000 90.460 63.140 ;
        RECT 89.800 62.910 90.060 63.000 ;
        RECT 90.320 62.210 90.460 63.000 ;
        RECT 90.260 61.890 90.520 62.210 ;
        RECT 91.180 54.750 91.440 55.070 ;
        RECT 91.240 54.050 91.380 54.750 ;
        RECT 91.180 53.730 91.440 54.050 ;
        RECT 90.720 50.330 90.980 50.650 ;
        RECT 88.880 45.570 89.140 45.890 ;
        RECT 89.330 45.035 89.610 45.405 ;
        RECT 87.960 44.550 88.220 44.870 ;
        RECT 87.500 41.830 87.760 42.150 ;
        RECT 87.040 36.730 87.300 37.050 ;
        RECT 86.580 31.630 86.840 31.950 ;
        RECT 87.560 31.270 87.700 41.830 ;
        RECT 88.020 38.750 88.160 44.550 ;
        RECT 88.420 41.150 88.680 41.470 ;
        RECT 88.480 39.430 88.620 41.150 ;
        RECT 89.400 39.430 89.540 45.035 ;
        RECT 89.800 42.510 90.060 42.830 ;
        RECT 88.420 39.110 88.680 39.430 ;
        RECT 88.880 39.110 89.140 39.430 ;
        RECT 89.340 39.110 89.600 39.430 ;
        RECT 87.960 38.430 88.220 38.750 ;
        RECT 88.480 37.050 88.620 39.110 ;
        RECT 88.420 36.730 88.680 37.050 ;
        RECT 88.940 33.990 89.080 39.110 ;
        RECT 89.400 36.370 89.540 39.110 ;
        RECT 89.860 37.730 90.000 42.510 ;
        RECT 89.800 37.410 90.060 37.730 ;
        RECT 89.800 36.390 90.060 36.710 ;
        RECT 89.340 36.050 89.600 36.370 ;
        RECT 89.860 35.010 90.000 36.390 ;
        RECT 89.800 34.690 90.060 35.010 ;
        RECT 88.880 33.670 89.140 33.990 ;
        RECT 88.940 32.290 89.080 33.670 ;
        RECT 89.340 32.990 89.600 33.310 ;
        RECT 88.880 31.970 89.140 32.290 ;
        RECT 87.500 31.010 87.760 31.270 ;
        RECT 87.100 30.950 87.760 31.010 ;
        RECT 87.100 30.870 87.700 30.950 ;
        RECT 84.280 30.270 84.540 30.590 ;
        RECT 84.340 28.550 84.480 30.270 ;
        RECT 87.100 28.890 87.240 30.870 ;
        RECT 87.960 30.270 88.220 30.590 ;
        RECT 88.020 28.890 88.160 30.270 ;
        RECT 88.940 29.570 89.080 31.970 ;
        RECT 89.400 31.610 89.540 32.990 ;
        RECT 89.860 31.610 90.000 34.690 ;
        RECT 90.780 33.650 90.920 50.330 ;
        RECT 91.170 45.035 91.450 45.405 ;
        RECT 91.240 44.870 91.380 45.035 ;
        RECT 91.180 44.550 91.440 44.870 ;
        RECT 91.640 44.550 91.900 44.870 ;
        RECT 91.180 43.870 91.440 44.190 ;
        RECT 91.240 43.170 91.380 43.870 ;
        RECT 91.180 42.850 91.440 43.170 ;
        RECT 91.240 39.430 91.380 42.850 ;
        RECT 91.700 41.380 91.840 44.550 ;
        RECT 92.160 43.170 92.300 74.470 ;
        RECT 93.540 70.370 93.680 74.810 ;
        RECT 93.940 74.130 94.200 74.450 ;
        RECT 93.480 70.050 93.740 70.370 ;
        RECT 92.560 69.370 92.820 69.690 ;
        RECT 92.620 66.630 92.760 69.370 ;
        RECT 92.560 66.310 92.820 66.630 ;
        RECT 93.020 63.590 93.280 63.910 ;
        RECT 93.080 61.530 93.220 63.590 ;
        RECT 94.000 62.170 94.140 74.130 ;
        RECT 94.920 74.110 95.060 82.970 ;
        RECT 95.840 75.810 95.980 107.450 ;
        RECT 97.160 104.390 97.420 104.710 ;
        RECT 97.620 104.390 97.880 104.710 ;
        RECT 96.700 103.710 96.960 104.030 ;
        RECT 96.760 102.670 96.900 103.710 ;
        RECT 97.220 103.010 97.360 104.390 ;
        RECT 97.160 102.690 97.420 103.010 ;
        RECT 96.700 102.350 96.960 102.670 ;
        RECT 96.240 102.010 96.500 102.330 ;
        RECT 96.300 97.085 96.440 102.010 ;
        RECT 96.230 96.715 96.510 97.085 ;
        RECT 96.700 90.110 96.960 90.430 ;
        RECT 96.760 88.390 96.900 90.110 ;
        RECT 96.700 88.070 96.960 88.390 ;
        RECT 97.160 88.070 97.420 88.390 ;
        RECT 96.760 82.690 96.900 88.070 ;
        RECT 97.220 83.630 97.360 88.070 ;
        RECT 97.160 83.310 97.420 83.630 ;
        RECT 96.760 82.550 97.360 82.690 ;
        RECT 96.700 81.950 96.960 82.270 ;
        RECT 96.760 80.910 96.900 81.950 ;
        RECT 96.700 80.590 96.960 80.910 ;
        RECT 97.220 77.850 97.360 82.550 ;
        RECT 97.680 81.250 97.820 104.390 ;
        RECT 98.140 99.690 98.280 109.150 ;
        RECT 99.060 108.450 99.200 109.490 ;
        RECT 99.000 108.130 99.260 108.450 ;
        RECT 99.520 107.170 99.660 110.850 ;
        RECT 104.120 109.810 104.260 111.870 ;
        RECT 104.060 109.490 104.320 109.810 ;
        RECT 98.540 106.770 98.800 107.090 ;
        RECT 99.060 107.030 99.660 107.170 ;
        RECT 98.600 105.730 98.740 106.770 ;
        RECT 98.540 105.410 98.800 105.730 ;
        RECT 98.140 99.550 98.740 99.690 ;
        RECT 98.080 98.950 98.340 99.270 ;
        RECT 98.140 97.570 98.280 98.950 ;
        RECT 98.080 97.250 98.340 97.570 ;
        RECT 98.140 94.170 98.280 97.250 ;
        RECT 98.080 93.850 98.340 94.170 ;
        RECT 98.140 91.450 98.280 93.850 ;
        RECT 98.080 91.130 98.340 91.450 ;
        RECT 98.140 83.290 98.280 91.130 ;
        RECT 98.080 82.970 98.340 83.290 ;
        RECT 97.620 80.930 97.880 81.250 ;
        RECT 98.140 80.230 98.280 82.970 ;
        RECT 98.080 79.910 98.340 80.230 ;
        RECT 97.620 79.230 97.880 79.550 ;
        RECT 97.160 77.530 97.420 77.850 ;
        RECT 97.680 76.830 97.820 79.230 ;
        RECT 98.140 77.510 98.280 79.910 ;
        RECT 98.080 77.190 98.340 77.510 ;
        RECT 97.620 76.510 97.880 76.830 ;
        RECT 95.780 75.490 96.040 75.810 ;
        RECT 95.320 74.810 95.580 75.130 ;
        RECT 96.700 74.810 96.960 75.130 ;
        RECT 94.400 73.790 94.660 74.110 ;
        RECT 94.860 73.790 95.120 74.110 ;
        RECT 94.460 73.090 94.600 73.790 ;
        RECT 94.400 72.770 94.660 73.090 ;
        RECT 94.400 71.070 94.660 71.390 ;
        RECT 94.460 69.010 94.600 71.070 ;
        RECT 94.400 68.690 94.660 69.010 ;
        RECT 94.460 66.630 94.600 68.690 ;
        RECT 95.380 67.650 95.520 74.810 ;
        RECT 96.760 72.750 96.900 74.810 ;
        RECT 97.160 74.470 97.420 74.790 ;
        RECT 96.700 72.430 96.960 72.750 ;
        RECT 96.240 69.370 96.500 69.690 ;
        RECT 95.780 68.350 96.040 68.670 ;
        RECT 95.320 67.330 95.580 67.650 ;
        RECT 95.840 66.630 95.980 68.350 ;
        RECT 94.400 66.310 94.660 66.630 ;
        RECT 95.780 66.310 96.040 66.630 ;
        RECT 96.300 65.950 96.440 69.370 ;
        RECT 96.700 66.310 96.960 66.630 ;
        RECT 95.320 65.630 95.580 65.950 ;
        RECT 96.240 65.630 96.500 65.950 ;
        RECT 95.380 64.590 95.520 65.630 ;
        RECT 95.320 64.270 95.580 64.590 ;
        RECT 96.760 62.210 96.900 66.310 ;
        RECT 93.540 62.030 94.140 62.170 ;
        RECT 93.020 61.210 93.280 61.530 ;
        RECT 92.560 60.190 92.820 60.510 ;
        RECT 92.620 55.070 92.760 60.190 ;
        RECT 92.560 54.750 92.820 55.070 ;
        RECT 92.560 53.050 92.820 53.370 ;
        RECT 92.620 50.990 92.760 53.050 ;
        RECT 92.560 50.670 92.820 50.990 ;
        RECT 92.100 42.850 92.360 43.170 ;
        RECT 92.100 41.380 92.360 41.470 ;
        RECT 91.700 41.240 92.360 41.380 ;
        RECT 92.100 41.150 92.360 41.240 ;
        RECT 92.160 39.430 92.300 41.150 ;
        RECT 92.560 39.450 92.820 39.770 ;
        RECT 91.180 39.110 91.440 39.430 ;
        RECT 92.100 39.110 92.360 39.430 ;
        RECT 91.240 38.490 91.380 39.110 ;
        RECT 91.240 38.350 92.300 38.490 ;
        RECT 92.160 37.050 92.300 38.350 ;
        RECT 92.100 36.730 92.360 37.050 ;
        RECT 92.620 36.710 92.760 39.450 ;
        RECT 93.540 37.730 93.680 62.030 ;
        RECT 96.700 61.890 96.960 62.210 ;
        RECT 96.700 61.210 96.960 61.530 ;
        RECT 96.760 56.770 96.900 61.210 ;
        RECT 96.700 56.450 96.960 56.770 ;
        RECT 97.220 56.170 97.360 74.470 ;
        RECT 97.680 72.410 97.820 76.510 ;
        RECT 98.600 75.470 98.740 99.550 ;
        RECT 99.060 75.810 99.200 107.030 ;
        RECT 99.580 105.895 101.460 106.265 ;
        RECT 104.580 104.710 104.720 112.890 ;
        RECT 105.960 110.490 106.100 128.790 ;
        RECT 107.280 114.930 107.540 115.250 ;
        RECT 107.340 113.890 107.480 114.930 ;
        RECT 107.280 113.570 107.540 113.890 ;
        RECT 105.900 110.170 106.160 110.490 ;
        RECT 110.560 108.450 110.700 128.280 ;
        RECT 116.540 116.610 116.680 128.280 ;
        RECT 116.480 116.290 116.740 116.610 ;
        RECT 110.500 108.130 110.760 108.450 ;
        RECT 104.980 107.790 105.240 108.110 ;
        RECT 105.040 105.730 105.180 107.790 ;
        RECT 104.980 105.410 105.240 105.730 ;
        RECT 104.520 104.390 104.780 104.710 ;
        RECT 102.220 102.350 102.480 102.670 ;
        RECT 99.580 100.455 101.460 100.825 ;
        RECT 99.920 98.610 100.180 98.930 ;
        RECT 99.980 97.570 100.120 98.610 ;
        RECT 99.920 97.250 100.180 97.570 ;
        RECT 102.280 96.890 102.420 102.350 ;
        RECT 106.360 102.010 106.620 102.330 ;
        RECT 102.680 100.990 102.940 101.310 ;
        RECT 104.520 100.990 104.780 101.310 ;
        RECT 102.740 99.270 102.880 100.990 ;
        RECT 104.580 99.610 104.720 100.990 ;
        RECT 104.060 99.290 104.320 99.610 ;
        RECT 104.520 99.290 104.780 99.610 ;
        RECT 102.680 98.950 102.940 99.270 ;
        RECT 102.220 96.570 102.480 96.890 ;
        RECT 99.580 95.015 101.460 95.385 ;
        RECT 102.280 94.850 102.420 96.570 ;
        RECT 104.120 96.290 104.260 99.290 ;
        RECT 106.420 97.570 106.560 102.010 ;
        RECT 107.280 100.990 107.540 101.310 ;
        RECT 107.340 98.930 107.480 100.990 ;
        RECT 107.280 98.610 107.540 98.930 ;
        RECT 106.360 97.250 106.620 97.570 ;
        RECT 104.520 96.290 104.780 96.550 ;
        RECT 104.120 96.230 104.780 96.290 ;
        RECT 104.980 96.230 105.240 96.550 ;
        RECT 104.120 96.150 104.720 96.230 ;
        RECT 102.220 94.530 102.480 94.850 ;
        RECT 99.580 89.575 101.460 89.945 ;
        RECT 102.280 88.390 102.420 94.530 ;
        RECT 104.580 88.730 104.720 96.150 ;
        RECT 105.040 94.170 105.180 96.230 ;
        RECT 104.980 93.850 105.240 94.170 ;
        RECT 105.040 92.130 105.180 93.850 ;
        RECT 110.500 93.510 110.760 93.830 ;
        RECT 106.360 92.830 106.620 93.150 ;
        RECT 104.980 91.810 105.240 92.130 ;
        RECT 104.520 88.410 104.780 88.730 ;
        RECT 102.220 88.070 102.480 88.390 ;
        RECT 103.600 87.390 103.860 87.710 ;
        RECT 99.580 84.135 101.460 84.505 ;
        RECT 103.660 83.970 103.800 87.390 ;
        RECT 103.600 83.650 103.860 83.970 ;
        RECT 103.600 80.250 103.860 80.570 ;
        RECT 101.760 79.910 102.020 80.230 ;
        RECT 99.580 78.695 101.460 79.065 ;
        RECT 101.820 78.530 101.960 79.910 ;
        RECT 102.680 79.230 102.940 79.550 ;
        RECT 101.760 78.210 102.020 78.530 ;
        RECT 102.740 77.850 102.880 79.230 ;
        RECT 103.660 77.850 103.800 80.250 ;
        RECT 104.580 78.530 104.720 88.410 ;
        RECT 105.040 88.390 105.180 91.810 ;
        RECT 106.420 89.070 106.560 92.830 ;
        RECT 110.560 91.450 110.700 93.510 ;
        RECT 110.040 91.130 110.300 91.450 ;
        RECT 110.500 91.130 110.760 91.450 ;
        RECT 108.660 90.110 108.920 90.430 ;
        RECT 106.360 88.750 106.620 89.070 ;
        RECT 104.980 88.070 105.240 88.390 ;
        RECT 108.720 88.050 108.860 90.110 ;
        RECT 110.100 89.410 110.240 91.130 ;
        RECT 110.040 89.090 110.300 89.410 ;
        RECT 108.660 87.730 108.920 88.050 ;
        RECT 105.900 83.650 106.160 83.970 ;
        RECT 104.520 78.210 104.780 78.530 ;
        RECT 102.680 77.530 102.940 77.850 ;
        RECT 103.600 77.530 103.860 77.850 ;
        RECT 103.660 75.810 103.800 77.530 ;
        RECT 99.000 75.490 99.260 75.810 ;
        RECT 103.600 75.490 103.860 75.810 ;
        RECT 98.540 75.150 98.800 75.470 ;
        RECT 98.080 74.810 98.340 75.130 ;
        RECT 97.620 72.090 97.880 72.410 ;
        RECT 98.140 67.650 98.280 74.810 ;
        RECT 104.580 74.790 104.720 78.210 ;
        RECT 105.960 75.810 106.100 83.650 ;
        RECT 106.360 82.970 106.620 83.290 ;
        RECT 106.420 81.250 106.560 82.970 ;
        RECT 106.360 80.930 106.620 81.250 ;
        RECT 110.560 80.570 110.700 91.130 ;
        RECT 110.960 82.290 111.220 82.610 ;
        RECT 111.020 81.250 111.160 82.290 ;
        RECT 110.960 80.930 111.220 81.250 ;
        RECT 107.280 80.250 107.540 80.570 ;
        RECT 110.500 80.250 110.760 80.570 ;
        RECT 107.340 75.810 107.480 80.250 ;
        RECT 107.740 79.230 108.000 79.550 ;
        RECT 107.800 77.170 107.940 79.230 ;
        RECT 107.740 76.850 108.000 77.170 ;
        RECT 105.900 75.490 106.160 75.810 ;
        RECT 107.280 75.490 107.540 75.810 ;
        RECT 104.520 74.470 104.780 74.790 ;
        RECT 99.580 73.255 101.460 73.625 ;
        RECT 99.000 69.370 99.260 69.690 ;
        RECT 104.520 69.370 104.780 69.690 ;
        RECT 98.540 69.030 98.800 69.350 ;
        RECT 97.620 67.330 97.880 67.650 ;
        RECT 98.080 67.330 98.340 67.650 ;
        RECT 97.680 66.630 97.820 67.330 ;
        RECT 97.620 66.310 97.880 66.630 ;
        RECT 98.600 64.590 98.740 69.030 ;
        RECT 99.060 66.370 99.200 69.370 ;
        RECT 101.760 68.350 102.020 68.670 ;
        RECT 104.060 68.350 104.320 68.670 ;
        RECT 99.580 67.815 101.460 68.185 ;
        RECT 101.820 66.970 101.960 68.350 ;
        RECT 101.760 66.650 102.020 66.970 ;
        RECT 99.060 66.230 99.660 66.370 ;
        RECT 99.920 66.310 100.180 66.630 ;
        RECT 99.000 64.610 99.260 64.930 ;
        RECT 98.540 64.270 98.800 64.590 ;
        RECT 97.620 61.890 97.880 62.210 ;
        RECT 97.680 58.130 97.820 61.890 ;
        RECT 99.060 61.190 99.200 64.610 ;
        RECT 99.520 63.570 99.660 66.230 ;
        RECT 99.980 64.930 100.120 66.310 ;
        RECT 103.140 65.630 103.400 65.950 ;
        RECT 99.920 64.610 100.180 64.930 ;
        RECT 103.200 64.590 103.340 65.630 ;
        RECT 103.140 64.270 103.400 64.590 ;
        RECT 99.460 63.250 99.720 63.570 ;
        RECT 102.220 63.250 102.480 63.570 ;
        RECT 99.580 62.375 101.460 62.745 ;
        RECT 102.280 61.870 102.420 63.250 ;
        RECT 102.220 61.550 102.480 61.870 ;
        RECT 99.000 60.870 99.260 61.190 ;
        RECT 97.620 57.810 97.880 58.130 ;
        RECT 96.760 56.030 97.360 56.170 ;
        RECT 94.400 54.750 94.660 55.070 ;
        RECT 94.460 47.330 94.600 54.750 ;
        RECT 94.860 52.030 95.120 52.350 ;
        RECT 94.920 48.270 95.060 52.030 ;
        RECT 94.860 47.950 95.120 48.270 ;
        RECT 94.860 47.330 95.120 47.590 ;
        RECT 94.460 47.270 95.120 47.330 ;
        RECT 94.460 47.190 95.060 47.270 ;
        RECT 94.390 45.035 94.670 45.405 ;
        RECT 94.460 42.490 94.600 45.035 ;
        RECT 96.240 44.725 96.500 44.870 ;
        RECT 96.230 44.355 96.510 44.725 ;
        RECT 94.400 42.170 94.660 42.490 ;
        RECT 94.860 42.170 95.120 42.490 ;
        RECT 95.780 42.170 96.040 42.490 ;
        RECT 94.920 39.770 95.060 42.170 ;
        RECT 95.840 41.810 95.980 42.170 ;
        RECT 95.780 41.490 96.040 41.810 ;
        RECT 96.760 40.450 96.900 56.030 ;
        RECT 97.160 55.430 97.420 55.750 ;
        RECT 97.220 51.330 97.360 55.430 ;
        RECT 97.160 51.010 97.420 51.330 ;
        RECT 97.680 49.970 97.820 57.810 ;
        RECT 98.540 57.470 98.800 57.790 ;
        RECT 98.600 55.750 98.740 57.470 ;
        RECT 99.060 55.750 99.200 60.870 ;
        RECT 102.280 58.810 102.420 61.550 ;
        RECT 104.120 61.530 104.260 68.350 ;
        RECT 104.580 64.930 104.720 69.370 ;
        RECT 109.580 68.690 109.840 69.010 ;
        RECT 105.440 68.350 105.700 68.670 ;
        RECT 105.500 66.290 105.640 68.350 ;
        RECT 105.900 67.330 106.160 67.650 ;
        RECT 105.440 65.970 105.700 66.290 ;
        RECT 105.960 64.930 106.100 67.330 ;
        RECT 109.640 66.630 109.780 68.690 ;
        RECT 109.580 66.310 109.840 66.630 ;
        RECT 104.520 64.610 104.780 64.930 ;
        RECT 105.900 64.610 106.160 64.930 ;
        RECT 105.960 62.210 106.100 64.610 ;
        RECT 105.900 61.890 106.160 62.210 ;
        RECT 104.060 61.210 104.320 61.530 ;
        RECT 105.960 59.490 106.100 61.890 ;
        RECT 105.900 59.170 106.160 59.490 ;
        RECT 109.640 58.810 109.780 66.310 ;
        RECT 110.040 65.630 110.300 65.950 ;
        RECT 110.100 60.850 110.240 65.630 ;
        RECT 110.040 60.530 110.300 60.850 ;
        RECT 102.220 58.490 102.480 58.810 ;
        RECT 109.580 58.490 109.840 58.810 ;
        RECT 99.580 56.935 101.460 57.305 ;
        RECT 98.540 55.430 98.800 55.750 ;
        RECT 99.000 55.430 99.260 55.750 ;
        RECT 98.080 54.750 98.340 55.070 ;
        RECT 98.140 53.370 98.280 54.750 ;
        RECT 98.080 53.050 98.340 53.370 ;
        RECT 99.060 53.030 99.200 55.430 ;
        RECT 99.000 52.710 99.260 53.030 ;
        RECT 97.620 49.650 97.880 49.970 ;
        RECT 99.060 47.930 99.200 52.710 ;
        RECT 99.580 51.495 101.460 51.865 ;
        RECT 102.280 50.650 102.420 58.490 ;
        RECT 103.140 58.150 103.400 58.470 ;
        RECT 103.200 56.770 103.340 58.150 ;
        RECT 105.440 57.470 105.700 57.790 ;
        RECT 103.140 56.450 103.400 56.770 ;
        RECT 102.680 52.030 102.940 52.350 ;
        RECT 102.220 50.330 102.480 50.650 ;
        RECT 102.740 49.970 102.880 52.030 ;
        RECT 103.200 50.310 103.340 56.450 ;
        RECT 105.500 55.410 105.640 57.470 ;
        RECT 109.640 55.750 109.780 58.490 ;
        RECT 109.580 55.430 109.840 55.750 ;
        RECT 105.440 55.090 105.700 55.410 ;
        RECT 110.040 54.750 110.300 55.070 ;
        RECT 110.100 53.710 110.240 54.750 ;
        RECT 110.040 53.390 110.300 53.710 ;
        RECT 103.140 49.990 103.400 50.310 ;
        RECT 102.680 49.650 102.940 49.970 ;
        RECT 99.000 47.610 99.260 47.930 ;
        RECT 99.060 45.890 99.200 47.610 ;
        RECT 99.580 46.055 101.460 46.425 ;
        RECT 99.000 45.570 99.260 45.890 ;
        RECT 102.680 45.570 102.940 45.890 ;
        RECT 97.620 41.830 97.880 42.150 ;
        RECT 96.700 40.130 96.960 40.450 ;
        RECT 94.860 39.450 95.120 39.770 ;
        RECT 93.940 38.430 94.200 38.750 ;
        RECT 93.480 37.410 93.740 37.730 ;
        RECT 94.000 37.050 94.140 38.430 ;
        RECT 94.920 37.050 95.060 39.450 ;
        RECT 96.700 38.430 96.960 38.750 ;
        RECT 96.760 37.390 96.900 38.430 ;
        RECT 97.680 37.730 97.820 41.830 ;
        RECT 99.580 40.615 101.460 40.985 ;
        RECT 102.220 39.680 102.480 39.770 ;
        RECT 102.740 39.680 102.880 45.570 ;
        RECT 103.140 41.490 103.400 41.810 ;
        RECT 102.220 39.540 102.880 39.680 ;
        RECT 102.220 39.450 102.480 39.540 ;
        RECT 102.680 38.770 102.940 39.090 ;
        RECT 97.620 37.410 97.880 37.730 ;
        RECT 102.740 37.390 102.880 38.770 ;
        RECT 96.700 37.070 96.960 37.390 ;
        RECT 102.680 37.070 102.940 37.390 ;
        RECT 93.940 36.730 94.200 37.050 ;
        RECT 94.860 36.730 95.120 37.050 ;
        RECT 92.560 36.450 92.820 36.710 ;
        RECT 91.700 36.390 92.820 36.450 ;
        RECT 91.700 36.310 92.760 36.390 ;
        RECT 91.700 34.330 91.840 36.310 ;
        RECT 91.640 34.010 91.900 34.330 ;
        RECT 95.320 34.010 95.580 34.330 ;
        RECT 90.720 33.330 90.980 33.650 ;
        RECT 89.340 31.290 89.600 31.610 ;
        RECT 89.800 31.290 90.060 31.610 ;
        RECT 91.700 30.930 91.840 34.010 ;
        RECT 93.480 32.990 93.740 33.310 ;
        RECT 93.540 31.950 93.680 32.990 ;
        RECT 95.380 32.290 95.520 34.010 ;
        RECT 96.760 33.990 96.900 37.070 ;
        RECT 103.200 37.050 103.340 41.490 ;
        RECT 104.060 38.770 104.320 39.090 ;
        RECT 104.120 37.730 104.260 38.770 ;
        RECT 104.060 37.410 104.320 37.730 ;
        RECT 102.220 36.730 102.480 37.050 ;
        RECT 103.140 36.730 103.400 37.050 ;
        RECT 99.580 35.175 101.460 35.545 ;
        RECT 102.280 35.010 102.420 36.730 ;
        RECT 102.220 34.690 102.480 35.010 ;
        RECT 96.700 33.670 96.960 33.990 ;
        RECT 95.320 31.970 95.580 32.290 ;
        RECT 93.480 31.630 93.740 31.950 ;
        RECT 102.280 31.610 102.420 34.690 ;
        RECT 102.220 31.290 102.480 31.610 ;
        RECT 91.640 30.610 91.900 30.930 ;
        RECT 90.720 30.270 90.980 30.590 ;
        RECT 88.880 29.250 89.140 29.570 ;
        RECT 87.040 28.570 87.300 28.890 ;
        RECT 87.960 28.570 88.220 28.890 ;
        RECT 80.140 28.230 80.400 28.550 ;
        RECT 81.060 28.230 81.320 28.550 ;
        RECT 84.280 28.230 84.540 28.550 ;
        RECT 81.980 27.550 82.240 27.870 ;
        RECT 83.360 27.550 83.620 27.870 ;
        RECT 78.300 23.810 78.560 24.130 ;
        RECT 82.040 22.770 82.180 27.550 ;
        RECT 83.420 23.450 83.560 27.550 ;
        RECT 84.580 27.015 86.460 27.385 ;
        RECT 87.100 23.450 87.240 28.570 ;
        RECT 90.780 28.210 90.920 30.270 ;
        RECT 99.580 29.735 101.460 30.105 ;
        RECT 90.720 27.890 90.980 28.210 ;
        RECT 99.580 24.295 101.460 24.665 ;
        RECT 83.360 23.130 83.620 23.450 ;
        RECT 87.040 23.130 87.300 23.450 ;
        RECT 81.980 22.450 82.240 22.770 ;
        RECT 84.580 21.575 86.460 21.945 ;
        RECT 72.320 20.410 72.580 20.730 ;
        RECT 72.380 18.690 72.520 20.410 ;
        RECT 99.580 18.855 101.460 19.225 ;
        RECT 72.320 18.370 72.580 18.690 ;
        RECT 71.860 17.350 72.120 17.670 ;
        RECT 84.580 16.135 86.460 16.505 ;
        RECT 63.120 15.310 63.380 15.630 ;
        RECT 46.560 13.950 46.820 14.270 ;
        RECT 59.900 13.950 60.160 14.270 ;
        RECT 9.580 13.415 11.460 13.785 ;
        RECT 39.580 13.415 41.460 13.785 ;
        RECT 69.580 13.415 71.460 13.785 ;
        RECT 99.580 13.415 101.460 13.785 ;
        RECT 24.580 10.695 26.460 11.065 ;
        RECT 54.580 10.695 56.460 11.065 ;
        RECT 84.580 10.695 86.460 11.065 ;
      LAYER met3 ;
        RECT 9.530 116.795 11.510 117.125 ;
        RECT 39.530 116.795 41.510 117.125 ;
        RECT 69.530 116.795 71.510 117.125 ;
        RECT 99.530 116.795 101.510 117.125 ;
        RECT 24.530 114.075 26.510 114.405 ;
        RECT 54.530 114.075 56.510 114.405 ;
        RECT 84.530 114.075 86.510 114.405 ;
        RECT 2.000 113.055 2.235 113.385 ;
        RECT 9.530 111.355 11.510 111.685 ;
        RECT 39.530 111.355 41.510 111.685 ;
        RECT 69.530 111.355 71.510 111.685 ;
        RECT 99.530 111.355 101.510 111.685 ;
        RECT 24.530 108.635 26.510 108.965 ;
        RECT 54.530 108.635 56.510 108.965 ;
        RECT 84.530 108.635 86.510 108.965 ;
        RECT 9.530 105.915 11.510 106.245 ;
        RECT 39.530 105.915 41.510 106.245 ;
        RECT 69.530 105.915 71.510 106.245 ;
        RECT 99.530 105.915 101.510 106.245 ;
        RECT 24.530 103.195 26.510 103.525 ;
        RECT 54.530 103.195 56.510 103.525 ;
        RECT 84.530 103.195 86.510 103.525 ;
        RECT 9.530 100.475 11.510 100.805 ;
        RECT 39.530 100.475 41.510 100.805 ;
        RECT 69.530 100.475 71.510 100.805 ;
        RECT 99.530 100.475 101.510 100.805 ;
        RECT 24.530 97.755 26.510 98.085 ;
        RECT 54.530 97.755 56.510 98.085 ;
        RECT 84.530 97.755 86.510 98.085 ;
        RECT 20.305 97.050 20.635 97.065 ;
        RECT 46.985 97.050 47.315 97.065 ;
        RECT 72.030 97.050 72.410 97.060 ;
        RECT 96.205 97.050 96.535 97.065 ;
        RECT 20.305 96.750 96.535 97.050 ;
        RECT 20.305 96.735 20.635 96.750 ;
        RECT 46.985 96.735 47.315 96.750 ;
        RECT 72.030 96.740 72.410 96.750 ;
        RECT 72.990 96.385 73.290 96.750 ;
        RECT 96.205 96.735 96.535 96.750 ;
        RECT 72.745 96.070 73.290 96.385 ;
        RECT 72.745 96.055 73.075 96.070 ;
        RECT 9.530 95.035 11.510 95.365 ;
        RECT 39.530 95.035 41.510 95.365 ;
        RECT 69.530 95.035 71.510 95.365 ;
        RECT 99.530 95.035 101.510 95.365 ;
        RECT 24.530 92.315 26.510 92.645 ;
        RECT 54.530 92.315 56.510 92.645 ;
        RECT 84.530 92.315 86.510 92.645 ;
        RECT 80.105 90.260 80.435 90.265 ;
        RECT 81.945 90.260 82.275 90.265 ;
        RECT 80.105 90.250 80.690 90.260 ;
        RECT 81.945 90.250 82.530 90.260 ;
        RECT 80.105 89.950 80.890 90.250 ;
        RECT 81.945 89.950 82.730 90.250 ;
        RECT 80.105 89.940 80.690 89.950 ;
        RECT 81.945 89.940 82.530 89.950 ;
        RECT 80.105 89.935 80.435 89.940 ;
        RECT 81.945 89.935 82.275 89.940 ;
        RECT 9.530 89.595 11.510 89.925 ;
        RECT 39.530 89.595 41.510 89.925 ;
        RECT 69.530 89.595 71.510 89.925 ;
        RECT 99.530 89.595 101.510 89.925 ;
        RECT 51.125 88.890 51.455 88.905 ;
        RECT 52.710 88.890 53.090 88.900 ;
        RECT 51.125 88.590 53.090 88.890 ;
        RECT 51.125 88.575 51.455 88.590 ;
        RECT 52.710 88.580 53.090 88.590 ;
        RECT 24.530 86.875 26.510 87.205 ;
        RECT 54.530 86.875 56.510 87.205 ;
        RECT 84.530 86.875 86.510 87.205 ;
        RECT 52.045 86.170 52.375 86.185 ;
        RECT 75.505 86.170 75.835 86.185 ;
        RECT 52.045 85.870 75.835 86.170 ;
        RECT 52.045 85.855 52.375 85.870 ;
        RECT 75.505 85.855 75.835 85.870 ;
        RECT 9.530 84.155 11.510 84.485 ;
        RECT 39.530 84.155 41.510 84.485 ;
        RECT 69.530 84.155 71.510 84.485 ;
        RECT 99.530 84.155 101.510 84.485 ;
        RECT 78.725 83.460 79.055 83.465 ;
        RECT 81.485 83.460 81.815 83.465 ;
        RECT 78.470 83.450 79.055 83.460 ;
        RECT 81.230 83.450 81.815 83.460 ;
        RECT 78.270 83.150 79.055 83.450 ;
        RECT 81.030 83.150 81.815 83.450 ;
        RECT 78.470 83.140 79.055 83.150 ;
        RECT 81.230 83.140 81.815 83.150 ;
        RECT 78.725 83.135 79.055 83.140 ;
        RECT 81.485 83.135 81.815 83.140 ;
        RECT 24.530 81.435 26.510 81.765 ;
        RECT 54.530 81.435 56.510 81.765 ;
        RECT 84.530 81.435 86.510 81.765 ;
        RECT 20.510 80.730 20.890 80.740 ;
        RECT 2.000 80.430 20.890 80.730 ;
        RECT 20.510 80.420 20.890 80.430 ;
        RECT 9.530 78.715 11.510 79.045 ;
        RECT 39.530 78.715 41.510 79.045 ;
        RECT 69.530 78.715 71.510 79.045 ;
        RECT 99.530 78.715 101.510 79.045 ;
        RECT 52.965 78.010 53.295 78.025 ;
        RECT 51.140 77.710 53.295 78.010 ;
        RECT 51.140 77.345 51.440 77.710 ;
        RECT 52.965 77.695 53.295 77.710 ;
        RECT 51.125 77.015 51.455 77.345 ;
        RECT 24.530 75.995 26.510 76.325 ;
        RECT 54.530 75.995 56.510 76.325 ;
        RECT 84.530 75.995 86.510 76.325 ;
        RECT 9.530 73.275 11.510 73.605 ;
        RECT 39.530 73.275 41.510 73.605 ;
        RECT 69.530 73.275 71.510 73.605 ;
        RECT 99.530 73.275 101.510 73.605 ;
        RECT 51.585 72.570 51.915 72.585 ;
        RECT 58.945 72.570 59.275 72.585 ;
        RECT 60.325 72.570 60.655 72.585 ;
        RECT 64.005 72.570 64.335 72.585 ;
        RECT 51.585 72.270 64.335 72.570 ;
        RECT 51.585 72.255 51.915 72.270 ;
        RECT 58.945 72.255 59.275 72.270 ;
        RECT 60.325 72.255 60.655 72.270 ;
        RECT 64.005 72.255 64.335 72.270 ;
        RECT 24.445 71.890 24.775 71.905 ;
        RECT 26.745 71.890 27.075 71.905 ;
        RECT 35.025 71.890 35.355 71.905 ;
        RECT 62.625 71.890 62.955 71.905 ;
        RECT 64.925 71.890 65.255 71.905 ;
        RECT 24.445 71.590 65.255 71.890 ;
        RECT 24.445 71.575 24.775 71.590 ;
        RECT 26.745 71.575 27.075 71.590 ;
        RECT 35.025 71.575 35.355 71.590 ;
        RECT 62.625 71.575 62.955 71.590 ;
        RECT 64.925 71.575 65.255 71.590 ;
        RECT 24.530 70.555 26.510 70.885 ;
        RECT 54.530 70.555 56.510 70.885 ;
        RECT 84.530 70.555 86.510 70.885 ;
        RECT 9.530 67.835 11.510 68.165 ;
        RECT 39.530 67.835 41.510 68.165 ;
        RECT 69.530 67.835 71.510 68.165 ;
        RECT 99.530 67.835 101.510 68.165 ;
        RECT 20.510 67.130 20.890 67.140 ;
        RECT 59.405 67.130 59.735 67.145 ;
        RECT 20.510 66.830 59.735 67.130 ;
        RECT 20.510 66.820 20.890 66.830 ;
        RECT 59.405 66.815 59.735 66.830 ;
        RECT 68.145 67.130 68.475 67.145 ;
        RECT 72.030 67.130 72.410 67.140 ;
        RECT 68.145 66.830 72.410 67.130 ;
        RECT 68.145 66.815 68.475 66.830 ;
        RECT 72.030 66.820 72.410 66.830 ;
        RECT 24.530 65.115 26.510 65.445 ;
        RECT 54.530 65.115 56.510 65.445 ;
        RECT 84.530 65.115 86.510 65.445 ;
        RECT 49.745 63.730 50.075 63.745 ;
        RECT 55.725 63.730 56.055 63.745 ;
        RECT 49.745 63.430 56.055 63.730 ;
        RECT 49.745 63.415 50.075 63.430 ;
        RECT 55.725 63.415 56.055 63.430 ;
        RECT 9.530 62.395 11.510 62.725 ;
        RECT 39.530 62.395 41.510 62.725 ;
        RECT 69.530 62.395 71.510 62.725 ;
        RECT 99.530 62.395 101.510 62.725 ;
        RECT 82.150 61.690 82.530 61.700 ;
        RECT 83.325 61.690 83.655 61.705 ;
        RECT 82.150 61.390 83.655 61.690 ;
        RECT 82.150 61.380 82.530 61.390 ;
        RECT 83.325 61.375 83.655 61.390 ;
        RECT 24.530 59.675 26.510 60.005 ;
        RECT 54.530 59.675 56.510 60.005 ;
        RECT 84.530 59.675 86.510 60.005 ;
        RECT 9.530 56.955 11.510 57.285 ;
        RECT 39.530 56.955 41.510 57.285 ;
        RECT 69.530 56.955 71.510 57.285 ;
        RECT 99.530 56.955 101.510 57.285 ;
        RECT 24.530 54.235 26.510 54.565 ;
        RECT 54.530 54.235 56.510 54.565 ;
        RECT 84.530 54.235 86.510 54.565 ;
        RECT 9.530 51.515 11.510 51.845 ;
        RECT 39.530 51.515 41.510 51.845 ;
        RECT 69.530 51.515 71.510 51.845 ;
        RECT 99.530 51.515 101.510 51.845 ;
        RECT 24.530 48.795 26.510 49.125 ;
        RECT 54.530 48.795 56.510 49.125 ;
        RECT 84.530 48.795 86.510 49.125 ;
        RECT 28.125 48.770 28.455 48.785 ;
        RECT 28.125 48.470 46.610 48.770 ;
        RECT 28.125 48.455 28.455 48.470 ;
        RECT 8.345 48.090 8.675 48.105 ;
        RECT 2.000 47.790 8.675 48.090 ;
        RECT 46.310 48.090 46.610 48.470 ;
        RECT 46.985 48.090 47.315 48.105 ;
        RECT 46.310 47.790 47.315 48.090 ;
        RECT 8.345 47.775 8.675 47.790 ;
        RECT 46.985 47.775 47.315 47.790 ;
        RECT 9.530 46.075 11.510 46.405 ;
        RECT 39.530 46.075 41.510 46.405 ;
        RECT 69.530 46.075 71.510 46.405 ;
        RECT 99.530 46.075 101.510 46.405 ;
        RECT 81.230 46.050 81.610 46.060 ;
        RECT 85.625 46.050 85.955 46.065 ;
        RECT 81.230 45.750 85.955 46.050 ;
        RECT 81.230 45.740 81.610 45.750 ;
        RECT 85.625 45.735 85.955 45.750 ;
        RECT 56.645 45.370 56.975 45.385 ;
        RECT 89.305 45.370 89.635 45.385 ;
        RECT 91.145 45.370 91.475 45.385 ;
        RECT 94.365 45.370 94.695 45.385 ;
        RECT 56.645 45.070 94.695 45.370 ;
        RECT 56.645 45.055 56.975 45.070 ;
        RECT 89.305 45.055 89.635 45.070 ;
        RECT 91.145 45.055 91.475 45.070 ;
        RECT 94.365 45.055 94.695 45.070 ;
        RECT 72.030 44.690 72.410 44.700 ;
        RECT 72.745 44.690 73.075 44.705 ;
        RECT 96.205 44.690 96.535 44.705 ;
        RECT 72.030 44.390 96.535 44.690 ;
        RECT 72.030 44.380 72.410 44.390 ;
        RECT 72.745 44.375 73.075 44.390 ;
        RECT 96.205 44.375 96.535 44.390 ;
        RECT 24.530 43.355 26.510 43.685 ;
        RECT 54.530 43.355 56.510 43.685 ;
        RECT 84.530 43.355 86.510 43.685 ;
        RECT 46.985 42.650 47.315 42.665 ;
        RECT 72.745 42.650 73.075 42.665 ;
        RECT 46.985 42.350 73.075 42.650 ;
        RECT 46.985 42.335 47.315 42.350 ;
        RECT 72.745 42.335 73.075 42.350 ;
        RECT 78.265 41.980 78.595 41.985 ;
        RECT 78.265 41.970 78.850 41.980 ;
        RECT 78.040 41.670 78.850 41.970 ;
        RECT 78.265 41.660 78.850 41.670 ;
        RECT 78.265 41.655 78.595 41.660 ;
        RECT 9.530 40.635 11.510 40.965 ;
        RECT 39.530 40.635 41.510 40.965 ;
        RECT 69.530 40.635 71.510 40.965 ;
        RECT 99.530 40.635 101.510 40.965 ;
        RECT 52.045 40.610 52.375 40.625 ;
        RECT 52.710 40.610 53.090 40.620 ;
        RECT 52.045 40.310 53.090 40.610 ;
        RECT 52.045 40.295 52.375 40.310 ;
        RECT 52.710 40.300 53.090 40.310 ;
        RECT 80.310 40.610 80.690 40.620 ;
        RECT 81.485 40.610 81.815 40.625 ;
        RECT 80.310 40.310 81.815 40.610 ;
        RECT 80.310 40.300 80.690 40.310 ;
        RECT 81.485 40.295 81.815 40.310 ;
        RECT 24.530 37.915 26.510 38.245 ;
        RECT 54.530 37.915 56.510 38.245 ;
        RECT 84.530 37.915 86.510 38.245 ;
        RECT 9.530 35.195 11.510 35.525 ;
        RECT 39.530 35.195 41.510 35.525 ;
        RECT 69.530 35.195 71.510 35.525 ;
        RECT 99.530 35.195 101.510 35.525 ;
        RECT 24.530 32.475 26.510 32.805 ;
        RECT 54.530 32.475 56.510 32.805 ;
        RECT 84.530 32.475 86.510 32.805 ;
        RECT 9.530 29.755 11.510 30.085 ;
        RECT 39.530 29.755 41.510 30.085 ;
        RECT 69.530 29.755 71.510 30.085 ;
        RECT 99.530 29.755 101.510 30.085 ;
        RECT 24.530 27.035 26.510 27.365 ;
        RECT 54.530 27.035 56.510 27.365 ;
        RECT 84.530 27.035 86.510 27.365 ;
        RECT 9.530 24.315 11.510 24.645 ;
        RECT 39.530 24.315 41.510 24.645 ;
        RECT 69.530 24.315 71.510 24.645 ;
        RECT 99.530 24.315 101.510 24.645 ;
        RECT 24.530 21.595 26.510 21.925 ;
        RECT 54.530 21.595 56.510 21.925 ;
        RECT 84.530 21.595 86.510 21.925 ;
        RECT 9.530 18.875 11.510 19.205 ;
        RECT 39.530 18.875 41.510 19.205 ;
        RECT 69.530 18.875 71.510 19.205 ;
        RECT 99.530 18.875 101.510 19.205 ;
        RECT 24.530 16.155 26.510 16.485 ;
        RECT 54.530 16.155 56.510 16.485 ;
        RECT 84.530 16.155 86.510 16.485 ;
        RECT 9.530 13.435 11.510 13.765 ;
        RECT 39.530 13.435 41.510 13.765 ;
        RECT 69.530 13.435 71.510 13.765 ;
        RECT 99.530 13.435 101.510 13.765 ;
        RECT 24.530 10.715 26.510 11.045 ;
        RECT 54.530 10.715 56.510 11.045 ;
        RECT 84.530 10.715 86.510 11.045 ;
      LAYER met4 ;
        RECT 72.055 96.735 72.385 97.065 ;
        RECT 52.735 88.575 53.065 88.905 ;
        RECT 20.535 80.415 20.865 80.745 ;
        RECT 20.550 67.145 20.850 80.415 ;
        RECT 20.535 66.815 20.865 67.145 ;
        RECT 52.750 40.625 53.050 88.575 ;
        RECT 72.070 67.145 72.370 96.735 ;
        RECT 80.335 89.935 80.665 90.265 ;
        RECT 82.175 89.935 82.505 90.265 ;
        RECT 78.495 83.135 78.825 83.465 ;
        RECT 72.055 66.815 72.385 67.145 ;
        RECT 72.070 44.705 72.370 66.815 ;
        RECT 72.055 44.375 72.385 44.705 ;
        RECT 78.510 41.985 78.810 83.135 ;
        RECT 78.495 41.655 78.825 41.985 ;
        RECT 80.350 40.625 80.650 89.935 ;
        RECT 81.255 83.135 81.585 83.465 ;
        RECT 81.270 46.065 81.570 83.135 ;
        RECT 82.190 61.705 82.490 89.935 ;
        RECT 82.175 61.375 82.505 61.705 ;
        RECT 81.255 45.735 81.585 46.065 ;
        RECT 52.735 40.295 53.065 40.625 ;
        RECT 80.335 40.295 80.665 40.625 ;
  END
END digital_top
END LIBRARY

