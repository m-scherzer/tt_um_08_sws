VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_08_sws
  CLASS BLOCK ;
  FOREIGN tt_um_08_sws ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER li1 ;
        RECT 75.440 155.565 75.755 156.125 ;
      LAYER met1 ;
        RECT 143.180 223.840 144.630 225.140 ;
        RECT 75.450 155.570 75.770 155.830 ;
        RECT 129.090 139.190 134.150 139.405 ;
        RECT 143.370 139.390 144.510 223.840 ;
        RECT 137.240 139.380 144.510 139.390 ;
        RECT 136.210 139.190 144.510 139.380 ;
        RECT 129.090 138.530 144.510 139.190 ;
        RECT 129.090 138.225 134.150 138.530 ;
        RECT 136.210 138.250 144.510 138.530 ;
        RECT 136.210 138.240 138.350 138.250 ;
      LAYER met2 ;
        RECT 143.230 223.790 144.580 225.190 ;
        RECT 75.480 155.540 75.740 155.860 ;
        RECT 75.540 154.015 75.680 155.540 ;
        RECT 75.470 153.645 75.750 154.015 ;
        RECT 129.140 138.175 134.100 139.455 ;
      LAYER met3 ;
        RECT 143.180 223.815 144.630 225.165 ;
        RECT 75.445 153.980 75.775 153.995 ;
        RECT 77.490 153.980 77.870 153.990 ;
        RECT 75.445 153.680 77.870 153.980 ;
        RECT 75.445 153.665 75.775 153.680 ;
        RECT 77.490 153.670 77.870 153.680 ;
        RECT 77.490 139.020 77.870 139.030 ;
        RECT 129.090 139.020 134.150 139.430 ;
        RECT 77.490 138.720 134.150 139.020 ;
        RECT 77.490 138.710 77.870 138.720 ;
        RECT 129.090 138.200 134.150 138.720 ;
      LAYER met4 ;
        RECT 143.830 225.145 144.130 225.760 ;
        RECT 143.225 223.835 144.585 225.145 ;
        RECT 77.515 153.665 77.845 153.995 ;
        RECT 77.530 139.035 77.830 153.665 ;
        RECT 77.515 138.705 77.845 139.035 ;
    END
  END clk
  PIN dem_dis
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 125.995 103.475 126.335 103.845 ;
      LAYER met1 ;
        RECT 135.340 223.880 136.790 225.180 ;
        RECT 135.635 174.550 136.775 223.880 ;
        RECT 135.580 173.430 136.830 174.550 ;
        RECT 135.635 173.420 136.775 173.430 ;
        RECT 135.580 165.470 136.830 166.590 ;
        RECT 135.635 141.220 136.775 165.470 ;
        RECT 135.580 140.230 136.830 141.220 ;
        RECT 135.635 140.155 136.775 140.230 ;
        RECT 135.660 134.480 136.800 134.510 ;
        RECT 135.590 133.400 136.850 134.480 ;
        RECT 135.660 106.690 136.800 133.400 ;
        RECT 133.100 106.600 136.850 106.690 ;
        RECT 129.700 105.630 136.850 106.600 ;
        RECT 133.100 105.500 136.850 105.630 ;
        RECT 126.065 103.750 126.355 103.795 ;
        RECT 126.510 103.750 126.830 103.810 ;
        RECT 126.065 103.610 126.830 103.750 ;
        RECT 126.065 103.565 126.355 103.610 ;
        RECT 126.510 103.550 126.830 103.610 ;
      LAYER met2 ;
        RECT 135.390 223.830 136.740 225.230 ;
        RECT 135.630 173.380 136.780 174.600 ;
        RECT 135.630 166.640 136.740 173.380 ;
        RECT 135.630 165.420 136.780 166.640 ;
        RECT 135.630 141.200 136.780 141.270 ;
        RECT 135.630 140.180 136.800 141.200 ;
        RECT 135.640 133.320 136.800 140.180 ;
        RECT 126.530 106.045 126.810 106.415 ;
        RECT 126.600 103.840 126.740 106.045 ;
        RECT 129.750 105.580 133.160 106.650 ;
        RECT 126.540 103.520 126.800 103.840 ;
      LAYER met3 ;
        RECT 135.340 223.855 136.790 225.205 ;
        RECT 129.700 106.530 133.210 106.625 ;
        RECT 126.505 106.380 126.835 106.395 ;
        RECT 129.340 106.380 133.340 106.530 ;
        RECT 126.505 106.080 133.340 106.380 ;
        RECT 126.505 106.065 126.835 106.080 ;
        RECT 129.340 105.930 133.340 106.080 ;
        RECT 129.700 105.605 133.210 105.930 ;
      LAYER met4 ;
        RECT 135.550 225.185 135.850 225.760 ;
        RECT 135.385 223.875 136.745 225.185 ;
    END
  END dem_dis
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN iop
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER li1 ;
        RECT 25.485 47.015 25.655 52.055 ;
        RECT 36.685 47.025 36.855 52.065 ;
        RECT 47.905 46.995 48.075 52.035 ;
        RECT 59.155 46.975 59.325 52.015 ;
        RECT 70.375 46.965 70.545 52.005 ;
        RECT 81.615 46.955 81.785 51.995 ;
        RECT 92.865 46.965 93.035 52.005 ;
        RECT 104.145 46.955 104.315 51.995 ;
        RECT 115.415 46.955 115.585 51.995 ;
        RECT 126.665 46.955 126.835 51.995 ;
        RECT 23.085 33.355 23.255 38.395 ;
        RECT 34.365 33.355 34.535 38.395 ;
        RECT 45.655 33.335 45.825 38.375 ;
        RECT 56.875 33.335 57.045 38.375 ;
        RECT 68.075 33.335 68.245 38.375 ;
        RECT 79.365 33.325 79.535 38.365 ;
        RECT 90.605 33.345 90.775 38.385 ;
        RECT 101.815 33.365 101.985 38.405 ;
        RECT 113.015 33.405 113.185 38.445 ;
        RECT 124.225 33.425 124.395 38.465 ;
      LAYER met1 ;
        RECT 25.455 51.980 25.685 52.035 ;
        RECT 36.655 51.990 36.885 52.045 ;
        RECT 25.305 47.010 25.735 51.980 ;
        RECT 36.505 47.020 36.935 51.990 ;
        RECT 47.875 51.960 48.105 52.015 ;
        RECT 47.725 46.990 48.155 51.960 ;
        RECT 59.125 51.940 59.355 51.995 ;
        RECT 58.975 46.970 59.405 51.940 ;
        RECT 70.345 51.930 70.575 51.985 ;
        RECT 70.195 46.960 70.625 51.930 ;
        RECT 81.585 51.920 81.815 51.975 ;
        RECT 92.835 51.930 93.065 51.985 ;
        RECT 81.435 46.950 81.865 51.920 ;
        RECT 92.685 46.960 93.115 51.930 ;
        RECT 104.115 51.920 104.345 51.975 ;
        RECT 115.385 51.920 115.615 51.975 ;
        RECT 126.635 51.920 126.865 51.975 ;
        RECT 103.965 46.950 104.395 51.920 ;
        RECT 115.235 46.950 115.665 51.920 ;
        RECT 126.485 46.950 126.915 51.920 ;
        RECT 29.055 45.020 41.225 45.030 ;
        RECT 17.855 45.005 41.225 45.020 ;
        RECT 15.900 45.000 41.225 45.005 ;
        RECT 15.900 44.980 52.445 45.000 ;
        RECT 15.900 44.970 63.695 44.980 ;
        RECT 15.900 44.960 74.915 44.970 ;
        RECT 85.235 44.960 97.405 44.970 ;
        RECT 15.900 43.880 131.205 44.960 ;
        RECT 15.900 43.870 30.025 43.880 ;
        RECT 15.900 43.855 18.690 43.870 ;
        RECT 15.900 41.620 17.050 43.855 ;
        RECT 40.275 43.850 131.205 43.880 ;
        RECT 51.525 43.830 131.205 43.850 ;
        RECT 62.745 43.820 131.205 43.830 ;
        RECT 73.985 43.810 86.155 43.820 ;
        RECT 96.515 43.810 131.205 43.820 ;
        RECT 15.900 41.540 19.685 41.620 ;
        RECT 141.160 41.610 146.210 41.640 ;
        RECT 119.855 41.590 146.210 41.610 ;
        RECT 108.645 41.550 146.210 41.590 ;
        RECT 15.900 41.520 42.165 41.540 ;
        RECT 97.445 41.530 146.210 41.550 ;
        RECT 15.900 41.510 75.875 41.520 ;
        RECT 86.235 41.510 146.210 41.530 ;
        RECT 15.900 40.500 146.210 41.510 ;
        RECT 15.900 40.470 142.250 40.500 ;
        RECT 18.715 40.460 142.250 40.470 ;
        RECT 18.715 40.440 120.815 40.460 ;
        RECT 18.715 40.400 109.615 40.440 ;
        RECT 18.715 40.390 98.405 40.400 ;
        RECT 41.285 40.380 98.405 40.390 ;
        RECT 41.285 40.370 87.165 40.380 ;
        RECT 74.995 40.360 87.165 40.370 ;
        RECT 23.005 33.430 23.435 38.400 ;
        RECT 34.285 33.430 34.715 38.400 ;
        RECT 23.055 33.375 23.285 33.430 ;
        RECT 34.335 33.375 34.565 33.430 ;
        RECT 45.575 33.410 46.005 38.380 ;
        RECT 56.795 33.410 57.225 38.380 ;
        RECT 67.995 33.410 68.425 38.380 ;
        RECT 45.625 33.355 45.855 33.410 ;
        RECT 56.845 33.355 57.075 33.410 ;
        RECT 68.045 33.355 68.275 33.410 ;
        RECT 79.285 33.400 79.715 38.370 ;
        RECT 90.525 33.420 90.955 38.390 ;
        RECT 101.735 33.440 102.165 38.410 ;
        RECT 112.935 33.480 113.365 38.450 ;
        RECT 124.145 33.500 124.575 38.470 ;
        RECT 79.335 33.345 79.565 33.400 ;
        RECT 90.575 33.365 90.805 33.420 ;
        RECT 101.785 33.385 102.015 33.440 ;
        RECT 112.985 33.425 113.215 33.480 ;
        RECT 124.195 33.445 124.425 33.500 ;
        RECT 145.070 18.880 146.210 40.500 ;
        RECT 145.030 17.960 146.250 18.880 ;
        RECT 145.020 14.870 146.160 14.980 ;
        RECT 144.980 13.950 146.200 14.870 ;
        RECT 145.020 6.630 146.160 13.950 ;
        RECT 93.650 5.490 146.160 6.630 ;
        RECT 93.650 1.480 94.790 5.490 ;
        RECT 93.500 0.230 94.890 1.480 ;
        RECT 93.650 0.150 94.790 0.230 ;
      LAYER met2 ;
        RECT 25.355 47.010 25.685 52.030 ;
        RECT 36.555 47.020 36.885 52.040 ;
        RECT 25.345 46.960 25.685 47.010 ;
        RECT 36.545 46.970 36.885 47.020 ;
        RECT 47.775 46.990 48.105 52.010 ;
        RECT 25.345 45.000 25.625 46.960 ;
        RECT 36.545 45.010 36.825 46.970 ;
        RECT 47.765 46.940 48.105 46.990 ;
        RECT 59.025 46.970 59.355 51.990 ;
        RECT 24.825 44.230 25.925 45.000 ;
        RECT 36.025 44.240 37.125 45.010 ;
        RECT 47.765 44.980 48.045 46.940 ;
        RECT 59.015 46.920 59.355 46.970 ;
        RECT 70.245 46.960 70.575 51.980 ;
        RECT 47.245 44.210 48.345 44.980 ;
        RECT 59.015 44.960 59.295 46.920 ;
        RECT 70.235 46.910 70.575 46.960 ;
        RECT 81.485 46.950 81.815 51.970 ;
        RECT 92.735 46.960 93.065 51.980 ;
        RECT 58.495 44.190 59.595 44.960 ;
        RECT 70.235 44.950 70.515 46.910 ;
        RECT 81.475 46.900 81.815 46.950 ;
        RECT 92.725 46.910 93.065 46.960 ;
        RECT 104.015 46.950 104.345 51.970 ;
        RECT 115.285 46.950 115.615 51.970 ;
        RECT 126.535 46.950 126.865 51.970 ;
        RECT 69.715 44.180 70.815 44.950 ;
        RECT 81.475 44.940 81.755 46.900 ;
        RECT 92.725 44.950 93.005 46.910 ;
        RECT 104.005 46.900 104.345 46.950 ;
        RECT 115.275 46.900 115.615 46.950 ;
        RECT 126.525 46.900 126.865 46.950 ;
        RECT 80.955 44.170 82.055 44.940 ;
        RECT 92.205 44.180 93.305 44.950 ;
        RECT 104.005 44.940 104.285 46.900 ;
        RECT 115.275 44.940 115.555 46.900 ;
        RECT 126.525 44.940 126.805 46.900 ;
        RECT 103.485 44.170 104.585 44.940 ;
        RECT 114.755 44.170 115.855 44.940 ;
        RECT 126.005 44.170 127.105 44.940 ;
        RECT 22.815 40.410 23.915 41.180 ;
        RECT 34.095 40.410 35.195 41.180 ;
        RECT 23.115 38.450 23.395 40.410 ;
        RECT 34.395 38.450 34.675 40.410 ;
        RECT 45.385 40.390 46.485 41.160 ;
        RECT 56.605 40.390 57.705 41.160 ;
        RECT 67.805 40.390 68.905 41.160 ;
        RECT 23.055 38.400 23.395 38.450 ;
        RECT 34.335 38.400 34.675 38.450 ;
        RECT 45.685 38.430 45.965 40.390 ;
        RECT 56.905 38.430 57.185 40.390 ;
        RECT 68.105 38.430 68.385 40.390 ;
        RECT 79.095 40.380 80.195 41.150 ;
        RECT 90.335 40.400 91.435 41.170 ;
        RECT 101.545 40.420 102.645 41.190 ;
        RECT 112.745 40.460 113.845 41.230 ;
        RECT 123.955 40.480 125.055 41.250 ;
        RECT 23.055 33.380 23.385 38.400 ;
        RECT 34.335 33.380 34.665 38.400 ;
        RECT 45.625 38.380 45.965 38.430 ;
        RECT 56.845 38.380 57.185 38.430 ;
        RECT 68.045 38.380 68.385 38.430 ;
        RECT 79.395 38.420 79.675 40.380 ;
        RECT 90.635 38.440 90.915 40.400 ;
        RECT 101.845 38.460 102.125 40.420 ;
        RECT 113.045 38.500 113.325 40.460 ;
        RECT 124.255 38.520 124.535 40.480 ;
        RECT 45.625 33.360 45.955 38.380 ;
        RECT 56.845 33.360 57.175 38.380 ;
        RECT 68.045 33.360 68.375 38.380 ;
        RECT 79.335 38.370 79.675 38.420 ;
        RECT 90.575 38.390 90.915 38.440 ;
        RECT 101.785 38.410 102.125 38.460 ;
        RECT 112.985 38.450 113.325 38.500 ;
        RECT 124.195 38.470 124.535 38.520 ;
        RECT 79.335 33.350 79.665 38.370 ;
        RECT 90.575 33.370 90.905 38.390 ;
        RECT 101.785 33.390 102.115 38.410 ;
        RECT 112.985 33.430 113.315 38.450 ;
        RECT 124.195 33.450 124.525 38.470 ;
        RECT 145.080 18.760 146.200 18.930 ;
        RECT 145.070 14.920 146.200 18.760 ;
        RECT 145.030 13.970 146.200 14.920 ;
        RECT 145.030 13.900 146.150 13.970 ;
        RECT 93.550 0.180 94.840 1.530 ;
      LAYER met3 ;
        RECT 93.500 0.205 94.890 1.505 ;
      LAYER met4 ;
        RECT 93.545 0.225 94.845 1.485 ;
        RECT 93.850 0.000 94.750 0.225 ;
    END
  END iop
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN reset
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER li1 ;
        RECT 122.895 168.515 123.255 169.095 ;
      LAYER met1 ;
        RECT 138.130 223.810 139.580 225.110 ;
        RECT 133.500 172.050 136.690 172.190 ;
        RECT 129.260 171.930 136.690 172.050 ;
        RECT 138.330 171.930 139.470 223.810 ;
        RECT 129.260 170.790 139.470 171.930 ;
        RECT 133.500 170.600 136.690 170.790 ;
        RECT 122.845 168.690 123.135 168.735 ;
        RECT 128.350 168.690 128.670 168.750 ;
        RECT 122.845 168.550 128.670 168.690 ;
        RECT 122.845 168.505 123.135 168.550 ;
        RECT 128.350 168.490 128.670 168.550 ;
      LAYER met2 ;
        RECT 138.180 223.760 139.530 225.160 ;
        RECT 128.370 171.325 128.650 171.695 ;
        RECT 128.440 168.780 128.580 171.325 ;
        RECT 129.310 170.740 133.650 172.100 ;
        RECT 128.380 168.460 128.640 168.780 ;
      LAYER met3 ;
        RECT 138.130 223.785 139.580 225.135 ;
        RECT 128.345 171.660 128.675 171.675 ;
        RECT 129.260 171.660 133.700 172.075 ;
        RECT 128.345 171.360 133.700 171.660 ;
        RECT 128.345 171.345 128.675 171.360 ;
        RECT 129.260 170.765 133.700 171.360 ;
      LAYER met4 ;
        RECT 138.310 225.115 138.610 225.760 ;
        RECT 138.175 223.805 139.535 225.115 ;
    END
  END reset
  PIN ua[0]
    ANTENNAGATEAREA 200.000000 ;
    PORT
      LAYER li1 ;
        RECT 27.895 65.555 28.895 65.725 ;
        RECT 39.095 65.565 40.095 65.735 ;
        RECT 50.315 65.535 51.315 65.705 ;
        RECT 61.565 65.515 62.565 65.685 ;
        RECT 72.785 65.505 73.785 65.675 ;
        RECT 84.025 65.495 85.025 65.665 ;
        RECT 95.275 65.505 96.275 65.675 ;
        RECT 106.555 65.495 107.555 65.665 ;
        RECT 117.825 65.495 118.825 65.665 ;
        RECT 129.075 65.495 130.075 65.665 ;
        RECT 19.845 19.685 20.845 19.855 ;
        RECT 31.125 19.685 32.125 19.855 ;
        RECT 42.415 19.665 43.415 19.835 ;
        RECT 53.635 19.665 54.635 19.835 ;
        RECT 64.835 19.665 65.835 19.835 ;
        RECT 76.125 19.655 77.125 19.825 ;
        RECT 87.365 19.675 88.365 19.845 ;
        RECT 98.575 19.695 99.575 19.865 ;
        RECT 109.775 19.735 110.775 19.905 ;
        RECT 120.985 19.755 121.985 19.925 ;
      LAYER met1 ;
        RECT 29.655 68.100 43.325 68.110 ;
        RECT 13.950 68.080 43.325 68.100 ;
        RECT 13.950 68.060 54.545 68.080 ;
        RECT 13.950 68.050 65.795 68.060 ;
        RECT 13.950 68.040 77.015 68.050 ;
        RECT 85.835 68.040 99.505 68.050 ;
        RECT 139.530 68.040 143.320 68.060 ;
        RECT 13.950 66.960 152.870 68.040 ;
        RECT 13.950 66.950 32.125 66.960 ;
        RECT 13.950 18.530 15.100 66.950 ;
        RECT 40.875 66.930 152.870 66.960 ;
        RECT 52.125 66.910 152.870 66.930 ;
        RECT 63.345 66.900 152.870 66.910 ;
        RECT 74.585 66.890 88.255 66.900 ;
        RECT 97.115 66.890 143.320 66.900 ;
        RECT 27.815 65.490 28.965 65.800 ;
        RECT 39.015 65.500 40.165 65.810 ;
        RECT 50.235 65.470 51.385 65.780 ;
        RECT 61.485 65.450 62.635 65.760 ;
        RECT 72.705 65.440 73.855 65.750 ;
        RECT 83.945 65.430 85.095 65.740 ;
        RECT 95.195 65.440 96.345 65.750 ;
        RECT 106.475 65.430 107.625 65.740 ;
        RECT 117.745 65.430 118.895 65.740 ;
        RECT 128.995 65.430 130.145 65.740 ;
        RECT 19.775 19.610 20.925 19.920 ;
        RECT 31.055 19.610 32.205 19.920 ;
        RECT 42.345 19.590 43.495 19.900 ;
        RECT 53.565 19.590 54.715 19.900 ;
        RECT 64.765 19.590 65.915 19.900 ;
        RECT 76.055 19.580 77.205 19.890 ;
        RECT 87.295 19.600 88.445 19.910 ;
        RECT 98.505 19.620 99.655 19.930 ;
        RECT 109.705 19.660 110.855 19.970 ;
        RECT 120.915 19.680 122.065 19.990 ;
        RECT 13.940 18.460 17.635 18.530 ;
        RECT 117.755 18.510 131.425 18.530 ;
        RECT 106.545 18.470 131.425 18.510 ;
        RECT 13.940 18.440 41.565 18.460 ;
        RECT 95.345 18.450 131.425 18.470 ;
        RECT 13.940 18.430 75.275 18.440 ;
        RECT 84.135 18.430 131.425 18.450 ;
        RECT 13.940 17.380 131.425 18.430 ;
        RECT 13.950 17.370 15.100 17.380 ;
        RECT 16.615 17.360 120.215 17.380 ;
        RECT 16.615 17.320 109.015 17.360 ;
        RECT 16.615 17.310 97.805 17.320 ;
        RECT 39.185 17.300 97.805 17.310 ;
        RECT 39.185 17.290 86.565 17.300 ;
        RECT 72.895 17.280 86.565 17.290 ;
        RECT 151.730 1.420 152.870 66.900 ;
        RECT 151.600 0.300 152.970 1.420 ;
      LAYER met2 ;
        RECT 27.795 67.130 28.915 67.810 ;
        RECT 38.995 67.140 40.115 67.820 ;
        RECT 28.075 65.850 28.745 67.130 ;
        RECT 39.275 65.860 39.945 67.140 ;
        RECT 50.215 67.110 51.335 67.790 ;
        RECT 27.865 65.440 28.915 65.850 ;
        RECT 39.065 65.450 40.115 65.860 ;
        RECT 50.495 65.830 51.165 67.110 ;
        RECT 61.465 67.090 62.585 67.770 ;
        RECT 50.285 65.420 51.335 65.830 ;
        RECT 61.745 65.810 62.415 67.090 ;
        RECT 72.685 67.080 73.805 67.760 ;
        RECT 61.535 65.400 62.585 65.810 ;
        RECT 72.965 65.800 73.635 67.080 ;
        RECT 83.925 67.070 85.045 67.750 ;
        RECT 95.175 67.080 96.295 67.760 ;
        RECT 72.755 65.390 73.805 65.800 ;
        RECT 84.205 65.790 84.875 67.070 ;
        RECT 95.455 65.800 96.125 67.080 ;
        RECT 106.455 67.070 107.575 67.750 ;
        RECT 117.725 67.070 118.845 67.750 ;
        RECT 128.975 67.070 130.095 67.750 ;
        RECT 83.995 65.380 85.045 65.790 ;
        RECT 95.245 65.390 96.295 65.800 ;
        RECT 106.735 65.790 107.405 67.070 ;
        RECT 118.005 65.790 118.675 67.070 ;
        RECT 129.255 65.790 129.925 67.070 ;
        RECT 106.525 65.380 107.575 65.790 ;
        RECT 117.795 65.380 118.845 65.790 ;
        RECT 129.045 65.380 130.095 65.790 ;
        RECT 19.825 19.560 20.875 19.970 ;
        RECT 31.105 19.560 32.155 19.970 ;
        RECT 19.995 18.280 20.665 19.560 ;
        RECT 31.275 18.280 31.945 19.560 ;
        RECT 42.395 19.540 43.445 19.950 ;
        RECT 53.615 19.540 54.665 19.950 ;
        RECT 64.815 19.540 65.865 19.950 ;
        RECT 19.825 17.600 20.945 18.280 ;
        RECT 31.105 17.600 32.225 18.280 ;
        RECT 42.565 18.260 43.235 19.540 ;
        RECT 53.785 18.260 54.455 19.540 ;
        RECT 64.985 18.260 65.655 19.540 ;
        RECT 76.105 19.530 77.155 19.940 ;
        RECT 87.345 19.550 88.395 19.960 ;
        RECT 98.555 19.570 99.605 19.980 ;
        RECT 109.755 19.610 110.805 20.020 ;
        RECT 120.965 19.630 122.015 20.040 ;
        RECT 42.395 17.580 43.515 18.260 ;
        RECT 53.615 17.580 54.735 18.260 ;
        RECT 64.815 17.580 65.935 18.260 ;
        RECT 76.275 18.250 76.945 19.530 ;
        RECT 87.515 18.270 88.185 19.550 ;
        RECT 98.725 18.290 99.395 19.570 ;
        RECT 109.925 18.330 110.595 19.610 ;
        RECT 121.135 18.350 121.805 19.630 ;
        RECT 76.105 17.570 77.225 18.250 ;
        RECT 87.345 17.590 88.465 18.270 ;
        RECT 98.555 17.610 99.675 18.290 ;
        RECT 109.755 17.650 110.875 18.330 ;
        RECT 120.965 17.670 122.085 18.350 ;
        RECT 151.650 0.250 152.920 1.470 ;
      LAYER met3 ;
        RECT 151.600 0.275 152.970 1.445 ;
      LAYER met4 ;
        RECT 151.645 0.295 152.925 1.425 ;
        RECT 151.810 0.000 152.710 0.295 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER li1 ;
        RECT 21.465 65.555 26.465 65.725 ;
        RECT 32.665 65.565 37.665 65.735 ;
        RECT 43.885 65.535 48.885 65.705 ;
        RECT 55.135 65.515 60.135 65.685 ;
        RECT 66.355 65.505 71.355 65.675 ;
        RECT 77.595 65.495 82.595 65.665 ;
        RECT 88.845 65.505 93.845 65.675 ;
        RECT 100.125 65.495 105.125 65.665 ;
        RECT 111.395 65.495 116.395 65.665 ;
        RECT 122.645 65.495 127.645 65.665 ;
        RECT 133.395 65.465 138.395 65.635 ;
        RECT 138.455 55.210 138.625 65.250 ;
      LAYER met1 ;
        RECT 29.645 69.670 43.315 69.680 ;
        RECT 18.445 69.650 43.315 69.670 ;
        RECT 18.445 69.630 54.535 69.650 ;
        RECT 18.445 69.620 65.785 69.630 ;
        RECT 139.590 69.620 150.610 69.640 ;
        RECT 18.445 69.610 77.005 69.620 ;
        RECT 85.825 69.610 99.495 69.620 ;
        RECT 132.155 69.610 150.610 69.620 ;
        RECT 18.445 69.570 150.610 69.610 ;
        RECT 18.445 68.530 150.740 69.570 ;
        RECT 18.445 68.520 32.115 68.530 ;
        RECT 40.865 68.500 150.740 68.530 ;
        RECT 52.115 68.490 143.320 68.500 ;
        RECT 52.115 68.480 140.670 68.490 ;
        RECT 63.335 68.470 140.670 68.480 ;
        RECT 149.360 68.470 150.740 68.500 ;
        RECT 74.575 68.460 88.245 68.470 ;
        RECT 97.105 68.460 133.295 68.470 ;
        RECT 21.405 65.510 26.555 65.790 ;
        RECT 32.605 65.520 37.755 65.800 ;
        RECT 43.825 65.490 48.975 65.770 ;
        RECT 149.460 65.760 150.600 65.780 ;
        RECT 55.075 65.470 60.225 65.750 ;
        RECT 66.295 65.460 71.445 65.740 ;
        RECT 77.535 65.450 82.685 65.730 ;
        RECT 88.785 65.460 93.935 65.740 ;
        RECT 100.065 65.450 105.215 65.730 ;
        RECT 111.335 65.450 116.485 65.730 ;
        RECT 122.585 65.450 127.735 65.730 ;
        RECT 133.315 65.430 138.455 65.690 ;
        RECT 138.425 65.100 138.655 65.230 ;
        RECT 138.345 55.130 138.725 65.100 ;
        RECT 149.340 64.660 150.720 65.760 ;
        RECT 149.460 2.770 150.600 64.660 ;
        RECT 131.940 1.880 150.600 2.770 ;
        RECT 131.800 1.630 150.600 1.880 ;
        RECT 131.800 1.380 133.490 1.630 ;
        RECT 131.800 0.430 133.540 1.380 ;
      LAYER met2 ;
        RECT 22.695 68.620 25.405 69.470 ;
        RECT 33.895 68.630 36.605 69.480 ;
        RECT 22.895 65.840 24.825 68.620 ;
        RECT 34.095 65.850 36.025 68.630 ;
        RECT 45.115 68.600 47.825 69.450 ;
        RECT 21.455 65.460 26.505 65.840 ;
        RECT 32.655 65.470 37.705 65.850 ;
        RECT 45.315 65.820 47.245 68.600 ;
        RECT 56.365 68.580 59.075 69.430 ;
        RECT 43.875 65.440 48.925 65.820 ;
        RECT 56.565 65.800 58.495 68.580 ;
        RECT 67.585 68.570 70.295 69.420 ;
        RECT 55.125 65.420 60.175 65.800 ;
        RECT 67.785 65.790 69.715 68.570 ;
        RECT 78.825 68.560 81.535 69.410 ;
        RECT 90.075 68.570 92.785 69.420 ;
        RECT 66.345 65.410 71.395 65.790 ;
        RECT 79.025 65.780 80.955 68.560 ;
        RECT 90.275 65.790 92.205 68.570 ;
        RECT 101.355 68.560 104.065 69.410 ;
        RECT 112.625 68.560 115.335 69.410 ;
        RECT 123.875 68.560 126.585 69.410 ;
        RECT 137.675 68.690 139.075 69.460 ;
        RECT 77.585 65.400 82.635 65.780 ;
        RECT 88.835 65.410 93.885 65.790 ;
        RECT 101.555 65.780 103.485 68.560 ;
        RECT 112.825 65.780 114.755 68.560 ;
        RECT 124.075 65.780 126.005 68.560 ;
        RECT 100.115 65.400 105.165 65.780 ;
        RECT 111.385 65.400 116.435 65.780 ;
        RECT 122.635 65.400 127.685 65.780 ;
        RECT 138.385 65.740 138.645 68.690 ;
        RECT 149.410 68.420 150.690 69.620 ;
        RECT 149.480 65.810 150.640 68.420 ;
        RECT 133.365 65.380 138.645 65.740 ;
        RECT 138.385 65.150 138.645 65.380 ;
        RECT 138.385 64.770 138.675 65.150 ;
        RECT 138.395 55.080 138.675 64.770 ;
        RECT 149.390 64.610 150.670 65.810 ;
        RECT 131.850 0.380 133.490 1.930 ;
      LAYER met3 ;
        RECT 131.800 0.405 133.540 1.905 ;
      LAYER met4 ;
        RECT 131.845 0.425 133.495 1.885 ;
        RECT 132.490 0.000 133.390 0.425 ;
    END
  END ua[1]
  PIN vdd
    ANTENNAGATEAREA 774.872986 ;
    ANTENNADIFFAREA 1141.909790 ;
    PORT
      LAYER nwell ;
        RECT 14.470 207.155 128.010 209.985 ;
        RECT 14.470 201.715 128.010 204.545 ;
        RECT 14.470 196.275 128.010 199.105 ;
        RECT 14.470 190.835 128.010 193.665 ;
        RECT 14.470 185.395 128.010 188.225 ;
        RECT 14.470 179.955 128.010 182.785 ;
        RECT 14.470 174.515 128.010 177.345 ;
        RECT 14.470 169.075 128.010 171.905 ;
        RECT 14.470 163.635 128.010 166.465 ;
        RECT 14.470 158.195 128.010 161.025 ;
        RECT 14.470 152.755 128.010 155.585 ;
        RECT 14.470 147.315 128.010 150.145 ;
        RECT 14.470 141.875 128.010 144.705 ;
        RECT 14.470 136.435 128.010 139.265 ;
        RECT 14.470 130.995 128.010 133.825 ;
        RECT 14.470 125.555 128.010 128.385 ;
        RECT 14.470 120.115 128.010 122.945 ;
        RECT 14.470 114.675 128.010 117.505 ;
        RECT 14.470 109.235 128.010 112.065 ;
        RECT 14.470 103.795 128.010 106.625 ;
        RECT 14.470 99.580 128.010 101.185 ;
        RECT 20.485 54.580 29.875 66.420 ;
        RECT 31.685 54.590 41.075 66.430 ;
        RECT 42.905 54.560 52.295 66.400 ;
        RECT 54.155 54.540 63.545 66.380 ;
        RECT 65.375 54.530 74.765 66.370 ;
        RECT 76.615 54.520 86.005 66.360 ;
        RECT 87.865 54.530 97.255 66.370 ;
        RECT 99.145 54.520 108.535 66.360 ;
        RECT 110.415 54.520 119.805 66.360 ;
        RECT 121.665 54.520 131.055 66.360 ;
        RECT 132.415 54.490 139.375 66.330 ;
        RECT 20.655 49.020 23.115 53.210 ;
        RECT 24.735 45.940 29.125 53.130 ;
        RECT 31.855 49.030 34.315 53.220 ;
        RECT 35.935 45.950 40.325 53.140 ;
        RECT 43.075 49.000 45.535 53.190 ;
        RECT 47.155 45.920 51.545 53.110 ;
        RECT 54.325 48.980 56.785 53.170 ;
        RECT 58.405 45.900 62.795 53.090 ;
        RECT 65.545 48.970 68.005 53.160 ;
        RECT 69.625 45.890 74.015 53.080 ;
        RECT 76.785 48.960 79.245 53.150 ;
        RECT 80.865 45.880 85.255 53.070 ;
        RECT 88.035 48.970 90.495 53.160 ;
        RECT 92.115 45.890 96.505 53.080 ;
        RECT 99.315 48.960 101.775 53.150 ;
        RECT 103.395 45.880 107.785 53.070 ;
        RECT 110.585 48.960 113.045 53.150 ;
        RECT 114.665 45.880 119.055 53.070 ;
        RECT 121.835 48.960 124.295 53.150 ;
        RECT 125.915 45.880 130.305 53.070 ;
        RECT 19.615 32.280 24.005 39.470 ;
        RECT 25.625 32.200 28.085 36.390 ;
        RECT 30.895 32.280 35.285 39.470 ;
        RECT 36.905 32.200 39.365 36.390 ;
        RECT 42.185 32.260 46.575 39.450 ;
        RECT 48.195 32.180 50.655 36.370 ;
        RECT 53.405 32.260 57.795 39.450 ;
        RECT 59.415 32.180 61.875 36.370 ;
        RECT 64.605 32.260 68.995 39.450 ;
        RECT 70.615 32.180 73.075 36.370 ;
        RECT 75.895 32.250 80.285 39.440 ;
        RECT 81.905 32.170 84.365 36.360 ;
        RECT 87.135 32.270 91.525 39.460 ;
        RECT 93.145 32.190 95.605 36.380 ;
        RECT 98.345 32.290 102.735 39.480 ;
        RECT 104.355 32.210 106.815 36.400 ;
        RECT 109.545 32.330 113.935 39.520 ;
        RECT 115.555 32.250 118.015 36.440 ;
        RECT 120.755 32.350 125.145 39.540 ;
        RECT 126.765 32.270 129.225 36.460 ;
        RECT 18.865 18.990 28.255 30.830 ;
        RECT 30.145 18.990 39.535 30.830 ;
        RECT 41.435 18.970 50.825 30.810 ;
        RECT 52.655 18.970 62.045 30.810 ;
        RECT 63.855 18.970 73.245 30.810 ;
        RECT 75.145 18.960 84.535 30.800 ;
        RECT 86.385 18.980 95.775 30.820 ;
        RECT 97.595 19.000 106.985 30.840 ;
        RECT 108.795 19.040 118.185 30.880 ;
        RECT 120.005 19.060 129.395 30.900 ;
        RECT 131.725 19.030 138.685 30.870 ;
      LAYER li1 ;
        RECT 15.435 209.745 15.955 210.285 ;
        RECT 14.745 208.655 15.955 209.745 ;
        RECT 16.125 209.745 17.335 210.265 ;
        RECT 16.125 208.655 18.715 209.745 ;
        RECT 20.480 209.090 20.830 210.340 ;
        RECT 18.890 208.655 24.235 209.090 ;
        RECT 24.405 208.655 24.695 209.820 ;
        RECT 24.865 209.745 25.385 210.285 ;
        RECT 24.865 208.655 26.075 209.745 ;
        RECT 27.840 209.090 28.190 210.340 ;
        RECT 33.360 209.090 33.710 210.340 ;
        RECT 26.250 208.655 31.595 209.090 ;
        RECT 31.770 208.655 37.115 209.090 ;
        RECT 37.285 208.655 37.575 209.820 ;
        RECT 37.745 209.745 38.265 210.285 ;
        RECT 37.745 208.655 38.955 209.745 ;
        RECT 40.720 209.090 41.070 210.340 ;
        RECT 46.240 209.090 46.590 210.340 ;
        RECT 39.130 208.655 44.475 209.090 ;
        RECT 44.650 208.655 49.995 209.090 ;
        RECT 50.165 208.655 50.455 209.820 ;
        RECT 50.625 209.745 51.145 210.285 ;
        RECT 50.625 208.655 51.835 209.745 ;
        RECT 53.600 209.090 53.950 210.340 ;
        RECT 59.120 209.090 59.470 210.340 ;
        RECT 52.010 208.655 57.355 209.090 ;
        RECT 57.530 208.655 62.875 209.090 ;
        RECT 63.045 208.655 63.335 209.820 ;
        RECT 63.505 209.745 64.025 210.285 ;
        RECT 63.505 208.655 64.715 209.745 ;
        RECT 66.480 209.090 66.830 210.340 ;
        RECT 72.000 209.090 72.350 210.340 ;
        RECT 64.890 208.655 70.235 209.090 ;
        RECT 70.410 208.655 75.755 209.090 ;
        RECT 75.925 208.655 76.215 209.820 ;
        RECT 76.385 209.745 76.905 210.285 ;
        RECT 76.385 208.655 77.595 209.745 ;
        RECT 79.360 209.090 79.710 210.340 ;
        RECT 84.880 209.090 85.230 210.340 ;
        RECT 77.770 208.655 83.115 209.090 ;
        RECT 83.290 208.655 88.635 209.090 ;
        RECT 88.805 208.655 89.095 209.820 ;
        RECT 89.265 209.745 89.785 210.285 ;
        RECT 89.265 208.655 90.475 209.745 ;
        RECT 92.240 209.090 92.590 210.340 ;
        RECT 97.760 209.090 98.110 210.340 ;
        RECT 90.650 208.655 95.995 209.090 ;
        RECT 96.170 208.655 101.515 209.090 ;
        RECT 101.685 208.655 101.975 209.820 ;
        RECT 102.145 209.745 102.665 210.285 ;
        RECT 102.145 208.655 103.355 209.745 ;
        RECT 105.120 209.090 105.470 210.340 ;
        RECT 110.640 209.090 110.990 210.340 ;
        RECT 103.530 208.655 108.875 209.090 ;
        RECT 109.050 208.655 114.395 209.090 ;
        RECT 114.565 208.655 114.855 209.820 ;
        RECT 117.080 209.090 117.430 210.340 ;
        RECT 122.600 209.090 122.950 210.340 ;
        RECT 126.525 209.745 127.045 210.285 ;
        RECT 115.490 208.655 120.835 209.090 ;
        RECT 121.010 208.655 126.355 209.090 ;
        RECT 126.525 208.655 127.735 209.745 ;
        RECT 14.660 208.485 127.820 208.655 ;
        RECT 14.745 207.395 15.955 208.485 ;
        RECT 15.435 206.855 15.955 207.395 ;
        RECT 16.125 207.395 18.715 208.485 ;
        RECT 18.890 208.050 24.235 208.485 ;
        RECT 16.125 206.875 17.335 207.395 ;
        RECT 20.480 206.800 20.830 208.050 ;
        RECT 24.405 207.320 24.695 208.485 ;
        RECT 25.325 207.395 27.915 208.485 ;
        RECT 28.090 208.050 33.435 208.485 ;
        RECT 33.610 208.050 38.955 208.485 ;
        RECT 39.130 208.050 44.475 208.485 ;
        RECT 44.650 208.050 49.995 208.485 ;
        RECT 25.325 206.875 26.535 207.395 ;
        RECT 29.680 206.800 30.030 208.050 ;
        RECT 35.200 206.800 35.550 208.050 ;
        RECT 40.720 206.800 41.070 208.050 ;
        RECT 46.240 206.800 46.590 208.050 ;
        RECT 50.165 207.320 50.455 208.485 ;
        RECT 50.625 207.395 52.295 208.485 ;
        RECT 52.470 208.050 57.815 208.485 ;
        RECT 57.990 208.050 63.335 208.485 ;
        RECT 63.510 208.050 68.855 208.485 ;
        RECT 69.030 208.050 74.375 208.485 ;
        RECT 50.625 206.875 51.375 207.395 ;
        RECT 54.060 206.800 54.410 208.050 ;
        RECT 59.580 206.800 59.930 208.050 ;
        RECT 65.100 206.800 65.450 208.050 ;
        RECT 70.620 206.800 70.970 208.050 ;
        RECT 74.585 207.345 74.815 208.485 ;
        RECT 75.485 207.345 75.695 208.485 ;
        RECT 75.925 207.320 76.215 208.485 ;
        RECT 76.385 207.395 77.595 208.485 ;
        RECT 77.785 207.975 78.085 208.485 ;
        RECT 79.215 207.975 79.845 208.485 ;
        RECT 80.515 207.975 80.815 208.485 ;
        RECT 81.445 207.395 84.955 208.485 ;
        RECT 85.130 208.050 90.475 208.485 ;
        RECT 90.650 208.050 95.995 208.485 ;
        RECT 96.170 208.050 101.515 208.485 ;
        RECT 76.385 206.855 76.905 207.395 ;
        RECT 81.445 206.875 83.135 207.395 ;
        RECT 86.720 206.800 87.070 208.050 ;
        RECT 92.240 206.800 92.590 208.050 ;
        RECT 97.760 206.800 98.110 208.050 ;
        RECT 101.685 207.320 101.975 208.485 ;
        RECT 102.605 207.395 104.275 208.485 ;
        RECT 104.450 208.050 109.795 208.485 ;
        RECT 109.970 208.050 115.315 208.485 ;
        RECT 115.490 208.050 120.835 208.485 ;
        RECT 121.010 208.050 126.355 208.485 ;
        RECT 102.605 206.875 103.355 207.395 ;
        RECT 106.040 206.800 106.390 208.050 ;
        RECT 111.560 206.800 111.910 208.050 ;
        RECT 117.080 206.800 117.430 208.050 ;
        RECT 122.600 206.800 122.950 208.050 ;
        RECT 126.525 207.395 127.735 208.485 ;
        RECT 126.525 206.855 127.045 207.395 ;
        RECT 15.435 204.305 15.955 204.845 ;
        RECT 14.745 203.215 15.955 204.305 ;
        RECT 17.045 204.305 18.735 204.825 ;
        RECT 17.045 203.215 20.555 204.305 ;
        RECT 22.320 203.650 22.670 204.900 ;
        RECT 27.840 203.650 28.190 204.900 ;
        RECT 33.360 203.650 33.710 204.900 ;
        RECT 20.730 203.215 26.075 203.650 ;
        RECT 26.250 203.215 31.595 203.650 ;
        RECT 31.770 203.215 37.115 203.650 ;
        RECT 37.285 203.215 37.575 204.380 ;
        RECT 38.205 204.305 39.415 204.825 ;
        RECT 38.205 203.215 40.795 204.305 ;
        RECT 42.560 203.650 42.910 204.900 ;
        RECT 48.080 203.650 48.430 204.900 ;
        RECT 53.600 203.650 53.950 204.900 ;
        RECT 59.120 203.650 59.470 204.900 ;
        RECT 40.970 203.215 46.315 203.650 ;
        RECT 46.490 203.215 51.835 203.650 ;
        RECT 52.010 203.215 57.355 203.650 ;
        RECT 57.530 203.215 62.875 203.650 ;
        RECT 63.045 203.215 63.335 204.380 ;
        RECT 63.505 204.305 64.255 204.825 ;
        RECT 63.505 203.215 65.175 204.305 ;
        RECT 65.405 203.215 65.615 204.355 ;
        RECT 66.285 203.215 66.515 204.355 ;
        RECT 67.225 203.215 67.455 204.355 ;
        RECT 68.125 203.215 68.335 204.355 ;
        RECT 68.995 203.215 69.300 204.355 ;
        RECT 69.640 203.215 69.970 203.595 ;
        RECT 70.490 203.215 70.740 203.675 ;
        RECT 72.355 203.215 72.725 203.675 ;
        RECT 73.360 203.215 73.690 203.645 ;
        RECT 75.580 203.215 75.830 203.675 ;
        RECT 76.835 203.215 77.165 203.715 ;
        RECT 78.195 203.215 78.500 204.355 ;
        RECT 86.965 204.305 87.715 204.825 ;
        RECT 78.840 203.215 79.170 203.595 ;
        RECT 79.690 203.215 79.940 203.675 ;
        RECT 81.555 203.215 81.925 203.675 ;
        RECT 82.560 203.215 82.890 203.645 ;
        RECT 84.780 203.215 85.030 203.675 ;
        RECT 86.035 203.215 86.365 203.715 ;
        RECT 86.965 203.215 88.635 204.305 ;
        RECT 88.805 203.215 89.095 204.380 ;
        RECT 89.725 204.305 90.935 204.825 ;
        RECT 89.725 203.215 92.315 204.305 ;
        RECT 94.080 203.650 94.430 204.900 ;
        RECT 99.600 203.650 99.950 204.900 ;
        RECT 105.120 203.650 105.470 204.900 ;
        RECT 110.640 203.650 110.990 204.900 ;
        RECT 92.490 203.215 97.835 203.650 ;
        RECT 98.010 203.215 103.355 203.650 ;
        RECT 103.530 203.215 108.875 203.650 ;
        RECT 109.050 203.215 114.395 203.650 ;
        RECT 114.565 203.215 114.855 204.380 ;
        RECT 117.080 203.650 117.430 204.900 ;
        RECT 122.600 203.650 122.950 204.900 ;
        RECT 126.525 204.305 127.045 204.845 ;
        RECT 115.490 203.215 120.835 203.650 ;
        RECT 121.010 203.215 126.355 203.650 ;
        RECT 126.525 203.215 127.735 204.305 ;
        RECT 14.660 203.045 127.820 203.215 ;
        RECT 14.745 201.955 15.955 203.045 ;
        RECT 15.435 201.415 15.955 201.955 ;
        RECT 16.125 201.955 18.715 203.045 ;
        RECT 18.890 202.610 24.235 203.045 ;
        RECT 16.125 201.435 17.335 201.955 ;
        RECT 20.480 201.360 20.830 202.610 ;
        RECT 24.405 201.880 24.695 203.045 ;
        RECT 25.325 201.955 27.915 203.045 ;
        RECT 28.090 202.610 33.435 203.045 ;
        RECT 33.610 202.610 38.955 203.045 ;
        RECT 39.130 202.610 44.475 203.045 ;
        RECT 44.650 202.610 49.995 203.045 ;
        RECT 25.325 201.435 26.535 201.955 ;
        RECT 29.680 201.360 30.030 202.610 ;
        RECT 35.200 201.360 35.550 202.610 ;
        RECT 40.720 201.360 41.070 202.610 ;
        RECT 46.240 201.360 46.590 202.610 ;
        RECT 50.165 201.880 50.455 203.045 ;
        RECT 51.085 201.955 54.595 203.045 ;
        RECT 54.770 202.610 60.115 203.045 ;
        RECT 51.085 201.435 52.775 201.955 ;
        RECT 56.360 201.360 56.710 202.610 ;
        RECT 60.715 202.545 61.045 203.045 ;
        RECT 62.050 202.585 62.300 203.045 ;
        RECT 64.190 202.615 64.520 203.045 ;
        RECT 65.155 202.585 65.525 203.045 ;
        RECT 67.140 202.585 67.390 203.045 ;
        RECT 67.910 202.665 68.240 203.045 ;
        RECT 68.535 201.985 68.705 203.045 ;
        RECT 69.375 202.205 69.545 203.045 ;
        RECT 70.215 202.205 70.385 203.045 ;
        RECT 71.305 202.265 71.635 203.045 ;
        RECT 72.195 202.620 72.530 203.045 ;
        RECT 73.180 202.285 73.510 203.045 ;
        RECT 74.110 201.895 74.370 203.045 ;
        RECT 74.545 201.955 75.755 203.045 ;
        RECT 74.545 201.415 75.065 201.955 ;
        RECT 75.925 201.880 76.215 203.045 ;
        RECT 76.825 202.265 77.155 203.045 ;
        RECT 77.715 202.620 78.050 203.045 ;
        RECT 78.665 202.285 78.995 203.045 ;
        RECT 80.035 201.905 80.340 203.045 ;
        RECT 80.680 202.665 81.010 203.045 ;
        RECT 81.530 202.585 81.780 203.045 ;
        RECT 83.395 202.585 83.765 203.045 ;
        RECT 84.400 202.615 84.730 203.045 ;
        RECT 86.620 202.585 86.870 203.045 ;
        RECT 87.875 202.545 88.205 203.045 ;
        RECT 88.805 201.955 90.475 203.045 ;
        RECT 90.650 202.610 95.995 203.045 ;
        RECT 96.170 202.610 101.515 203.045 ;
        RECT 88.805 201.435 89.555 201.955 ;
        RECT 92.240 201.360 92.590 202.610 ;
        RECT 97.760 201.360 98.110 202.610 ;
        RECT 101.685 201.880 101.975 203.045 ;
        RECT 102.605 201.955 104.275 203.045 ;
        RECT 104.450 202.610 109.795 203.045 ;
        RECT 109.970 202.610 115.315 203.045 ;
        RECT 115.490 202.610 120.835 203.045 ;
        RECT 121.010 202.610 126.355 203.045 ;
        RECT 102.605 201.435 103.355 201.955 ;
        RECT 106.040 201.360 106.390 202.610 ;
        RECT 111.560 201.360 111.910 202.610 ;
        RECT 117.080 201.360 117.430 202.610 ;
        RECT 122.600 201.360 122.950 202.610 ;
        RECT 126.525 201.955 127.735 203.045 ;
        RECT 126.525 201.415 127.045 201.955 ;
        RECT 15.435 198.865 15.955 199.405 ;
        RECT 14.745 197.775 15.955 198.865 ;
        RECT 17.045 198.865 18.735 199.385 ;
        RECT 17.045 197.775 20.555 198.865 ;
        RECT 22.320 198.210 22.670 199.460 ;
        RECT 27.840 198.210 28.190 199.460 ;
        RECT 33.360 198.210 33.710 199.460 ;
        RECT 20.730 197.775 26.075 198.210 ;
        RECT 26.250 197.775 31.595 198.210 ;
        RECT 31.770 197.775 37.115 198.210 ;
        RECT 37.285 197.775 37.575 198.940 ;
        RECT 38.205 198.865 39.415 199.385 ;
        RECT 38.205 197.775 40.795 198.865 ;
        RECT 42.560 198.210 42.910 199.460 ;
        RECT 48.080 198.210 48.430 199.460 ;
        RECT 53.600 198.210 53.950 199.460 ;
        RECT 59.120 198.210 59.470 199.460 ;
        RECT 40.970 197.775 46.315 198.210 ;
        RECT 46.490 197.775 51.835 198.210 ;
        RECT 52.010 197.775 57.355 198.210 ;
        RECT 57.530 197.775 62.875 198.210 ;
        RECT 63.045 197.775 63.335 198.940 ;
        RECT 63.965 198.865 64.715 199.385 ;
        RECT 63.965 197.775 65.635 198.865 ;
        RECT 66.245 197.775 66.575 198.535 ;
        RECT 80.515 198.455 80.845 198.700 ;
        RECT 80.660 198.430 80.845 198.455 ;
        RECT 80.660 198.330 81.275 198.430 ;
        RECT 67.640 197.775 67.970 198.185 ;
        RECT 68.555 197.775 69.225 198.185 ;
        RECT 69.935 197.775 70.265 198.215 ;
        RECT 71.295 197.775 71.625 198.155 ;
        RECT 72.480 197.775 72.810 198.155 ;
        RECT 73.385 197.775 73.715 198.155 ;
        RECT 74.395 197.775 74.725 198.155 ;
        RECT 76.020 197.775 76.345 198.235 ;
        RECT 78.135 197.775 78.405 198.235 ;
        RECT 79.590 197.775 79.845 198.320 ;
        RECT 80.670 197.775 81.275 198.330 ;
        RECT 81.445 197.775 81.705 198.915 ;
        RECT 82.375 197.775 82.655 198.915 ;
        RECT 82.885 197.775 83.095 198.915 ;
        RECT 83.765 197.775 83.995 198.915 ;
        RECT 84.245 197.775 84.475 198.915 ;
        RECT 85.145 197.775 85.355 198.915 ;
        RECT 86.045 198.865 87.255 199.385 ;
        RECT 86.045 197.775 88.635 198.865 ;
        RECT 88.805 197.775 89.095 198.940 ;
        RECT 89.725 198.865 90.935 199.385 ;
        RECT 89.725 197.775 92.315 198.865 ;
        RECT 94.080 198.210 94.430 199.460 ;
        RECT 99.600 198.210 99.950 199.460 ;
        RECT 105.120 198.210 105.470 199.460 ;
        RECT 110.640 198.210 110.990 199.460 ;
        RECT 92.490 197.775 97.835 198.210 ;
        RECT 98.010 197.775 103.355 198.210 ;
        RECT 103.530 197.775 108.875 198.210 ;
        RECT 109.050 197.775 114.395 198.210 ;
        RECT 114.565 197.775 114.855 198.940 ;
        RECT 117.080 198.210 117.430 199.460 ;
        RECT 122.600 198.210 122.950 199.460 ;
        RECT 126.525 198.865 127.045 199.405 ;
        RECT 115.490 197.775 120.835 198.210 ;
        RECT 121.010 197.775 126.355 198.210 ;
        RECT 126.525 197.775 127.735 198.865 ;
        RECT 14.660 197.605 127.820 197.775 ;
        RECT 14.745 196.515 15.955 197.605 ;
        RECT 15.435 195.975 15.955 196.515 ;
        RECT 16.125 196.515 18.715 197.605 ;
        RECT 18.890 197.170 24.235 197.605 ;
        RECT 16.125 195.995 17.335 196.515 ;
        RECT 20.480 195.920 20.830 197.170 ;
        RECT 24.405 196.440 24.695 197.605 ;
        RECT 25.325 196.515 27.915 197.605 ;
        RECT 28.090 197.170 33.435 197.605 ;
        RECT 33.610 197.170 38.955 197.605 ;
        RECT 39.130 197.170 44.475 197.605 ;
        RECT 44.650 197.170 49.995 197.605 ;
        RECT 25.325 195.995 26.535 196.515 ;
        RECT 29.680 195.920 30.030 197.170 ;
        RECT 35.200 195.920 35.550 197.170 ;
        RECT 40.720 195.920 41.070 197.170 ;
        RECT 46.240 195.920 46.590 197.170 ;
        RECT 50.165 196.440 50.455 197.605 ;
        RECT 50.625 196.515 52.295 197.605 ;
        RECT 50.625 195.995 51.375 196.515 ;
        RECT 52.525 196.465 52.735 197.605 ;
        RECT 53.405 196.465 53.635 197.605 ;
        RECT 53.845 196.515 55.515 197.605 ;
        RECT 53.845 195.995 54.595 196.515 ;
        RECT 55.745 196.465 55.955 197.605 ;
        RECT 56.625 196.465 56.855 197.605 ;
        RECT 57.065 196.515 58.275 197.605 ;
        RECT 58.450 197.170 63.795 197.605 ;
        RECT 63.970 197.170 69.315 197.605 ;
        RECT 57.065 195.975 57.585 196.515 ;
        RECT 60.040 195.920 60.390 197.170 ;
        RECT 65.560 195.920 65.910 197.170 ;
        RECT 69.930 197.060 70.185 197.605 ;
        RECT 71.010 197.050 71.615 197.605 ;
        RECT 71.000 196.950 71.615 197.050 ;
        RECT 71.000 196.925 71.185 196.950 ;
        RECT 70.855 196.680 71.185 196.925 ;
        RECT 72.295 196.465 72.545 197.605 ;
        RECT 73.215 197.135 73.545 197.605 ;
        RECT 75.925 196.440 76.215 197.605 ;
        RECT 78.365 196.805 78.695 197.605 ;
        RECT 79.610 197.170 84.955 197.605 ;
        RECT 85.130 197.170 90.475 197.605 ;
        RECT 90.650 197.170 95.995 197.605 ;
        RECT 96.170 197.170 101.515 197.605 ;
        RECT 81.200 195.920 81.550 197.170 ;
        RECT 86.720 195.920 87.070 197.170 ;
        RECT 92.240 195.920 92.590 197.170 ;
        RECT 97.760 195.920 98.110 197.170 ;
        RECT 101.685 196.440 101.975 197.605 ;
        RECT 102.150 197.170 107.495 197.605 ;
        RECT 103.740 195.920 104.090 197.170 ;
        RECT 107.705 196.465 107.935 197.605 ;
        RECT 108.605 196.465 108.815 197.605 ;
        RECT 109.475 196.465 109.780 197.605 ;
        RECT 110.120 197.225 110.450 197.605 ;
        RECT 110.970 197.145 111.220 197.605 ;
        RECT 112.835 197.145 113.205 197.605 ;
        RECT 113.840 197.175 114.170 197.605 ;
        RECT 116.060 197.145 116.310 197.605 ;
        RECT 117.315 197.105 117.645 197.605 ;
        RECT 118.245 196.515 120.835 197.605 ;
        RECT 121.010 197.170 126.355 197.605 ;
        RECT 118.245 195.995 119.455 196.515 ;
        RECT 122.600 195.920 122.950 197.170 ;
        RECT 126.525 196.515 127.735 197.605 ;
        RECT 126.525 195.975 127.045 196.515 ;
        RECT 15.435 193.425 15.955 193.965 ;
        RECT 14.745 192.335 15.955 193.425 ;
        RECT 17.045 193.425 18.735 193.945 ;
        RECT 17.045 192.335 20.555 193.425 ;
        RECT 22.320 192.770 22.670 194.020 ;
        RECT 27.840 192.770 28.190 194.020 ;
        RECT 33.360 192.770 33.710 194.020 ;
        RECT 20.730 192.335 26.075 192.770 ;
        RECT 26.250 192.335 31.595 192.770 ;
        RECT 31.770 192.335 37.115 192.770 ;
        RECT 37.285 192.335 37.575 193.500 ;
        RECT 39.800 192.770 40.150 194.020 ;
        RECT 38.210 192.335 43.555 192.770 ;
        RECT 44.155 192.335 44.485 192.835 ;
        RECT 45.490 192.335 45.740 192.795 ;
        RECT 47.630 192.335 47.960 192.765 ;
        RECT 48.595 192.335 48.965 192.795 ;
        RECT 50.580 192.335 50.830 192.795 ;
        RECT 51.350 192.335 51.680 192.715 ;
        RECT 52.020 192.335 52.325 193.475 ;
        RECT 53.355 192.335 53.660 193.475 ;
        RECT 54.000 192.335 54.330 192.715 ;
        RECT 54.850 192.335 55.100 192.795 ;
        RECT 56.715 192.335 57.085 192.795 ;
        RECT 57.720 192.335 58.050 192.765 ;
        RECT 59.940 192.335 60.190 192.795 ;
        RECT 61.195 192.335 61.525 192.835 ;
        RECT 63.045 192.335 63.335 193.500 ;
        RECT 63.965 193.425 64.715 193.945 ;
        RECT 63.965 192.335 65.635 193.425 ;
        RECT 65.865 192.335 66.075 193.475 ;
        RECT 66.745 192.335 66.975 193.475 ;
        RECT 67.185 193.425 67.705 193.965 ;
        RECT 68.565 193.425 70.255 193.945 ;
        RECT 67.185 192.335 68.395 193.425 ;
        RECT 68.565 192.335 72.075 193.425 ;
        RECT 72.245 192.335 72.505 193.475 ;
        RECT 74.530 192.335 74.810 193.135 ;
        RECT 75.950 192.335 76.230 193.135 ;
        RECT 78.255 192.335 78.515 193.475 ;
        RECT 80.740 192.770 81.090 194.020 ;
        RECT 79.150 192.335 84.495 192.770 ;
        RECT 85.415 192.335 85.585 193.095 ;
        RECT 87.955 192.335 88.125 193.475 ;
        RECT 88.805 192.335 89.095 193.500 ;
        RECT 89.785 192.335 89.995 193.475 ;
        RECT 90.665 192.335 90.895 193.475 ;
        RECT 93.405 193.425 94.615 193.945 ;
        RECT 92.005 192.335 92.335 193.095 ;
        RECT 93.405 192.335 95.995 193.425 ;
        RECT 96.205 192.335 96.435 193.475 ;
        RECT 97.105 192.335 97.315 193.475 ;
        RECT 97.975 192.335 98.280 193.475 ;
        RECT 98.620 192.335 98.950 192.715 ;
        RECT 99.470 192.335 99.720 192.795 ;
        RECT 101.335 192.335 101.705 192.795 ;
        RECT 102.340 192.335 102.670 192.765 ;
        RECT 104.560 192.335 104.810 192.795 ;
        RECT 105.815 192.335 106.145 192.835 ;
        RECT 107.300 192.335 107.625 192.795 ;
        RECT 109.415 192.335 109.685 192.795 ;
        RECT 111.175 192.335 111.345 193.095 ;
        RECT 113.715 192.335 113.885 193.475 ;
        RECT 114.565 192.335 114.855 193.500 ;
        RECT 115.085 192.335 115.295 193.475 ;
        RECT 115.965 192.335 116.195 193.475 ;
        RECT 117.325 193.425 119.015 193.945 ;
        RECT 117.325 192.335 120.835 193.425 ;
        RECT 122.600 192.770 122.950 194.020 ;
        RECT 126.525 193.425 127.045 193.965 ;
        RECT 121.010 192.335 126.355 192.770 ;
        RECT 126.525 192.335 127.735 193.425 ;
        RECT 14.660 192.165 127.820 192.335 ;
        RECT 14.745 191.075 15.955 192.165 ;
        RECT 15.435 190.535 15.955 191.075 ;
        RECT 16.125 191.075 18.715 192.165 ;
        RECT 18.890 191.730 24.235 192.165 ;
        RECT 16.125 190.555 17.335 191.075 ;
        RECT 20.480 190.480 20.830 191.730 ;
        RECT 24.405 191.000 24.695 192.165 ;
        RECT 24.865 191.075 26.535 192.165 ;
        RECT 26.710 191.730 32.055 192.165 ;
        RECT 32.230 191.730 37.575 192.165 ;
        RECT 24.865 190.555 25.615 191.075 ;
        RECT 28.300 190.480 28.650 191.730 ;
        RECT 33.820 190.480 34.170 191.730 ;
        RECT 38.175 191.025 38.480 192.165 ;
        RECT 38.820 191.785 39.150 192.165 ;
        RECT 39.670 191.705 39.920 192.165 ;
        RECT 41.535 191.705 41.905 192.165 ;
        RECT 42.540 191.735 42.870 192.165 ;
        RECT 44.760 191.705 45.010 192.165 ;
        RECT 46.015 191.665 46.345 192.165 ;
        RECT 47.405 191.075 49.995 192.165 ;
        RECT 47.405 190.555 48.615 191.075 ;
        RECT 50.165 191.000 50.455 192.165 ;
        RECT 51.985 191.405 52.315 192.165 ;
        RECT 53.675 191.405 53.845 192.165 ;
        RECT 56.215 191.025 56.385 192.165 ;
        RECT 58.425 191.405 58.755 192.165 ;
        RECT 59.365 191.075 61.955 192.165 ;
        RECT 62.555 191.665 62.885 192.165 ;
        RECT 63.890 191.705 64.140 192.165 ;
        RECT 66.030 191.735 66.360 192.165 ;
        RECT 66.995 191.705 67.365 192.165 ;
        RECT 68.980 191.705 69.230 192.165 ;
        RECT 69.750 191.785 70.080 192.165 ;
        RECT 59.365 190.555 60.575 191.075 ;
        RECT 70.420 191.025 70.725 192.165 ;
        RECT 71.345 191.655 71.645 192.165 ;
        RECT 72.775 191.655 73.405 192.165 ;
        RECT 74.075 191.655 74.375 192.165 ;
        RECT 74.545 191.075 75.755 192.165 ;
        RECT 74.545 190.535 75.065 191.075 ;
        RECT 75.925 191.000 76.215 192.165 ;
        RECT 76.405 191.365 76.685 192.165 ;
        RECT 77.415 191.365 77.585 192.165 ;
        RECT 78.255 191.025 78.515 192.165 ;
        RECT 78.685 191.075 80.355 192.165 ;
        RECT 80.530 191.730 85.875 192.165 ;
        RECT 78.685 190.555 79.435 191.075 ;
        RECT 82.120 190.480 82.470 191.730 ;
        RECT 86.855 191.365 87.140 192.165 ;
        RECT 88.260 191.475 88.590 192.165 ;
        RECT 89.260 191.785 89.680 192.165 ;
        RECT 90.960 191.785 91.290 192.165 ;
        RECT 91.810 191.785 92.190 192.165 ;
        RECT 93.835 191.665 94.165 192.165 ;
        RECT 94.775 191.665 95.105 192.165 ;
        RECT 95.705 191.075 97.375 192.165 ;
        RECT 98.295 191.405 98.465 192.165 ;
        RECT 95.705 190.555 96.455 191.075 ;
        RECT 100.835 191.025 101.005 192.165 ;
        RECT 101.685 191.000 101.975 192.165 ;
        RECT 103.045 191.405 103.375 192.165 ;
        RECT 104.445 191.075 106.115 192.165 ;
        RECT 107.035 191.405 107.205 192.165 ;
        RECT 104.445 190.555 105.195 191.075 ;
        RECT 109.575 191.025 109.745 192.165 ;
        RECT 110.855 191.025 111.160 192.165 ;
        RECT 111.500 191.785 111.830 192.165 ;
        RECT 112.350 191.705 112.600 192.165 ;
        RECT 114.215 191.705 114.585 192.165 ;
        RECT 115.220 191.735 115.550 192.165 ;
        RECT 117.440 191.705 117.690 192.165 ;
        RECT 118.695 191.665 119.025 192.165 ;
        RECT 119.625 191.075 120.835 192.165 ;
        RECT 121.010 191.730 126.355 192.165 ;
        RECT 119.625 190.535 120.145 191.075 ;
        RECT 122.600 190.480 122.950 191.730 ;
        RECT 126.525 191.075 127.735 192.165 ;
        RECT 126.525 190.535 127.045 191.075 ;
        RECT 15.435 187.985 15.955 188.525 ;
        RECT 14.745 186.895 15.955 187.985 ;
        RECT 16.125 187.985 16.875 188.505 ;
        RECT 16.125 186.895 17.795 187.985 ;
        RECT 19.560 187.330 19.910 188.580 ;
        RECT 25.080 187.330 25.430 188.580 ;
        RECT 17.970 186.895 23.315 187.330 ;
        RECT 23.490 186.895 28.835 187.330 ;
        RECT 29.065 186.895 29.275 188.035 ;
        RECT 29.945 186.895 30.175 188.035 ;
        RECT 30.845 187.985 32.535 188.505 ;
        RECT 30.845 186.895 34.355 187.985 ;
        RECT 34.565 186.895 34.795 188.035 ;
        RECT 35.465 186.895 35.675 188.035 ;
        RECT 36.345 186.895 36.675 187.655 ;
        RECT 37.285 186.895 37.575 188.060 ;
        RECT 38.175 186.895 38.505 187.395 ;
        RECT 39.115 186.895 39.445 187.395 ;
        RECT 41.090 186.895 41.470 187.275 ;
        RECT 41.990 186.895 42.320 187.275 ;
        RECT 43.600 186.895 44.020 187.275 ;
        RECT 44.690 186.895 45.020 187.585 ;
        RECT 46.140 186.895 46.425 187.695 ;
        RECT 48.155 186.895 48.325 187.655 ;
        RECT 50.695 186.895 50.865 188.035 ;
        RECT 55.685 187.985 56.435 188.505 ;
        RECT 52.115 186.895 52.385 187.355 ;
        RECT 54.175 186.895 54.500 187.355 ;
        RECT 55.685 186.895 57.355 187.985 ;
        RECT 59.120 187.330 59.470 188.580 ;
        RECT 57.530 186.895 62.875 187.330 ;
        RECT 63.045 186.895 63.335 188.060 ;
        RECT 63.505 187.985 64.025 188.525 ;
        RECT 64.885 187.985 66.575 188.505 ;
        RECT 72.245 187.985 72.765 188.525 ;
        RECT 63.505 186.895 64.715 187.985 ;
        RECT 64.885 186.895 68.395 187.985 ;
        RECT 69.135 186.895 69.405 187.355 ;
        RECT 71.195 186.895 71.520 187.355 ;
        RECT 72.245 186.895 73.455 187.985 ;
        RECT 75.220 187.330 75.570 188.580 ;
        RECT 73.630 186.895 78.975 187.330 ;
        RECT 79.955 186.895 80.240 187.695 ;
        RECT 81.360 186.895 81.690 187.585 ;
        RECT 82.360 186.895 82.780 187.275 ;
        RECT 84.060 186.895 84.390 187.275 ;
        RECT 84.910 186.895 85.290 187.275 ;
        RECT 86.935 186.895 87.265 187.395 ;
        RECT 87.875 186.895 88.205 187.395 ;
        RECT 88.805 186.895 89.095 188.060 ;
        RECT 89.325 186.895 89.535 188.035 ;
        RECT 90.205 186.895 90.435 188.035 ;
        RECT 92.025 187.985 93.235 188.505 ;
        RECT 91.085 186.895 91.415 187.655 ;
        RECT 92.025 186.895 94.615 187.985 ;
        RECT 95.355 186.895 95.625 187.355 ;
        RECT 97.415 186.895 97.740 187.355 ;
        RECT 98.895 186.895 99.200 188.035 ;
        RECT 99.540 186.895 99.870 187.275 ;
        RECT 100.390 186.895 100.640 187.355 ;
        RECT 102.255 186.895 102.625 187.355 ;
        RECT 103.260 186.895 103.590 187.325 ;
        RECT 105.480 186.895 105.730 187.355 ;
        RECT 106.735 186.895 107.065 187.395 ;
        RECT 109.260 187.330 109.610 188.580 ;
        RECT 107.670 186.895 113.015 187.330 ;
        RECT 113.625 186.895 113.955 187.655 ;
        RECT 114.565 186.895 114.855 188.060 ;
        RECT 117.325 187.985 119.015 188.505 ;
        RECT 116.385 186.895 116.715 187.655 ;
        RECT 117.325 186.895 120.835 187.985 ;
        RECT 122.600 187.330 122.950 188.580 ;
        RECT 126.525 187.985 127.045 188.525 ;
        RECT 121.010 186.895 126.355 187.330 ;
        RECT 126.525 186.895 127.735 187.985 ;
        RECT 14.660 186.725 127.820 186.895 ;
        RECT 14.745 185.635 15.955 186.725 ;
        RECT 15.435 185.095 15.955 185.635 ;
        RECT 16.125 185.635 18.715 186.725 ;
        RECT 18.890 186.290 24.235 186.725 ;
        RECT 16.125 185.115 17.335 185.635 ;
        RECT 20.480 185.040 20.830 186.290 ;
        RECT 24.405 185.560 24.695 186.725 ;
        RECT 26.215 186.225 26.545 186.725 ;
        RECT 27.550 186.265 27.800 186.725 ;
        RECT 29.690 186.295 30.020 186.725 ;
        RECT 30.655 186.265 31.025 186.725 ;
        RECT 32.640 186.265 32.890 186.725 ;
        RECT 33.410 186.345 33.740 186.725 ;
        RECT 34.080 185.585 34.385 186.725 ;
        RECT 34.985 185.635 37.575 186.725 ;
        RECT 34.985 185.115 36.195 185.635 ;
        RECT 37.785 185.585 38.015 186.725 ;
        RECT 38.685 185.585 38.895 186.725 ;
        RECT 39.635 185.585 39.805 186.725 ;
        RECT 42.175 185.965 42.345 186.725 ;
        RECT 44.695 185.585 44.865 186.725 ;
        RECT 47.235 185.965 47.405 186.725 ;
        RECT 48.845 185.585 49.055 186.725 ;
        RECT 49.725 185.585 49.955 186.725 ;
        RECT 50.165 185.560 50.455 186.725 ;
        RECT 51.055 185.585 51.360 186.725 ;
        RECT 51.700 186.345 52.030 186.725 ;
        RECT 52.550 186.265 52.800 186.725 ;
        RECT 54.415 186.265 54.785 186.725 ;
        RECT 55.420 186.295 55.750 186.725 ;
        RECT 57.640 186.265 57.890 186.725 ;
        RECT 58.895 186.225 59.225 186.725 ;
        RECT 59.825 185.635 61.035 186.725 ;
        RECT 61.205 185.635 64.715 186.725 ;
        RECT 64.890 186.290 70.235 186.725 ;
        RECT 70.410 186.290 75.755 186.725 ;
        RECT 59.825 185.095 60.345 185.635 ;
        RECT 61.205 185.115 62.895 185.635 ;
        RECT 66.480 185.040 66.830 186.290 ;
        RECT 72.000 185.040 72.350 186.290 ;
        RECT 75.925 185.560 76.215 186.725 ;
        RECT 76.845 185.635 79.435 186.725 ;
        RECT 80.175 186.265 80.445 186.725 ;
        RECT 82.235 186.265 82.560 186.725 ;
        RECT 83.285 185.635 84.955 186.725 ;
        RECT 85.875 185.965 86.045 186.725 ;
        RECT 76.845 185.115 78.055 185.635 ;
        RECT 83.285 185.115 84.035 185.635 ;
        RECT 88.415 185.585 88.585 186.725 ;
        RECT 89.325 185.585 89.535 186.725 ;
        RECT 90.205 185.585 90.435 186.725 ;
        RECT 90.645 185.635 92.315 186.725 ;
        RECT 93.055 186.265 93.325 186.725 ;
        RECT 95.115 186.265 95.440 186.725 ;
        RECT 96.915 185.965 97.085 186.725 ;
        RECT 90.645 185.115 91.395 185.635 ;
        RECT 99.455 185.585 99.625 186.725 ;
        RECT 100.745 185.965 101.075 186.725 ;
        RECT 101.685 185.560 101.975 186.725 ;
        RECT 102.205 185.585 102.415 186.725 ;
        RECT 103.085 185.585 103.315 186.725 ;
        RECT 103.985 185.635 107.495 186.725 ;
        RECT 108.235 186.265 108.505 186.725 ;
        RECT 110.295 186.265 110.620 186.725 ;
        RECT 111.805 185.635 115.315 186.725 ;
        RECT 115.490 186.290 120.835 186.725 ;
        RECT 121.010 186.290 126.355 186.725 ;
        RECT 103.985 185.115 105.675 185.635 ;
        RECT 111.805 185.115 113.495 185.635 ;
        RECT 117.080 185.040 117.430 186.290 ;
        RECT 122.600 185.040 122.950 186.290 ;
        RECT 126.525 185.635 127.735 186.725 ;
        RECT 126.525 185.095 127.045 185.635 ;
        RECT 15.435 182.545 15.955 183.085 ;
        RECT 14.745 181.455 15.955 182.545 ;
        RECT 18.180 181.890 18.530 183.140 ;
        RECT 16.590 181.455 21.935 181.890 ;
        RECT 22.545 181.455 22.875 182.215 ;
        RECT 24.040 181.455 24.365 181.915 ;
        RECT 26.155 181.455 26.425 181.915 ;
        RECT 27.735 181.455 28.005 181.915 ;
        RECT 29.795 181.455 30.120 181.915 ;
        RECT 31.355 181.455 31.525 182.595 ;
        RECT 35.445 182.545 36.195 183.065 ;
        RECT 33.895 181.455 34.065 182.215 ;
        RECT 35.445 181.455 37.115 182.545 ;
        RECT 37.285 181.455 37.575 182.620 ;
        RECT 38.315 181.455 38.585 181.915 ;
        RECT 40.375 181.455 40.700 181.915 ;
        RECT 42.325 181.455 42.655 182.215 ;
        RECT 43.835 181.455 44.105 181.915 ;
        RECT 45.895 181.455 46.220 181.915 ;
        RECT 47.515 181.455 47.785 181.915 ;
        RECT 49.575 181.455 49.900 181.915 ;
        RECT 51.135 181.455 51.305 182.595 ;
        RECT 53.675 181.455 53.845 182.215 ;
        RECT 55.265 181.455 55.495 182.595 ;
        RECT 56.165 181.455 56.375 182.595 ;
        RECT 57.175 181.455 57.445 181.915 ;
        RECT 59.235 181.455 59.560 181.915 ;
        RECT 60.725 181.455 61.055 182.215 ;
        RECT 62.105 181.455 62.435 182.215 ;
        RECT 63.045 181.455 63.335 182.620 ;
        RECT 63.965 182.545 65.175 183.065 ;
        RECT 63.965 181.455 66.555 182.545 ;
        RECT 68.320 181.890 68.670 183.140 ;
        RECT 66.730 181.455 72.075 181.890 ;
        RECT 74.255 181.455 74.585 181.905 ;
        RECT 76.630 181.455 76.960 182.255 ;
        RECT 78.235 181.455 78.485 182.255 ;
        RECT 78.755 181.455 78.925 182.595 ;
        RECT 80.035 181.455 80.340 182.595 ;
        RECT 80.680 181.455 81.010 181.835 ;
        RECT 81.530 181.455 81.780 181.915 ;
        RECT 83.395 181.455 83.765 181.915 ;
        RECT 84.400 181.455 84.730 181.885 ;
        RECT 86.620 181.455 86.870 181.915 ;
        RECT 87.875 181.455 88.205 181.955 ;
        RECT 88.805 181.455 89.095 182.620 ;
        RECT 90.625 181.455 90.955 182.215 ;
        RECT 92.915 181.455 93.220 182.595 ;
        RECT 93.560 181.455 93.890 181.835 ;
        RECT 94.410 181.455 94.660 181.915 ;
        RECT 96.275 181.455 96.645 181.915 ;
        RECT 97.280 181.455 97.610 181.885 ;
        RECT 99.500 181.455 99.750 181.915 ;
        RECT 100.755 181.455 101.085 181.955 ;
        RECT 103.115 181.455 103.285 182.595 ;
        RECT 105.655 181.455 105.825 182.215 ;
        RECT 107.300 181.455 107.625 181.915 ;
        RECT 109.415 181.455 109.685 181.915 ;
        RECT 111.175 181.455 111.345 182.215 ;
        RECT 113.715 181.455 113.885 182.595 ;
        RECT 114.565 181.455 114.855 182.620 ;
        RECT 115.915 181.455 116.220 182.595 ;
        RECT 124.685 182.545 125.435 183.065 ;
        RECT 126.525 182.545 127.045 183.085 ;
        RECT 116.560 181.455 116.890 181.835 ;
        RECT 117.410 181.455 117.660 181.915 ;
        RECT 119.275 181.455 119.645 181.915 ;
        RECT 120.280 181.455 120.610 181.885 ;
        RECT 122.500 181.455 122.750 181.915 ;
        RECT 123.755 181.455 124.085 181.955 ;
        RECT 124.685 181.455 126.355 182.545 ;
        RECT 126.525 181.455 127.735 182.545 ;
        RECT 14.660 181.285 127.820 181.455 ;
        RECT 14.745 180.195 15.955 181.285 ;
        RECT 15.435 179.655 15.955 180.195 ;
        RECT 16.125 180.195 18.715 181.285 ;
        RECT 18.890 180.850 24.235 181.285 ;
        RECT 16.125 179.675 17.335 180.195 ;
        RECT 20.480 179.600 20.830 180.850 ;
        RECT 24.405 180.120 24.695 181.285 ;
        RECT 25.295 180.785 25.625 181.285 ;
        RECT 26.630 180.825 26.880 181.285 ;
        RECT 28.770 180.855 29.100 181.285 ;
        RECT 29.735 180.825 30.105 181.285 ;
        RECT 31.720 180.825 31.970 181.285 ;
        RECT 32.490 180.905 32.820 181.285 ;
        RECT 33.160 180.145 33.465 181.285 ;
        RECT 35.095 180.825 35.365 181.285 ;
        RECT 37.155 180.825 37.480 181.285 ;
        RECT 39.105 180.525 39.435 181.285 ;
        RECT 40.970 180.850 46.315 181.285 ;
        RECT 42.560 179.600 42.910 180.850 ;
        RECT 47.055 180.825 47.325 181.285 ;
        RECT 49.115 180.825 49.440 181.285 ;
        RECT 50.165 180.120 50.455 181.285 ;
        RECT 52.115 180.825 52.385 181.285 ;
        RECT 54.175 180.825 54.500 181.285 ;
        RECT 55.655 180.145 55.960 181.285 ;
        RECT 56.300 180.905 56.630 181.285 ;
        RECT 57.150 180.825 57.400 181.285 ;
        RECT 59.015 180.825 59.385 181.285 ;
        RECT 60.020 180.855 60.350 181.285 ;
        RECT 62.240 180.825 62.490 181.285 ;
        RECT 63.495 180.785 63.825 181.285 ;
        RECT 64.945 180.145 65.155 181.285 ;
        RECT 65.825 180.145 66.055 181.285 ;
        RECT 66.270 180.135 66.530 181.285 ;
        RECT 67.130 180.525 67.460 181.285 ;
        RECT 70.115 180.835 70.445 181.285 ;
        RECT 71.755 180.905 72.085 181.285 ;
        RECT 72.940 180.905 73.270 181.285 ;
        RECT 73.845 180.905 74.175 181.285 ;
        RECT 74.855 180.905 75.185 181.285 ;
        RECT 75.925 180.120 76.215 181.285 ;
        RECT 78.395 180.835 78.725 181.285 ;
        RECT 80.355 180.525 80.525 181.285 ;
        RECT 82.895 180.145 83.065 181.285 ;
        RECT 83.755 180.475 84.050 181.285 ;
        RECT 84.650 180.475 84.910 181.285 ;
        RECT 85.510 181.280 91.785 181.285 ;
        RECT 85.510 180.485 85.770 181.280 ;
        RECT 86.370 180.555 86.630 181.280 ;
        RECT 87.230 180.555 87.490 181.280 ;
        RECT 88.090 180.555 88.350 181.280 ;
        RECT 88.950 180.555 89.195 181.280 ;
        RECT 89.810 180.555 90.055 181.280 ;
        RECT 90.670 180.555 90.915 181.280 ;
        RECT 91.530 180.555 91.785 181.280 ;
        RECT 92.415 180.540 92.685 181.285 ;
        RECT 92.945 180.195 94.155 181.285 ;
        RECT 94.895 180.825 95.165 181.285 ;
        RECT 96.955 180.825 97.280 181.285 ;
        RECT 98.575 180.825 98.845 181.285 ;
        RECT 100.635 180.825 100.960 181.285 ;
        RECT 92.945 179.655 93.465 180.195 ;
        RECT 101.685 180.120 101.975 181.285 ;
        RECT 102.585 180.525 102.915 181.285 ;
        RECT 104.495 180.145 104.665 181.285 ;
        RECT 104.935 180.485 105.185 181.285 ;
        RECT 106.460 180.485 106.790 181.285 ;
        RECT 108.415 180.525 108.585 181.285 ;
        RECT 110.955 180.145 111.125 181.285 ;
        RECT 112.235 180.145 112.540 181.285 ;
        RECT 112.880 180.905 113.210 181.285 ;
        RECT 113.730 180.825 113.980 181.285 ;
        RECT 115.595 180.825 115.965 181.285 ;
        RECT 116.600 180.855 116.930 181.285 ;
        RECT 118.820 180.825 119.070 181.285 ;
        RECT 120.075 180.785 120.405 181.285 ;
        RECT 121.445 180.525 121.775 181.285 ;
        RECT 122.825 180.525 123.155 181.285 ;
        RECT 123.765 180.195 126.355 181.285 ;
        RECT 126.525 180.195 127.735 181.285 ;
        RECT 123.765 179.675 124.975 180.195 ;
        RECT 126.525 179.655 127.045 180.195 ;
        RECT 15.435 177.105 15.955 177.645 ;
        RECT 14.745 176.015 15.955 177.105 ;
        RECT 16.125 177.105 17.815 177.625 ;
        RECT 16.125 176.015 19.635 177.105 ;
        RECT 21.400 176.450 21.750 177.700 ;
        RECT 19.810 176.015 25.155 176.450 ;
        RECT 25.385 176.015 25.595 177.155 ;
        RECT 26.265 176.015 26.495 177.155 ;
        RECT 27.145 176.015 27.475 176.775 ;
        RECT 28.515 176.015 28.820 177.155 ;
        RECT 29.160 176.015 29.490 176.395 ;
        RECT 30.010 176.015 30.260 176.475 ;
        RECT 31.875 176.015 32.245 176.475 ;
        RECT 32.880 176.015 33.210 176.445 ;
        RECT 35.100 176.015 35.350 176.475 ;
        RECT 36.355 176.015 36.685 176.515 ;
        RECT 37.285 176.015 37.575 177.180 ;
        RECT 38.255 176.015 38.425 177.155 ;
        RECT 41.885 177.105 42.635 177.625 ;
        RECT 40.795 176.015 40.965 176.775 ;
        RECT 41.885 176.015 43.555 177.105 ;
        RECT 44.430 176.015 44.760 176.815 ;
        RECT 46.035 176.015 46.285 176.815 ;
        RECT 46.555 176.015 46.725 177.155 ;
        RECT 48.375 176.015 48.545 177.155 ;
        RECT 48.815 176.015 49.065 176.815 ;
        RECT 50.340 176.015 50.670 176.815 ;
        RECT 52.055 176.015 52.225 177.155 ;
        RECT 52.495 176.015 52.745 176.815 ;
        RECT 54.020 176.015 54.350 176.815 ;
        RECT 56.435 176.015 56.605 176.775 ;
        RECT 58.975 176.015 59.145 177.155 ;
        RECT 60.340 176.015 60.625 176.885 ;
        RECT 61.230 176.015 61.485 176.475 ;
        RECT 62.085 176.015 62.395 176.815 ;
        RECT 63.045 176.015 63.335 177.180 ;
        RECT 63.970 176.015 64.230 177.165 ;
        RECT 64.830 176.015 65.160 176.775 ;
        RECT 65.810 176.015 66.070 177.165 ;
        RECT 66.670 176.015 67.000 176.775 ;
        RECT 68.115 176.015 68.445 177.075 ;
        RECT 69.465 176.015 69.795 176.375 ;
        RECT 72.875 176.015 73.205 176.465 ;
        RECT 74.790 176.015 75.120 176.815 ;
        RECT 76.395 176.015 76.645 176.815 ;
        RECT 76.915 176.015 77.085 177.155 ;
        RECT 77.875 176.015 78.045 176.815 ;
        RECT 78.715 176.015 78.885 176.815 ;
        RECT 79.555 176.015 79.725 176.815 ;
        RECT 80.395 176.015 80.565 176.815 ;
        RECT 81.235 176.015 81.405 176.815 ;
        RECT 82.075 176.015 82.245 176.815 ;
        RECT 82.915 176.015 83.085 176.815 ;
        RECT 83.755 176.015 83.925 176.815 ;
        RECT 84.595 176.015 84.765 176.815 ;
        RECT 85.435 176.015 85.605 176.815 ;
        RECT 86.275 176.015 86.445 176.815 ;
        RECT 87.115 176.015 87.285 176.865 ;
        RECT 87.955 176.015 88.125 176.865 ;
        RECT 88.805 176.015 89.095 177.180 ;
        RECT 91.780 176.450 92.130 177.700 ;
        RECT 90.190 176.015 95.535 176.450 ;
        RECT 95.765 176.015 95.975 177.155 ;
        RECT 96.645 176.015 96.875 177.155 ;
        RECT 97.085 177.105 97.835 177.625 ;
        RECT 97.085 176.015 98.755 177.105 ;
        RECT 99.435 176.015 99.605 177.155 ;
        RECT 102.605 177.105 103.815 177.625 ;
        RECT 99.875 176.015 100.125 176.815 ;
        RECT 101.400 176.015 101.730 176.815 ;
        RECT 102.605 176.015 105.195 177.105 ;
        RECT 105.875 176.015 106.045 177.155 ;
        RECT 106.315 176.015 106.565 176.815 ;
        RECT 107.840 176.015 108.170 176.815 ;
        RECT 109.600 176.015 109.925 176.475 ;
        RECT 111.715 176.015 111.985 176.475 ;
        RECT 113.225 176.015 113.455 177.155 ;
        RECT 114.125 176.015 114.335 177.155 ;
        RECT 114.565 176.015 114.855 177.180 ;
        RECT 115.025 177.105 115.775 177.625 ;
        RECT 115.025 176.015 116.695 177.105 ;
        RECT 116.905 176.015 117.135 177.155 ;
        RECT 117.805 176.015 118.015 177.155 ;
        RECT 118.245 177.105 119.455 177.625 ;
        RECT 118.245 176.015 120.835 177.105 ;
        RECT 122.600 176.450 122.950 177.700 ;
        RECT 126.525 177.105 127.045 177.645 ;
        RECT 121.010 176.015 126.355 176.450 ;
        RECT 126.525 176.015 127.735 177.105 ;
        RECT 14.660 175.845 127.820 176.015 ;
        RECT 14.745 174.755 15.955 175.845 ;
        RECT 15.435 174.215 15.955 174.755 ;
        RECT 16.125 174.755 18.715 175.845 ;
        RECT 18.890 175.410 24.235 175.845 ;
        RECT 16.125 174.235 17.335 174.755 ;
        RECT 20.480 174.160 20.830 175.410 ;
        RECT 24.405 174.680 24.695 175.845 ;
        RECT 25.845 174.705 26.055 175.845 ;
        RECT 26.725 174.705 26.955 175.845 ;
        RECT 27.735 175.385 28.005 175.845 ;
        RECT 29.795 175.385 30.120 175.845 ;
        RECT 31.815 174.705 31.985 175.845 ;
        RECT 34.355 175.085 34.525 175.845 ;
        RECT 36.150 175.045 36.480 175.845 ;
        RECT 37.755 175.045 38.005 175.845 ;
        RECT 38.275 174.705 38.445 175.845 ;
        RECT 39.635 174.705 39.805 175.845 ;
        RECT 40.075 175.045 40.325 175.845 ;
        RECT 41.600 175.045 41.930 175.845 ;
        RECT 43.510 175.045 43.840 175.845 ;
        RECT 45.115 175.045 45.365 175.845 ;
        RECT 45.635 174.705 45.805 175.845 ;
        RECT 46.995 174.705 47.165 175.845 ;
        RECT 47.435 175.045 47.685 175.845 ;
        RECT 48.960 175.045 49.290 175.845 ;
        RECT 50.165 174.680 50.455 175.845 ;
        RECT 50.625 174.755 51.835 175.845 ;
        RECT 52.575 175.385 52.845 175.845 ;
        RECT 54.635 175.385 54.960 175.845 ;
        RECT 57.355 175.085 57.525 175.845 ;
        RECT 50.625 174.215 51.145 174.755 ;
        RECT 59.895 174.705 60.065 175.845 ;
        RECT 60.745 174.755 62.415 175.845 ;
        RECT 63.025 175.085 63.355 175.845 ;
        RECT 64.425 174.755 67.935 175.845 ;
        RECT 68.615 175.045 68.855 175.845 ;
        RECT 69.375 175.045 69.705 175.845 ;
        RECT 60.745 174.235 61.495 174.755 ;
        RECT 64.425 174.235 66.115 174.755 ;
        RECT 70.215 174.695 70.545 175.845 ;
        RECT 71.330 174.695 71.590 175.845 ;
        RECT 72.190 175.085 72.520 175.845 ;
        RECT 73.640 175.085 73.970 175.845 ;
        RECT 74.570 174.695 74.830 175.845 ;
        RECT 75.925 174.680 76.215 175.845 ;
        RECT 78.010 175.045 78.340 175.845 ;
        RECT 79.615 175.045 79.865 175.845 ;
        RECT 80.135 174.705 80.305 175.845 ;
        RECT 81.495 174.705 81.665 175.845 ;
        RECT 81.935 175.045 82.185 175.845 ;
        RECT 83.460 175.045 83.790 175.845 ;
        RECT 85.220 175.385 85.545 175.845 ;
        RECT 87.335 175.385 87.605 175.845 ;
        RECT 88.825 175.045 89.135 175.845 ;
        RECT 89.735 175.385 89.990 175.845 ;
        RECT 90.595 174.975 90.880 175.845 ;
        RECT 91.105 174.755 92.315 175.845 ;
        RECT 92.485 174.755 95.995 175.845 ;
        RECT 96.170 175.410 101.515 175.845 ;
        RECT 91.105 174.215 91.625 174.755 ;
        RECT 92.485 174.235 94.175 174.755 ;
        RECT 97.760 174.160 98.110 175.410 ;
        RECT 101.685 174.680 101.975 175.845 ;
        RECT 102.155 175.035 102.450 175.845 ;
        RECT 103.050 175.035 103.310 175.845 ;
        RECT 103.910 175.840 110.185 175.845 ;
        RECT 103.910 175.045 104.170 175.840 ;
        RECT 104.770 175.115 105.030 175.840 ;
        RECT 105.630 175.115 105.890 175.840 ;
        RECT 106.490 175.115 106.750 175.840 ;
        RECT 107.350 175.115 107.595 175.840 ;
        RECT 108.210 175.115 108.455 175.840 ;
        RECT 109.070 175.115 109.315 175.840 ;
        RECT 109.930 175.115 110.185 175.840 ;
        RECT 110.815 175.100 111.085 175.845 ;
        RECT 111.855 174.705 112.025 175.845 ;
        RECT 112.295 175.045 112.545 175.845 ;
        RECT 113.820 175.045 114.150 175.845 ;
        RECT 115.730 175.045 116.060 175.845 ;
        RECT 117.335 175.045 117.585 175.845 ;
        RECT 117.855 174.705 118.025 175.845 ;
        RECT 118.765 174.705 118.975 175.845 ;
        RECT 119.645 174.705 119.875 175.845 ;
        RECT 121.010 175.410 126.355 175.845 ;
        RECT 122.600 174.160 122.950 175.410 ;
        RECT 126.525 174.755 127.735 175.845 ;
        RECT 126.525 174.215 127.045 174.755 ;
        RECT 15.435 171.665 15.955 172.205 ;
        RECT 14.745 170.575 15.955 171.665 ;
        RECT 18.640 171.010 18.990 172.260 ;
        RECT 24.160 171.010 24.510 172.260 ;
        RECT 29.680 171.010 30.030 172.260 ;
        RECT 17.050 170.575 22.395 171.010 ;
        RECT 22.570 170.575 27.915 171.010 ;
        RECT 28.090 170.575 33.435 171.010 ;
        RECT 34.310 170.575 34.640 171.375 ;
        RECT 35.915 170.575 36.165 171.375 ;
        RECT 36.435 170.575 36.605 171.715 ;
        RECT 37.285 170.575 37.575 171.740 ;
        RECT 38.715 170.575 38.885 171.715 ;
        RECT 41.885 171.665 43.095 172.185 ;
        RECT 39.155 170.575 39.405 171.375 ;
        RECT 40.680 170.575 41.010 171.375 ;
        RECT 41.885 170.575 44.475 171.665 ;
        RECT 44.735 170.575 45.005 171.320 ;
        RECT 45.635 170.580 45.890 171.305 ;
        RECT 46.505 170.580 46.750 171.305 ;
        RECT 47.365 170.580 47.610 171.305 ;
        RECT 48.225 170.580 48.470 171.305 ;
        RECT 49.070 170.580 49.330 171.305 ;
        RECT 49.930 170.580 50.190 171.305 ;
        RECT 50.790 170.580 51.050 171.305 ;
        RECT 51.650 170.580 51.910 171.375 ;
        RECT 45.635 170.575 51.910 170.580 ;
        RECT 52.510 170.575 52.770 171.385 ;
        RECT 53.370 170.575 53.665 171.385 ;
        RECT 54.275 170.575 54.580 171.715 ;
        RECT 54.920 170.575 55.250 170.955 ;
        RECT 55.770 170.575 56.020 171.035 ;
        RECT 57.635 170.575 58.005 171.035 ;
        RECT 58.640 170.575 58.970 171.005 ;
        RECT 60.860 170.575 61.110 171.035 ;
        RECT 62.115 170.575 62.445 171.075 ;
        RECT 63.045 170.575 63.335 171.740 ;
        RECT 63.565 170.575 63.775 171.715 ;
        RECT 64.445 170.575 64.675 171.715 ;
        RECT 67.400 171.010 67.750 172.260 ;
        RECT 72.920 171.010 73.270 172.260 ;
        RECT 78.440 171.010 78.790 172.260 ;
        RECT 65.810 170.575 71.155 171.010 ;
        RECT 71.330 170.575 76.675 171.010 ;
        RECT 76.850 170.575 82.195 171.010 ;
        RECT 82.875 170.575 83.115 171.375 ;
        RECT 83.635 170.575 83.965 171.375 ;
        RECT 84.475 170.575 84.805 171.725 ;
        RECT 85.695 170.575 85.965 171.035 ;
        RECT 87.755 170.575 88.080 171.035 ;
        RECT 88.805 170.575 89.095 171.740 ;
        RECT 89.765 170.575 89.995 171.715 ;
        RECT 90.665 170.575 90.875 171.715 ;
        RECT 91.535 170.575 91.840 171.715 ;
        RECT 101.225 171.665 102.915 172.185 ;
        RECT 92.180 170.575 92.510 170.955 ;
        RECT 93.030 170.575 93.280 171.035 ;
        RECT 94.895 170.575 95.265 171.035 ;
        RECT 95.900 170.575 96.230 171.005 ;
        RECT 98.120 170.575 98.370 171.035 ;
        RECT 99.375 170.575 99.705 171.075 ;
        RECT 101.225 170.575 104.735 171.665 ;
        RECT 104.905 170.575 105.290 171.410 ;
        RECT 105.890 170.575 106.150 171.410 ;
        RECT 106.750 170.575 107.010 171.410 ;
        RECT 107.610 170.575 107.955 171.410 ;
        RECT 108.635 170.575 108.805 171.715 ;
        RECT 111.805 171.665 112.325 172.205 ;
        RECT 109.075 170.575 109.325 171.375 ;
        RECT 110.600 170.575 110.930 171.375 ;
        RECT 111.805 170.575 113.015 171.665 ;
        RECT 113.225 170.575 113.455 171.715 ;
        RECT 114.125 170.575 114.335 171.715 ;
        RECT 114.565 170.575 114.855 171.740 ;
        RECT 116.375 170.575 116.680 171.715 ;
        RECT 125.145 171.665 125.665 172.205 ;
        RECT 126.525 171.665 127.045 172.205 ;
        RECT 117.020 170.575 117.350 170.955 ;
        RECT 117.870 170.575 118.120 171.035 ;
        RECT 119.735 170.575 120.105 171.035 ;
        RECT 120.740 170.575 121.070 171.005 ;
        RECT 122.960 170.575 123.210 171.035 ;
        RECT 124.215 170.575 124.545 171.075 ;
        RECT 125.145 170.575 126.355 171.665 ;
        RECT 126.525 170.575 127.735 171.665 ;
        RECT 14.660 170.405 127.820 170.575 ;
        RECT 14.745 169.315 15.955 170.405 ;
        RECT 15.435 168.775 15.955 169.315 ;
        RECT 16.125 169.315 18.715 170.405 ;
        RECT 18.890 169.970 24.235 170.405 ;
        RECT 16.125 168.795 17.335 169.315 ;
        RECT 20.480 168.720 20.830 169.970 ;
        RECT 24.405 169.240 24.695 170.405 ;
        RECT 25.325 169.315 26.995 170.405 ;
        RECT 25.325 168.795 26.075 169.315 ;
        RECT 27.225 169.265 27.435 170.405 ;
        RECT 28.105 169.265 28.335 170.405 ;
        RECT 28.545 169.315 30.215 170.405 ;
        RECT 28.545 168.795 29.295 169.315 ;
        RECT 30.445 169.265 30.655 170.405 ;
        RECT 31.325 169.265 31.555 170.405 ;
        RECT 32.335 169.945 32.605 170.405 ;
        RECT 34.395 169.945 34.720 170.405 ;
        RECT 35.575 169.235 35.905 170.405 ;
        RECT 36.635 169.235 36.965 170.405 ;
        RECT 37.695 169.265 38.025 170.405 ;
        RECT 38.205 169.315 39.875 170.405 ;
        RECT 40.050 169.970 45.395 170.405 ;
        RECT 38.205 168.795 38.955 169.315 ;
        RECT 41.640 168.720 41.990 169.970 ;
        RECT 46.075 169.265 46.245 170.405 ;
        RECT 46.515 169.605 46.765 170.405 ;
        RECT 48.040 169.605 48.370 170.405 ;
        RECT 50.165 169.240 50.455 170.405 ;
        RECT 50.625 169.315 52.295 170.405 ;
        RECT 52.465 169.570 52.850 170.405 ;
        RECT 53.450 169.570 53.710 170.405 ;
        RECT 54.310 169.570 54.570 170.405 ;
        RECT 55.170 169.570 55.515 170.405 ;
        RECT 55.685 169.315 57.355 170.405 ;
        RECT 57.530 169.970 62.875 170.405 ;
        RECT 63.050 169.970 68.395 170.405 ;
        RECT 50.625 168.795 51.375 169.315 ;
        RECT 55.685 168.795 56.435 169.315 ;
        RECT 59.120 168.720 59.470 169.970 ;
        RECT 64.640 168.720 64.990 169.970 ;
        RECT 69.040 169.645 69.370 170.405 ;
        RECT 69.970 169.255 70.230 170.405 ;
        RECT 70.410 169.255 70.670 170.405 ;
        RECT 71.270 169.645 71.600 170.405 ;
        RECT 73.185 169.605 73.495 170.405 ;
        RECT 74.095 169.945 74.350 170.405 ;
        RECT 74.955 169.535 75.240 170.405 ;
        RECT 75.925 169.240 76.215 170.405 ;
        RECT 77.135 169.645 77.305 170.405 ;
        RECT 79.675 169.265 79.845 170.405 ;
        RECT 81.335 169.605 81.620 170.405 ;
        RECT 82.740 169.715 83.070 170.405 ;
        RECT 83.740 170.025 84.160 170.405 ;
        RECT 85.440 170.025 85.770 170.405 ;
        RECT 86.290 170.025 86.670 170.405 ;
        RECT 88.315 169.905 88.645 170.405 ;
        RECT 89.255 169.905 89.585 170.405 ;
        RECT 91.855 169.645 92.025 170.405 ;
        RECT 94.395 169.265 94.565 170.405 ;
        RECT 96.605 169.645 96.935 170.405 ;
        RECT 98.005 169.315 101.515 170.405 ;
        RECT 98.005 168.795 99.695 169.315 ;
        RECT 101.685 169.240 101.975 170.405 ;
        RECT 103.035 169.265 103.340 170.405 ;
        RECT 103.680 170.025 104.010 170.405 ;
        RECT 104.530 169.945 104.780 170.405 ;
        RECT 106.395 169.945 106.765 170.405 ;
        RECT 107.400 169.975 107.730 170.405 ;
        RECT 109.620 169.945 109.870 170.405 ;
        RECT 110.875 169.905 111.205 170.405 ;
        RECT 113.235 169.265 113.405 170.405 ;
        RECT 115.775 169.645 115.945 170.405 ;
        RECT 117.420 169.945 117.745 170.405 ;
        RECT 119.535 169.945 119.805 170.405 ;
        RECT 120.585 169.265 120.815 170.405 ;
        RECT 121.485 169.265 121.695 170.405 ;
        RECT 121.930 169.980 122.265 170.405 ;
        RECT 122.825 169.625 123.155 170.405 ;
        RECT 124.205 169.645 124.535 170.405 ;
        RECT 125.145 169.315 126.355 170.405 ;
        RECT 126.525 169.315 127.735 170.405 ;
        RECT 125.145 168.775 125.665 169.315 ;
        RECT 126.525 168.775 127.045 169.315 ;
        RECT 15.435 166.225 15.955 166.765 ;
        RECT 14.745 165.135 15.955 166.225 ;
        RECT 16.585 166.225 17.335 166.745 ;
        RECT 16.585 165.135 18.255 166.225 ;
        RECT 18.855 165.135 19.160 166.275 ;
        RECT 19.500 165.135 19.830 165.515 ;
        RECT 20.350 165.135 20.600 165.595 ;
        RECT 22.215 165.135 22.585 165.595 ;
        RECT 23.220 165.135 23.550 165.565 ;
        RECT 25.440 165.135 25.690 165.595 ;
        RECT 26.695 165.135 27.025 165.635 ;
        RECT 27.715 165.135 27.985 165.880 ;
        RECT 28.615 165.140 28.870 165.865 ;
        RECT 29.485 165.140 29.730 165.865 ;
        RECT 30.345 165.140 30.590 165.865 ;
        RECT 31.205 165.140 31.450 165.865 ;
        RECT 32.050 165.140 32.310 165.865 ;
        RECT 32.910 165.140 33.170 165.865 ;
        RECT 33.770 165.140 34.030 165.865 ;
        RECT 34.630 165.140 34.890 165.935 ;
        RECT 28.615 165.135 34.890 165.140 ;
        RECT 35.490 165.135 35.750 165.945 ;
        RECT 36.350 165.135 36.645 165.945 ;
        RECT 37.285 165.135 37.575 166.300 ;
        RECT 38.185 165.135 38.515 165.895 ;
        RECT 39.185 165.135 39.395 166.275 ;
        RECT 40.065 165.135 40.295 166.275 ;
        RECT 41.405 165.135 41.735 165.895 ;
        RECT 42.385 165.135 42.615 166.275 ;
        RECT 43.285 165.135 43.495 166.275 ;
        RECT 44.295 165.135 44.565 165.595 ;
        RECT 46.355 165.135 46.680 165.595 ;
        RECT 47.835 165.135 48.140 166.275 ;
        RECT 48.480 165.135 48.810 165.515 ;
        RECT 49.330 165.135 49.580 165.595 ;
        RECT 51.195 165.135 51.565 165.595 ;
        RECT 52.200 165.135 52.530 165.565 ;
        RECT 54.420 165.135 54.670 165.595 ;
        RECT 55.675 165.135 56.005 165.635 ;
        RECT 57.585 165.135 57.795 166.275 ;
        RECT 58.465 165.135 58.695 166.275 ;
        RECT 59.975 165.135 60.305 166.285 ;
        RECT 60.815 165.135 61.145 165.935 ;
        RECT 61.665 165.135 61.905 165.935 ;
        RECT 63.045 165.135 63.335 166.300 ;
        RECT 64.575 165.135 64.905 166.285 ;
        RECT 69.945 166.225 70.465 166.765 ;
        RECT 74.085 166.225 74.605 166.765 ;
        RECT 65.415 165.135 65.745 165.935 ;
        RECT 66.265 165.135 66.505 165.935 ;
        RECT 67.240 165.135 67.525 166.005 ;
        RECT 68.130 165.135 68.385 165.595 ;
        RECT 68.985 165.135 69.295 165.935 ;
        RECT 69.945 165.135 71.155 166.225 ;
        RECT 71.335 165.135 71.665 166.195 ;
        RECT 72.685 165.135 73.015 165.495 ;
        RECT 74.085 165.135 75.295 166.225 ;
        RECT 76.275 165.135 76.560 165.935 ;
        RECT 77.680 165.135 78.010 165.825 ;
        RECT 78.680 165.135 79.100 165.515 ;
        RECT 80.380 165.135 80.710 165.515 ;
        RECT 81.230 165.135 81.610 165.515 ;
        RECT 83.255 165.135 83.585 165.635 ;
        RECT 84.195 165.135 84.525 165.635 ;
        RECT 85.185 165.135 85.395 166.275 ;
        RECT 86.065 165.135 86.295 166.275 ;
        RECT 86.565 165.135 86.775 166.275 ;
        RECT 87.445 165.135 87.675 166.275 ;
        RECT 88.805 165.135 89.095 166.300 ;
        RECT 89.725 166.225 90.475 166.745 ;
        RECT 89.725 165.135 91.395 166.225 ;
        RECT 93.160 165.570 93.510 166.820 ;
        RECT 91.570 165.135 96.915 165.570 ;
        RECT 97.895 165.135 98.180 165.935 ;
        RECT 99.300 165.135 99.630 165.825 ;
        RECT 100.300 165.135 100.720 165.515 ;
        RECT 102.000 165.135 102.330 165.515 ;
        RECT 102.850 165.135 103.230 165.515 ;
        RECT 104.875 165.135 105.205 165.635 ;
        RECT 105.815 165.135 106.145 165.635 ;
        RECT 107.775 165.135 108.045 165.595 ;
        RECT 109.835 165.135 110.160 165.595 ;
        RECT 111.440 165.135 111.765 165.595 ;
        RECT 113.555 165.135 113.825 165.595 ;
        RECT 114.565 165.135 114.855 166.300 ;
        RECT 116.375 165.135 116.680 166.275 ;
        RECT 125.145 166.225 125.665 166.765 ;
        RECT 126.525 166.225 127.045 166.765 ;
        RECT 117.020 165.135 117.350 165.515 ;
        RECT 117.870 165.135 118.120 165.595 ;
        RECT 119.735 165.135 120.105 165.595 ;
        RECT 120.740 165.135 121.070 165.565 ;
        RECT 122.960 165.135 123.210 165.595 ;
        RECT 124.215 165.135 124.545 165.635 ;
        RECT 125.145 165.135 126.355 166.225 ;
        RECT 126.525 165.135 127.735 166.225 ;
        RECT 14.660 164.965 127.820 165.135 ;
        RECT 14.745 163.875 15.955 164.965 ;
        RECT 15.435 163.335 15.955 163.875 ;
        RECT 16.125 163.875 18.715 164.965 ;
        RECT 18.890 164.530 24.235 164.965 ;
        RECT 16.125 163.355 17.335 163.875 ;
        RECT 20.480 163.280 20.830 164.530 ;
        RECT 24.405 163.800 24.695 164.965 ;
        RECT 26.225 164.205 26.555 164.965 ;
        RECT 27.595 163.825 27.900 164.965 ;
        RECT 28.240 164.585 28.570 164.965 ;
        RECT 29.090 164.505 29.340 164.965 ;
        RECT 30.955 164.505 31.325 164.965 ;
        RECT 31.960 164.535 32.290 164.965 ;
        RECT 34.180 164.505 34.430 164.965 ;
        RECT 35.435 164.465 35.765 164.965 ;
        RECT 36.795 163.825 37.100 164.965 ;
        RECT 37.440 164.585 37.770 164.965 ;
        RECT 38.290 164.505 38.540 164.965 ;
        RECT 40.155 164.505 40.525 164.965 ;
        RECT 41.160 164.535 41.490 164.965 ;
        RECT 43.380 164.505 43.630 164.965 ;
        RECT 44.635 164.465 44.965 164.965 ;
        RECT 46.075 163.825 46.245 164.965 ;
        RECT 48.615 164.205 48.785 164.965 ;
        RECT 50.165 163.800 50.455 164.965 ;
        RECT 51.375 164.205 51.545 164.965 ;
        RECT 53.915 163.825 54.085 164.965 ;
        RECT 55.195 163.825 55.500 164.965 ;
        RECT 55.840 164.585 56.170 164.965 ;
        RECT 56.690 164.505 56.940 164.965 ;
        RECT 58.555 164.505 58.925 164.965 ;
        RECT 59.560 164.535 59.890 164.965 ;
        RECT 61.780 164.505 62.030 164.965 ;
        RECT 63.035 164.465 63.365 164.965 ;
        RECT 64.425 163.875 67.015 164.965 ;
        RECT 67.240 164.095 67.525 164.965 ;
        RECT 68.130 164.505 68.385 164.965 ;
        RECT 68.985 164.165 69.295 164.965 ;
        RECT 70.410 164.530 75.755 164.965 ;
        RECT 64.425 163.355 65.635 163.875 ;
        RECT 72.000 163.280 72.350 164.530 ;
        RECT 75.925 163.800 76.215 164.965 ;
        RECT 76.385 163.875 78.055 164.965 ;
        RECT 78.975 164.205 79.145 164.965 ;
        RECT 76.385 163.355 77.135 163.875 ;
        RECT 81.515 163.825 81.685 164.965 ;
        RECT 82.805 164.205 83.135 164.965 ;
        RECT 83.745 163.875 85.415 164.965 ;
        RECT 86.025 164.205 86.355 164.965 ;
        RECT 87.890 164.530 93.235 164.965 ;
        RECT 83.745 163.355 84.495 163.875 ;
        RECT 89.480 163.280 89.830 164.530 ;
        RECT 94.155 164.205 94.325 164.965 ;
        RECT 96.695 163.825 96.865 164.965 ;
        RECT 98.295 164.205 98.465 164.965 ;
        RECT 100.835 163.825 101.005 164.965 ;
        RECT 101.685 163.800 101.975 164.965 ;
        RECT 102.700 164.505 103.025 164.965 ;
        RECT 104.815 164.505 105.085 164.965 ;
        RECT 107.255 163.825 107.425 164.965 ;
        RECT 109.795 164.205 109.965 164.965 ;
        RECT 110.945 163.825 111.155 164.965 ;
        RECT 111.825 163.825 112.055 164.965 ;
        RECT 113.615 163.825 113.920 164.965 ;
        RECT 114.260 164.585 114.590 164.965 ;
        RECT 115.110 164.505 115.360 164.965 ;
        RECT 116.975 164.505 117.345 164.965 ;
        RECT 117.980 164.535 118.310 164.965 ;
        RECT 120.200 164.505 120.450 164.965 ;
        RECT 121.455 164.465 121.785 164.965 ;
        RECT 122.825 164.205 123.155 164.965 ;
        RECT 123.765 163.875 126.355 164.965 ;
        RECT 126.525 163.875 127.735 164.965 ;
        RECT 123.765 163.355 124.975 163.875 ;
        RECT 126.525 163.335 127.045 163.875 ;
        RECT 15.435 160.785 15.955 161.325 ;
        RECT 14.745 159.695 15.955 160.785 ;
        RECT 16.125 160.785 16.875 161.305 ;
        RECT 16.125 159.695 17.795 160.785 ;
        RECT 18.775 159.695 19.060 160.495 ;
        RECT 20.180 159.695 20.510 160.385 ;
        RECT 21.180 159.695 21.600 160.075 ;
        RECT 22.880 159.695 23.210 160.075 ;
        RECT 23.730 159.695 24.110 160.075 ;
        RECT 25.755 159.695 26.085 160.195 ;
        RECT 26.695 159.695 27.025 160.195 ;
        RECT 28.135 159.695 28.305 160.835 ;
        RECT 31.765 160.785 32.285 161.325 ;
        RECT 30.675 159.695 30.845 160.455 ;
        RECT 31.765 159.695 32.975 160.785 ;
        RECT 33.895 159.695 34.065 160.455 ;
        RECT 36.435 159.695 36.605 160.835 ;
        RECT 37.285 159.695 37.575 160.860 ;
        RECT 38.205 160.785 39.895 161.305 ;
        RECT 45.565 160.785 46.085 161.325 ;
        RECT 38.205 159.695 41.715 160.785 ;
        RECT 42.440 159.695 42.765 160.155 ;
        RECT 44.555 159.695 44.825 160.155 ;
        RECT 45.565 159.695 46.775 160.785 ;
        RECT 47.515 159.695 47.785 160.155 ;
        RECT 49.575 159.695 49.900 160.155 ;
        RECT 51.375 159.695 51.545 160.455 ;
        RECT 53.915 159.695 54.085 160.835 ;
        RECT 60.285 160.785 61.495 161.305 ;
        RECT 55.335 159.695 55.605 160.155 ;
        RECT 57.395 159.695 57.720 160.155 ;
        RECT 59.345 159.695 59.675 160.455 ;
        RECT 60.285 159.695 62.875 160.785 ;
        RECT 63.045 159.695 63.335 160.860 ;
        RECT 63.505 160.785 64.025 161.325 ;
        RECT 63.505 159.695 64.715 160.785 ;
        RECT 64.890 159.695 65.150 160.845 ;
        RECT 65.750 159.695 66.080 160.455 ;
        RECT 66.730 159.695 66.990 160.845 ;
        RECT 67.590 159.695 67.920 160.455 ;
        RECT 69.040 159.695 69.370 160.455 ;
        RECT 69.970 159.695 70.230 160.845 ;
        RECT 70.880 159.695 71.210 160.455 ;
        RECT 71.810 159.695 72.070 160.845 ;
        RECT 72.245 160.785 73.455 161.305 ;
        RECT 72.245 159.695 74.835 160.785 ;
        RECT 76.600 160.130 76.950 161.380 ;
        RECT 75.010 159.695 80.355 160.130 ;
        RECT 80.585 159.695 80.795 160.835 ;
        RECT 81.465 159.695 81.695 160.835 ;
        RECT 82.655 159.695 82.825 160.455 ;
        RECT 85.195 159.695 85.365 160.835 ;
        RECT 86.945 159.695 87.275 160.455 ;
        RECT 88.805 159.695 89.095 160.860 ;
        RECT 90.075 159.695 90.360 160.495 ;
        RECT 91.480 159.695 91.810 160.385 ;
        RECT 92.480 159.695 92.900 160.075 ;
        RECT 94.180 159.695 94.510 160.075 ;
        RECT 95.030 159.695 95.410 160.075 ;
        RECT 97.055 159.695 97.385 160.195 ;
        RECT 97.995 159.695 98.325 160.195 ;
        RECT 100.285 159.695 100.615 160.455 ;
        RECT 101.285 159.695 101.495 160.835 ;
        RECT 102.165 159.695 102.395 160.835 ;
        RECT 103.160 159.695 103.485 160.155 ;
        RECT 105.275 159.695 105.545 160.155 ;
        RECT 107.315 159.695 107.585 160.155 ;
        RECT 109.375 159.695 109.700 160.155 ;
        RECT 111.175 159.695 111.345 160.455 ;
        RECT 113.715 159.695 113.885 160.835 ;
        RECT 114.565 159.695 114.855 160.860 ;
        RECT 115.775 159.695 115.945 160.455 ;
        RECT 118.315 159.695 118.485 160.835 ;
        RECT 124.685 160.785 125.435 161.305 ;
        RECT 126.525 160.785 127.045 161.325 ;
        RECT 119.735 159.695 120.005 160.155 ;
        RECT 121.795 159.695 122.120 160.155 ;
        RECT 123.285 159.695 123.615 160.455 ;
        RECT 124.685 159.695 126.355 160.785 ;
        RECT 126.525 159.695 127.735 160.785 ;
        RECT 14.660 159.525 127.820 159.695 ;
        RECT 14.745 158.435 15.955 159.525 ;
        RECT 15.435 157.895 15.955 158.435 ;
        RECT 16.125 158.435 17.335 159.525 ;
        RECT 16.125 157.895 16.645 158.435 ;
        RECT 17.565 158.385 17.775 159.525 ;
        RECT 18.445 158.385 18.675 159.525 ;
        RECT 18.925 158.385 19.155 159.525 ;
        RECT 19.825 158.385 20.035 159.525 ;
        RECT 21.015 158.765 21.185 159.525 ;
        RECT 23.555 158.385 23.725 159.525 ;
        RECT 24.405 158.360 24.695 159.525 ;
        RECT 25.305 158.765 25.635 159.525 ;
        RECT 26.710 159.090 32.055 159.525 ;
        RECT 28.300 157.840 28.650 159.090 ;
        RECT 32.780 159.065 33.105 159.525 ;
        RECT 34.895 159.065 35.165 159.525 ;
        RECT 35.905 158.435 37.115 159.525 ;
        RECT 37.290 159.090 42.635 159.525 ;
        RECT 35.905 157.895 36.425 158.435 ;
        RECT 38.880 157.840 39.230 159.090 ;
        RECT 43.510 158.725 43.840 159.525 ;
        RECT 45.115 158.725 45.365 159.525 ;
        RECT 45.635 158.385 45.805 159.525 ;
        RECT 46.995 158.385 47.165 159.525 ;
        RECT 47.435 158.725 47.685 159.525 ;
        RECT 48.960 158.725 49.290 159.525 ;
        RECT 50.165 158.360 50.455 159.525 ;
        RECT 51.135 158.385 51.305 159.525 ;
        RECT 51.575 158.725 51.825 159.525 ;
        RECT 53.100 158.725 53.430 159.525 ;
        RECT 55.205 158.765 55.535 159.525 ;
        RECT 56.150 159.090 61.495 159.525 ;
        RECT 57.740 157.840 58.090 159.090 ;
        RECT 61.815 158.375 62.145 159.525 ;
        RECT 62.655 158.725 62.985 159.525 ;
        RECT 63.505 158.725 63.745 159.525 ;
        RECT 64.885 158.435 68.395 159.525 ;
        RECT 69.040 158.765 69.370 159.525 ;
        RECT 64.885 157.915 66.575 158.435 ;
        RECT 69.970 158.375 70.230 159.525 ;
        RECT 70.880 158.765 71.210 159.525 ;
        RECT 71.810 158.375 72.070 159.525 ;
        RECT 72.950 158.725 73.280 159.525 ;
        RECT 74.555 158.725 74.805 159.525 ;
        RECT 75.075 158.385 75.245 159.525 ;
        RECT 75.925 158.360 76.215 159.525 ;
        RECT 77.355 158.385 77.525 159.525 ;
        RECT 77.795 158.725 78.045 159.525 ;
        RECT 79.320 158.725 79.650 159.525 ;
        RECT 81.335 158.725 81.620 159.525 ;
        RECT 82.740 158.835 83.070 159.525 ;
        RECT 83.740 159.145 84.160 159.525 ;
        RECT 85.440 159.145 85.770 159.525 ;
        RECT 86.290 159.145 86.670 159.525 ;
        RECT 88.315 159.025 88.645 159.525 ;
        RECT 89.255 159.025 89.585 159.525 ;
        RECT 90.185 158.435 92.775 159.525 ;
        RECT 90.185 157.915 91.395 158.435 ;
        RECT 93.005 158.385 93.215 159.525 ;
        RECT 93.885 158.385 94.115 159.525 ;
        RECT 94.325 158.435 95.995 159.525 ;
        RECT 96.605 158.765 96.935 159.525 ;
        RECT 98.005 158.435 101.515 159.525 ;
        RECT 94.325 157.915 95.075 158.435 ;
        RECT 98.005 157.915 99.695 158.435 ;
        RECT 101.685 158.360 101.975 159.525 ;
        RECT 102.605 158.435 105.195 159.525 ;
        RECT 105.805 158.765 106.135 159.525 ;
        RECT 106.745 158.435 107.955 159.525 ;
        RECT 108.130 159.090 113.475 159.525 ;
        RECT 113.650 159.090 118.995 159.525 ;
        RECT 102.605 157.915 103.815 158.435 ;
        RECT 106.745 157.895 107.265 158.435 ;
        RECT 109.720 157.840 110.070 159.090 ;
        RECT 115.240 157.840 115.590 159.090 ;
        RECT 119.315 158.375 119.645 159.525 ;
        RECT 120.155 158.725 120.485 159.525 ;
        RECT 121.005 158.725 121.245 159.525 ;
        RECT 122.845 158.435 126.355 159.525 ;
        RECT 126.525 158.435 127.735 159.525 ;
        RECT 122.845 157.915 124.535 158.435 ;
        RECT 126.525 157.895 127.045 158.435 ;
        RECT 15.435 155.345 15.955 155.885 ;
        RECT 14.745 154.255 15.955 155.345 ;
        RECT 28.545 155.345 30.235 155.865 ;
        RECT 35.905 155.345 36.425 155.885 ;
        RECT 17.395 154.255 17.680 155.055 ;
        RECT 18.800 154.255 19.130 154.945 ;
        RECT 19.800 154.255 20.220 154.635 ;
        RECT 21.500 154.255 21.830 154.635 ;
        RECT 22.350 154.255 22.730 154.635 ;
        RECT 24.375 154.255 24.705 154.755 ;
        RECT 25.315 154.255 25.645 154.755 ;
        RECT 26.685 154.255 27.015 155.015 ;
        RECT 28.545 154.255 32.055 155.345 ;
        RECT 32.795 154.255 33.065 154.715 ;
        RECT 34.855 154.255 35.180 154.715 ;
        RECT 35.905 154.255 37.115 155.345 ;
        RECT 37.285 154.255 37.575 155.420 ;
        RECT 38.205 155.345 38.955 155.865 ;
        RECT 38.205 154.255 39.875 155.345 ;
        RECT 40.555 154.255 40.725 155.395 ;
        RECT 40.995 154.255 41.245 155.055 ;
        RECT 42.520 154.255 42.850 155.055 ;
        RECT 44.235 154.255 44.405 155.395 ;
        RECT 44.675 154.255 44.925 155.055 ;
        RECT 46.200 154.255 46.530 155.055 ;
        RECT 48.110 154.255 48.440 155.055 ;
        RECT 49.715 154.255 49.965 155.055 ;
        RECT 50.235 154.255 50.405 155.395 ;
        RECT 51.545 155.345 52.295 155.865 ;
        RECT 51.545 154.255 53.215 155.345 ;
        RECT 54.195 154.255 54.480 155.055 ;
        RECT 55.600 154.255 55.930 154.945 ;
        RECT 56.600 154.255 57.020 154.635 ;
        RECT 58.300 154.255 58.630 154.635 ;
        RECT 59.150 154.255 59.530 154.635 ;
        RECT 61.175 154.255 61.505 154.755 ;
        RECT 62.115 154.255 62.445 154.755 ;
        RECT 63.045 154.255 63.335 155.420 ;
        RECT 63.545 154.255 63.775 155.395 ;
        RECT 64.445 154.255 64.655 155.395 ;
        RECT 64.885 155.345 65.635 155.865 ;
        RECT 64.885 154.255 66.555 155.345 ;
        RECT 66.815 154.255 67.085 155.000 ;
        RECT 67.715 154.260 67.970 154.985 ;
        RECT 68.585 154.260 68.830 154.985 ;
        RECT 69.445 154.260 69.690 154.985 ;
        RECT 70.305 154.260 70.550 154.985 ;
        RECT 71.150 154.260 71.410 154.985 ;
        RECT 72.010 154.260 72.270 154.985 ;
        RECT 72.870 154.260 73.130 154.985 ;
        RECT 73.730 154.260 73.990 155.055 ;
        RECT 67.715 154.255 73.990 154.260 ;
        RECT 74.590 154.255 74.850 155.065 ;
        RECT 75.450 154.255 75.745 155.065 ;
        RECT 76.630 154.255 76.960 155.055 ;
        RECT 78.235 154.255 78.485 155.055 ;
        RECT 78.755 154.255 78.925 155.395 ;
        RECT 81.035 154.255 81.205 155.395 ;
        RECT 85.125 155.345 86.815 155.865 ;
        RECT 81.475 154.255 81.725 155.055 ;
        RECT 83.000 154.255 83.330 155.055 ;
        RECT 85.125 154.255 88.635 155.345 ;
        RECT 88.805 154.255 89.095 155.420 ;
        RECT 89.265 155.345 90.475 155.865 ;
        RECT 89.265 154.255 91.855 155.345 ;
        RECT 93.620 154.690 93.970 155.940 ;
        RECT 92.030 154.255 97.375 154.690 ;
        RECT 98.055 154.255 98.225 155.395 ;
        RECT 101.685 155.345 102.435 155.865 ;
        RECT 98.495 154.255 98.745 155.055 ;
        RECT 100.020 154.255 100.350 155.055 ;
        RECT 101.685 154.255 103.355 155.345 ;
        RECT 104.230 154.255 104.560 155.055 ;
        RECT 105.835 154.255 106.085 155.055 ;
        RECT 106.355 154.255 106.525 155.395 ;
        RECT 107.910 154.255 108.240 155.055 ;
        RECT 109.515 154.255 109.765 155.055 ;
        RECT 110.035 154.255 110.205 155.395 ;
        RECT 111.395 154.255 111.565 155.395 ;
        RECT 111.835 154.255 112.085 155.055 ;
        RECT 113.360 154.255 113.690 155.055 ;
        RECT 114.565 154.255 114.855 155.420 ;
        RECT 115.025 155.345 115.545 155.885 ;
        RECT 115.025 154.255 116.235 155.345 ;
        RECT 116.915 154.255 117.155 155.055 ;
        RECT 117.675 154.255 118.005 155.055 ;
        RECT 118.515 154.255 118.845 155.405 ;
        RECT 119.165 155.345 119.915 155.865 ;
        RECT 119.165 154.255 120.835 155.345 ;
        RECT 122.600 154.690 122.950 155.940 ;
        RECT 126.525 155.345 127.045 155.885 ;
        RECT 121.010 154.255 126.355 154.690 ;
        RECT 126.525 154.255 127.735 155.345 ;
        RECT 14.660 154.085 127.820 154.255 ;
        RECT 14.745 152.995 15.955 154.085 ;
        RECT 15.435 152.455 15.955 152.995 ;
        RECT 16.585 152.995 20.095 154.085 ;
        RECT 21.015 153.325 21.185 154.085 ;
        RECT 16.585 152.475 18.275 152.995 ;
        RECT 23.555 152.945 23.725 154.085 ;
        RECT 24.405 152.920 24.695 154.085 ;
        RECT 25.330 153.650 30.675 154.085 ;
        RECT 26.920 152.400 27.270 153.650 ;
        RECT 30.885 152.945 31.115 154.085 ;
        RECT 31.785 152.945 31.995 154.085 ;
        RECT 32.665 153.325 32.995 154.085 ;
        RECT 34.115 152.945 34.285 154.085 ;
        RECT 36.655 153.325 36.825 154.085 ;
        RECT 38.255 152.945 38.425 154.085 ;
        RECT 38.695 153.285 38.945 154.085 ;
        RECT 40.220 153.285 40.550 154.085 ;
        RECT 41.885 152.995 44.475 154.085 ;
        RECT 44.650 153.650 49.995 154.085 ;
        RECT 41.885 152.475 43.095 152.995 ;
        RECT 46.240 152.400 46.590 153.650 ;
        RECT 50.165 152.920 50.455 154.085 ;
        RECT 51.550 153.650 56.895 154.085 ;
        RECT 53.140 152.400 53.490 153.650 ;
        RECT 57.105 152.945 57.335 154.085 ;
        RECT 58.005 152.945 58.215 154.085 ;
        RECT 59.255 153.285 59.540 154.085 ;
        RECT 60.660 153.395 60.990 154.085 ;
        RECT 61.660 153.705 62.080 154.085 ;
        RECT 63.360 153.705 63.690 154.085 ;
        RECT 64.210 153.705 64.590 154.085 ;
        RECT 66.235 153.585 66.565 154.085 ;
        RECT 67.175 153.585 67.505 154.085 ;
        RECT 68.565 152.995 71.155 154.085 ;
        RECT 71.800 153.325 72.130 154.085 ;
        RECT 68.565 152.475 69.775 152.995 ;
        RECT 72.730 152.935 72.990 154.085 ;
        RECT 73.175 153.025 73.505 154.085 ;
        RECT 74.525 153.725 74.855 154.085 ;
        RECT 75.925 152.920 76.215 154.085 ;
        RECT 76.845 152.995 79.435 154.085 ;
        RECT 79.610 153.650 84.955 154.085 ;
        RECT 85.130 153.650 90.475 154.085 ;
        RECT 76.845 152.475 78.055 152.995 ;
        RECT 81.200 152.400 81.550 153.650 ;
        RECT 86.720 152.400 87.070 153.650 ;
        RECT 90.685 152.945 90.915 154.085 ;
        RECT 91.585 152.945 91.795 154.085 ;
        RECT 92.485 152.995 95.995 154.085 ;
        RECT 96.170 153.650 101.515 154.085 ;
        RECT 92.485 152.475 94.175 152.995 ;
        RECT 97.760 152.400 98.110 153.650 ;
        RECT 101.685 152.920 101.975 154.085 ;
        RECT 102.605 152.995 105.195 154.085 ;
        RECT 102.605 152.475 103.815 152.995 ;
        RECT 105.875 152.945 106.045 154.085 ;
        RECT 106.315 153.285 106.565 154.085 ;
        RECT 107.840 153.285 108.170 154.085 ;
        RECT 109.555 152.945 109.725 154.085 ;
        RECT 109.995 153.285 110.245 154.085 ;
        RECT 111.520 153.285 111.850 154.085 ;
        RECT 113.190 153.650 118.535 154.085 ;
        RECT 114.780 152.400 115.130 153.650 ;
        RECT 118.765 152.945 118.975 154.085 ;
        RECT 119.645 152.945 119.875 154.085 ;
        RECT 120.985 153.325 121.315 154.085 ;
        RECT 122.845 152.995 126.355 154.085 ;
        RECT 126.525 152.995 127.735 154.085 ;
        RECT 122.845 152.475 124.535 152.995 ;
        RECT 126.525 152.455 127.045 152.995 ;
        RECT 15.435 149.905 15.955 150.445 ;
        RECT 14.745 148.815 15.955 149.905 ;
        RECT 25.785 149.905 26.535 150.425 ;
        RECT 16.935 148.815 17.220 149.615 ;
        RECT 18.340 148.815 18.670 149.505 ;
        RECT 19.340 148.815 19.760 149.195 ;
        RECT 21.040 148.815 21.370 149.195 ;
        RECT 21.890 148.815 22.270 149.195 ;
        RECT 23.915 148.815 24.245 149.315 ;
        RECT 24.855 148.815 25.185 149.315 ;
        RECT 25.785 148.815 27.455 149.905 ;
        RECT 28.435 148.815 28.720 149.615 ;
        RECT 29.840 148.815 30.170 149.505 ;
        RECT 30.840 148.815 31.260 149.195 ;
        RECT 32.540 148.815 32.870 149.195 ;
        RECT 33.390 148.815 33.770 149.195 ;
        RECT 35.415 148.815 35.745 149.315 ;
        RECT 36.355 148.815 36.685 149.315 ;
        RECT 37.285 148.815 37.575 149.980 ;
        RECT 38.205 149.905 39.415 150.425 ;
        RECT 38.205 148.815 40.795 149.905 ;
        RECT 41.670 148.815 42.000 149.615 ;
        RECT 43.275 148.815 43.525 149.615 ;
        RECT 43.795 148.815 43.965 149.955 ;
        RECT 44.645 149.905 45.165 150.445 ;
        RECT 44.645 148.815 45.855 149.905 ;
        RECT 47.855 148.815 48.135 149.615 ;
        RECT 50.615 148.815 50.895 149.615 ;
        RECT 52.055 148.815 52.225 149.955 ;
        RECT 55.685 149.905 56.435 150.425 ;
        RECT 52.495 148.815 52.745 149.615 ;
        RECT 54.020 148.815 54.350 149.615 ;
        RECT 55.685 148.815 57.355 149.905 ;
        RECT 58.275 148.815 58.445 149.575 ;
        RECT 60.815 148.815 60.985 149.955 ;
        RECT 62.105 148.815 62.435 149.575 ;
        RECT 63.045 148.815 63.335 149.980 ;
        RECT 65.805 149.905 66.555 150.425 ;
        RECT 64.405 148.815 64.735 149.575 ;
        RECT 65.805 148.815 67.475 149.905 ;
        RECT 68.120 148.815 68.450 149.575 ;
        RECT 69.050 148.815 69.310 149.965 ;
        RECT 69.490 148.815 69.750 149.965 ;
        RECT 80.985 149.905 82.675 150.425 ;
        RECT 70.350 148.815 70.680 149.575 ;
        RECT 71.380 148.815 71.665 149.685 ;
        RECT 72.270 148.815 72.525 149.275 ;
        RECT 73.125 148.815 73.435 149.615 ;
        RECT 75.485 148.815 75.795 149.615 ;
        RECT 76.395 148.815 76.650 149.275 ;
        RECT 77.255 148.815 77.540 149.685 ;
        RECT 79.595 148.815 79.875 149.615 ;
        RECT 80.985 148.815 84.495 149.905 ;
        RECT 85.415 148.815 85.585 149.575 ;
        RECT 87.955 148.815 88.125 149.955 ;
        RECT 88.805 148.815 89.095 149.980 ;
        RECT 89.695 148.815 90.025 149.315 ;
        RECT 90.635 148.815 90.965 149.315 ;
        RECT 92.610 148.815 92.990 149.195 ;
        RECT 93.510 148.815 93.840 149.195 ;
        RECT 95.120 148.815 95.540 149.195 ;
        RECT 96.210 148.815 96.540 149.505 ;
        RECT 97.660 148.815 97.945 149.615 ;
        RECT 100.520 149.250 100.870 150.500 ;
        RECT 98.930 148.815 104.275 149.250 ;
        RECT 104.925 148.815 105.205 149.615 ;
        RECT 107.715 148.815 107.885 149.955 ;
        RECT 108.155 148.815 108.405 149.615 ;
        RECT 109.680 148.815 110.010 149.615 ;
        RECT 111.455 148.815 111.725 149.275 ;
        RECT 113.515 148.815 113.840 149.275 ;
        RECT 114.565 148.815 114.855 149.980 ;
        RECT 116.375 148.815 116.680 149.955 ;
        RECT 125.145 149.905 125.665 150.445 ;
        RECT 126.525 149.905 127.045 150.445 ;
        RECT 117.020 148.815 117.350 149.195 ;
        RECT 117.870 148.815 118.120 149.275 ;
        RECT 119.735 148.815 120.105 149.275 ;
        RECT 120.740 148.815 121.070 149.245 ;
        RECT 122.960 148.815 123.210 149.275 ;
        RECT 124.215 148.815 124.545 149.315 ;
        RECT 125.145 148.815 126.355 149.905 ;
        RECT 126.525 148.815 127.735 149.905 ;
        RECT 14.660 148.645 127.820 148.815 ;
        RECT 14.745 147.555 15.955 148.645 ;
        RECT 15.435 147.015 15.955 147.555 ;
        RECT 16.585 147.555 20.095 148.645 ;
        RECT 21.015 147.885 21.185 148.645 ;
        RECT 16.585 147.035 18.275 147.555 ;
        RECT 23.555 147.505 23.725 148.645 ;
        RECT 24.405 147.480 24.695 148.645 ;
        RECT 25.365 147.505 25.595 148.645 ;
        RECT 26.265 147.505 26.475 148.645 ;
        RECT 27.145 147.885 27.475 148.645 ;
        RECT 28.525 147.885 28.855 148.645 ;
        RECT 29.975 147.505 30.145 148.645 ;
        RECT 32.515 147.885 32.685 148.645 ;
        RECT 34.065 147.555 35.735 148.645 ;
        RECT 36.610 147.845 36.940 148.645 ;
        RECT 38.215 147.845 38.465 148.645 ;
        RECT 34.065 147.035 34.815 147.555 ;
        RECT 38.735 147.505 38.905 148.645 ;
        RECT 40.095 147.505 40.265 148.645 ;
        RECT 40.535 147.845 40.785 148.645 ;
        RECT 42.060 147.845 42.390 148.645 ;
        RECT 43.265 147.555 44.475 148.645 ;
        RECT 44.650 148.210 49.995 148.645 ;
        RECT 43.265 147.015 43.785 147.555 ;
        RECT 46.240 146.960 46.590 148.210 ;
        RECT 50.165 147.480 50.455 148.645 ;
        RECT 52.055 147.505 52.225 148.645 ;
        RECT 54.595 147.885 54.765 148.645 ;
        RECT 56.195 147.505 56.365 148.645 ;
        RECT 56.635 147.845 56.885 148.645 ;
        RECT 58.160 147.845 58.490 148.645 ;
        RECT 60.575 147.885 60.745 148.645 ;
        RECT 63.115 147.505 63.285 148.645 ;
        RECT 63.965 147.555 65.175 148.645 ;
        RECT 65.350 148.210 70.695 148.645 ;
        RECT 63.965 147.015 64.485 147.555 ;
        RECT 66.940 146.960 67.290 148.210 ;
        RECT 70.870 147.495 71.130 148.645 ;
        RECT 71.730 147.885 72.060 148.645 ;
        RECT 73.180 147.885 73.510 148.645 ;
        RECT 74.110 147.495 74.370 148.645 ;
        RECT 74.545 147.555 75.755 148.645 ;
        RECT 74.545 147.015 75.065 147.555 ;
        RECT 75.925 147.480 76.215 148.645 ;
        RECT 77.090 147.845 77.420 148.645 ;
        RECT 78.695 147.845 78.945 148.645 ;
        RECT 79.215 147.505 79.385 148.645 ;
        RECT 80.575 147.505 80.745 148.645 ;
        RECT 81.015 147.845 81.265 148.645 ;
        RECT 82.540 147.845 82.870 148.645 ;
        RECT 83.805 147.505 84.015 148.645 ;
        RECT 84.685 147.505 84.915 148.645 ;
        RECT 85.935 147.845 86.220 148.645 ;
        RECT 87.340 147.955 87.670 148.645 ;
        RECT 88.340 148.265 88.760 148.645 ;
        RECT 90.040 148.265 90.370 148.645 ;
        RECT 90.890 148.265 91.270 148.645 ;
        RECT 92.915 148.145 93.245 148.645 ;
        RECT 93.855 148.145 94.185 148.645 ;
        RECT 95.745 147.505 95.975 148.645 ;
        RECT 96.645 147.505 96.855 148.645 ;
        RECT 97.835 147.885 98.005 148.645 ;
        RECT 100.375 147.505 100.545 148.645 ;
        RECT 101.685 147.480 101.975 148.645 ;
        RECT 102.585 147.885 102.915 148.645 ;
        RECT 104.465 147.845 104.745 148.645 ;
        RECT 107.255 147.505 107.425 148.645 ;
        RECT 107.695 147.845 107.945 148.645 ;
        RECT 109.220 147.845 109.550 148.645 ;
        RECT 110.425 147.555 112.095 148.645 ;
        RECT 113.015 147.885 113.185 148.645 ;
        RECT 110.425 147.035 111.175 147.555 ;
        RECT 115.555 147.505 115.725 148.645 ;
        RECT 117.215 147.845 117.500 148.645 ;
        RECT 118.620 147.955 118.950 148.645 ;
        RECT 119.620 148.265 120.040 148.645 ;
        RECT 121.320 148.265 121.650 148.645 ;
        RECT 122.170 148.265 122.550 148.645 ;
        RECT 124.195 148.145 124.525 148.645 ;
        RECT 125.135 148.145 125.465 148.645 ;
        RECT 126.525 147.555 127.735 148.645 ;
        RECT 126.525 147.015 127.045 147.555 ;
        RECT 15.435 144.465 15.955 145.005 ;
        RECT 14.745 143.375 15.955 144.465 ;
        RECT 16.585 144.465 18.275 144.985 ;
        RECT 16.585 143.375 20.095 144.465 ;
        RECT 20.325 143.375 20.535 144.515 ;
        RECT 21.205 143.375 21.435 144.515 ;
        RECT 22.915 143.375 23.200 144.175 ;
        RECT 24.320 143.375 24.650 144.065 ;
        RECT 25.320 143.375 25.740 143.755 ;
        RECT 27.020 143.375 27.350 143.755 ;
        RECT 27.870 143.375 28.250 143.755 ;
        RECT 29.895 143.375 30.225 143.875 ;
        RECT 30.835 143.375 31.165 143.875 ;
        RECT 33.360 143.810 33.710 145.060 ;
        RECT 31.770 143.375 37.115 143.810 ;
        RECT 37.285 143.375 37.575 144.540 ;
        RECT 38.205 144.465 39.415 144.985 ;
        RECT 38.205 143.375 40.795 144.465 ;
        RECT 41.005 143.375 41.235 144.515 ;
        RECT 41.905 143.375 42.115 144.515 ;
        RECT 53.385 144.465 53.905 145.005 ;
        RECT 54.765 144.465 56.455 144.985 ;
        RECT 42.775 143.375 43.105 143.875 ;
        RECT 43.715 143.375 44.045 143.875 ;
        RECT 45.690 143.375 46.070 143.755 ;
        RECT 46.590 143.375 46.920 143.755 ;
        RECT 48.200 143.375 48.620 143.755 ;
        RECT 49.290 143.375 49.620 144.065 ;
        RECT 50.740 143.375 51.025 144.175 ;
        RECT 52.445 143.375 52.775 144.135 ;
        RECT 53.385 143.375 54.595 144.465 ;
        RECT 54.765 143.375 58.275 144.465 ;
        RECT 58.485 143.375 58.715 144.515 ;
        RECT 59.385 143.375 59.595 144.515 ;
        RECT 60.285 144.465 61.495 144.985 ;
        RECT 60.285 143.375 62.875 144.465 ;
        RECT 63.045 143.375 63.335 144.540 ;
        RECT 64.715 143.375 64.885 144.135 ;
        RECT 67.255 143.375 67.425 144.515 ;
        RECT 70.160 143.810 70.510 145.060 ;
        RECT 75.680 143.810 76.030 145.060 ;
        RECT 82.825 144.465 83.575 144.985 ;
        RECT 68.570 143.375 73.915 143.810 ;
        RECT 74.090 143.375 79.435 143.810 ;
        RECT 81.435 143.375 81.715 144.175 ;
        RECT 82.825 143.375 84.495 144.465 ;
        RECT 85.415 143.375 85.585 144.135 ;
        RECT 87.955 143.375 88.125 144.515 ;
        RECT 88.805 143.375 89.095 144.540 ;
        RECT 90.625 143.375 90.955 144.135 ;
        RECT 92.005 143.375 92.335 144.135 ;
        RECT 93.515 143.375 93.785 143.835 ;
        RECT 95.575 143.375 95.900 143.835 ;
        RECT 97.055 143.375 97.360 144.515 ;
        RECT 106.285 144.465 107.975 144.985 ;
        RECT 97.700 143.375 98.030 143.755 ;
        RECT 98.550 143.375 98.800 143.835 ;
        RECT 100.415 143.375 100.785 143.835 ;
        RECT 101.420 143.375 101.750 143.805 ;
        RECT 103.640 143.375 103.890 143.835 ;
        RECT 104.895 143.375 105.225 143.875 ;
        RECT 106.285 143.375 109.795 144.465 ;
        RECT 110.670 143.375 111.000 144.175 ;
        RECT 112.275 143.375 112.525 144.175 ;
        RECT 112.795 143.375 112.965 144.515 ;
        RECT 114.565 143.375 114.855 144.540 ;
        RECT 116.235 143.375 116.405 144.135 ;
        RECT 118.775 143.375 118.945 144.515 ;
        RECT 119.665 143.375 119.895 144.515 ;
        RECT 120.565 143.375 120.775 144.515 ;
        RECT 122.845 144.465 124.535 144.985 ;
        RECT 126.525 144.465 127.045 145.005 ;
        RECT 121.905 143.375 122.235 144.135 ;
        RECT 122.845 143.375 126.355 144.465 ;
        RECT 126.525 143.375 127.735 144.465 ;
        RECT 14.660 143.205 127.820 143.375 ;
        RECT 14.745 142.115 15.955 143.205 ;
        RECT 15.435 141.575 15.955 142.115 ;
        RECT 16.125 142.115 18.715 143.205 ;
        RECT 18.890 142.770 24.235 143.205 ;
        RECT 16.125 141.595 17.335 142.115 ;
        RECT 20.480 141.520 20.830 142.770 ;
        RECT 24.405 142.040 24.695 143.205 ;
        RECT 25.325 142.115 28.835 143.205 ;
        RECT 29.010 142.770 34.355 143.205 ;
        RECT 25.325 141.595 27.015 142.115 ;
        RECT 30.600 141.520 30.950 142.770 ;
        RECT 35.005 142.405 35.285 143.205 ;
        RECT 38.205 142.115 41.715 143.205 ;
        RECT 41.890 142.770 47.235 143.205 ;
        RECT 38.205 141.595 39.895 142.115 ;
        RECT 43.480 141.520 43.830 142.770 ;
        RECT 49.235 142.405 49.515 143.205 ;
        RECT 50.165 142.040 50.455 143.205 ;
        RECT 50.625 142.115 52.295 143.205 ;
        RECT 50.625 141.595 51.375 142.115 ;
        RECT 52.975 142.065 53.145 143.205 ;
        RECT 53.415 142.405 53.665 143.205 ;
        RECT 54.940 142.405 55.270 143.205 ;
        RECT 56.715 142.745 56.985 143.205 ;
        RECT 58.775 142.745 59.100 143.205 ;
        RECT 60.255 142.065 60.560 143.205 ;
        RECT 60.900 142.825 61.230 143.205 ;
        RECT 61.750 142.745 62.000 143.205 ;
        RECT 63.615 142.745 63.985 143.205 ;
        RECT 64.620 142.775 64.950 143.205 ;
        RECT 66.840 142.745 67.090 143.205 ;
        RECT 68.095 142.705 68.425 143.205 ;
        RECT 69.465 142.445 69.795 143.205 ;
        RECT 70.405 142.115 71.615 143.205 ;
        RECT 70.405 141.575 70.925 142.115 ;
        RECT 71.825 142.065 72.055 143.205 ;
        RECT 72.725 142.065 72.935 143.205 ;
        RECT 73.165 142.115 75.755 143.205 ;
        RECT 73.165 141.595 74.375 142.115 ;
        RECT 75.925 142.040 76.215 143.205 ;
        RECT 76.845 142.115 79.435 143.205 ;
        RECT 79.610 142.770 84.955 143.205 ;
        RECT 85.130 142.770 90.475 143.205 ;
        RECT 90.650 142.770 95.995 143.205 ;
        RECT 96.170 142.770 101.515 143.205 ;
        RECT 76.845 141.595 78.055 142.115 ;
        RECT 81.200 141.520 81.550 142.770 ;
        RECT 86.720 141.520 87.070 142.770 ;
        RECT 92.240 141.520 92.590 142.770 ;
        RECT 97.760 141.520 98.110 142.770 ;
        RECT 101.685 142.040 101.975 143.205 ;
        RECT 103.070 142.770 108.415 143.205 ;
        RECT 104.660 141.520 105.010 142.770 ;
        RECT 110.415 142.405 110.695 143.205 ;
        RECT 112.265 142.115 115.775 143.205 ;
        RECT 116.695 142.445 116.865 143.205 ;
        RECT 112.265 141.595 113.955 142.115 ;
        RECT 119.235 142.065 119.405 143.205 ;
        RECT 120.125 142.065 120.355 143.205 ;
        RECT 121.025 142.065 121.235 143.205 ;
        RECT 121.465 142.115 122.675 143.205 ;
        RECT 122.845 142.115 126.355 143.205 ;
        RECT 126.525 142.115 127.735 143.205 ;
        RECT 121.465 141.575 121.985 142.115 ;
        RECT 122.845 141.595 124.535 142.115 ;
        RECT 126.525 141.575 127.045 142.115 ;
        RECT 15.435 139.025 15.955 139.565 ;
        RECT 14.745 137.935 15.955 139.025 ;
        RECT 25.785 139.025 26.995 139.545 ;
        RECT 16.935 137.935 17.220 138.735 ;
        RECT 18.340 137.935 18.670 138.625 ;
        RECT 19.340 137.935 19.760 138.315 ;
        RECT 21.040 137.935 21.370 138.315 ;
        RECT 21.890 137.935 22.270 138.315 ;
        RECT 23.915 137.935 24.245 138.435 ;
        RECT 24.855 137.935 25.185 138.435 ;
        RECT 25.785 137.935 28.375 139.025 ;
        RECT 30.140 138.370 30.490 139.620 ;
        RECT 28.550 137.935 33.895 138.370 ;
        RECT 34.265 137.935 34.545 138.605 ;
        RECT 35.215 137.935 35.545 138.655 ;
        RECT 37.285 137.935 37.575 139.100 ;
        RECT 39.145 137.935 39.425 138.735 ;
        RECT 43.020 138.370 43.370 139.620 ;
        RECT 41.430 137.935 46.775 138.370 ;
        RECT 48.775 137.935 49.055 138.735 ;
        RECT 50.215 137.935 50.385 139.075 ;
        RECT 53.385 139.025 54.135 139.545 ;
        RECT 50.655 137.935 50.905 138.735 ;
        RECT 52.180 137.935 52.510 138.735 ;
        RECT 53.385 137.935 55.055 139.025 ;
        RECT 55.265 137.935 55.495 139.075 ;
        RECT 56.165 137.935 56.375 139.075 ;
        RECT 56.605 139.025 57.815 139.545 ;
        RECT 56.605 137.935 59.195 139.025 ;
        RECT 59.875 137.935 60.045 139.075 ;
        RECT 60.315 137.935 60.565 138.735 ;
        RECT 61.840 137.935 62.170 138.735 ;
        RECT 63.045 137.935 63.335 139.100 ;
        RECT 64.475 137.935 64.645 139.075 ;
        RECT 77.305 139.025 78.515 139.545 ;
        RECT 64.915 137.935 65.165 138.735 ;
        RECT 66.440 137.935 66.770 138.735 ;
        RECT 68.075 137.935 68.405 138.435 ;
        RECT 69.015 137.935 69.345 138.435 ;
        RECT 70.990 137.935 71.370 138.315 ;
        RECT 71.890 137.935 72.220 138.315 ;
        RECT 73.500 137.935 73.920 138.315 ;
        RECT 74.590 137.935 74.920 138.625 ;
        RECT 76.040 137.935 76.325 138.735 ;
        RECT 77.305 137.935 79.895 139.025 ;
        RECT 80.575 137.935 80.745 139.075 ;
        RECT 81.015 137.935 81.265 138.735 ;
        RECT 82.540 137.935 82.870 138.735 ;
        RECT 85.415 137.935 85.585 138.695 ;
        RECT 87.955 137.935 88.125 139.075 ;
        RECT 88.805 137.935 89.095 139.100 ;
        RECT 92.025 139.025 93.715 139.545 ;
        RECT 90.165 137.935 90.495 138.695 ;
        RECT 92.025 137.935 95.535 139.025 ;
        RECT 97.300 138.370 97.650 139.620 ;
        RECT 95.710 137.935 101.055 138.370 ;
        RECT 101.265 137.935 101.495 139.075 ;
        RECT 102.165 137.935 102.375 139.075 ;
        RECT 102.605 139.025 104.295 139.545 ;
        RECT 102.605 137.935 106.115 139.025 ;
        RECT 106.795 137.935 106.965 139.075 ;
        RECT 107.235 137.935 107.485 138.735 ;
        RECT 108.760 137.935 109.090 138.735 ;
        RECT 110.670 137.935 111.000 138.735 ;
        RECT 112.275 137.935 112.525 138.735 ;
        RECT 112.795 137.935 112.965 139.075 ;
        RECT 114.565 137.935 114.855 139.100 ;
        RECT 115.525 137.935 115.755 139.075 ;
        RECT 116.425 137.935 116.635 139.075 ;
        RECT 126.525 139.025 127.045 139.565 ;
        RECT 117.675 137.935 117.960 138.735 ;
        RECT 119.080 137.935 119.410 138.625 ;
        RECT 120.080 137.935 120.500 138.315 ;
        RECT 121.780 137.935 122.110 138.315 ;
        RECT 122.630 137.935 123.010 138.315 ;
        RECT 124.655 137.935 124.985 138.435 ;
        RECT 125.595 137.935 125.925 138.435 ;
        RECT 126.525 137.935 127.735 139.025 ;
        RECT 14.660 137.765 127.820 137.935 ;
        RECT 14.745 136.675 15.955 137.765 ;
        RECT 16.130 137.330 21.475 137.765 ;
        RECT 15.435 136.135 15.955 136.675 ;
        RECT 17.720 136.080 18.070 137.330 ;
        RECT 22.085 137.005 22.415 137.765 ;
        RECT 23.065 136.625 23.295 137.765 ;
        RECT 23.965 136.625 24.175 137.765 ;
        RECT 24.405 136.600 24.695 137.765 ;
        RECT 25.325 136.675 28.835 137.765 ;
        RECT 29.755 137.005 29.925 137.765 ;
        RECT 25.325 136.155 27.015 136.675 ;
        RECT 32.295 136.625 32.465 137.765 ;
        RECT 33.145 136.675 34.815 137.765 ;
        RECT 35.465 136.965 35.745 137.765 ;
        RECT 37.945 137.095 38.225 137.765 ;
        RECT 38.895 137.045 39.225 137.765 ;
        RECT 40.045 136.675 43.555 137.765 ;
        RECT 44.205 136.965 44.485 137.765 ;
        RECT 46.485 136.675 49.995 137.765 ;
        RECT 33.145 136.155 33.895 136.675 ;
        RECT 40.045 136.155 41.735 136.675 ;
        RECT 46.485 136.155 48.175 136.675 ;
        RECT 50.165 136.600 50.455 137.765 ;
        RECT 51.085 136.675 52.755 137.765 ;
        RECT 53.675 137.005 53.845 137.765 ;
        RECT 51.085 136.155 51.835 136.675 ;
        RECT 56.215 136.625 56.385 137.765 ;
        RECT 57.965 137.005 58.295 137.765 ;
        RECT 59.365 136.675 61.035 137.765 ;
        RECT 59.365 136.155 60.115 136.675 ;
        RECT 61.715 136.625 61.885 137.765 ;
        RECT 62.155 136.965 62.405 137.765 ;
        RECT 63.680 136.965 64.010 137.765 ;
        RECT 65.345 136.675 67.015 137.765 ;
        RECT 67.615 136.985 67.865 137.765 ;
        RECT 68.535 137.385 68.890 137.765 ;
        RECT 70.960 137.305 71.285 137.765 ;
        RECT 73.075 137.305 73.345 137.765 ;
        RECT 74.085 136.675 75.755 137.765 ;
        RECT 65.345 136.155 66.095 136.675 ;
        RECT 74.085 136.155 74.835 136.675 ;
        RECT 75.925 136.600 76.215 137.765 ;
        RECT 77.785 136.965 78.065 137.765 ;
        RECT 80.575 136.625 80.745 137.765 ;
        RECT 81.015 136.965 81.265 137.765 ;
        RECT 82.540 136.965 82.870 137.765 ;
        RECT 84.555 136.965 84.840 137.765 ;
        RECT 85.960 137.075 86.290 137.765 ;
        RECT 86.960 137.385 87.380 137.765 ;
        RECT 88.660 137.385 88.990 137.765 ;
        RECT 89.510 137.385 89.890 137.765 ;
        RECT 91.535 137.265 91.865 137.765 ;
        RECT 92.475 137.265 92.805 137.765 ;
        RECT 94.155 137.005 94.325 137.765 ;
        RECT 96.695 136.625 96.865 137.765 ;
        RECT 98.710 136.965 99.040 137.765 ;
        RECT 100.315 136.965 100.565 137.765 ;
        RECT 100.835 136.625 101.005 137.765 ;
        RECT 101.685 136.600 101.975 137.765 ;
        RECT 103.815 137.005 103.985 137.765 ;
        RECT 106.355 136.625 106.525 137.765 ;
        RECT 107.645 137.005 107.975 137.765 ;
        RECT 110.255 137.005 110.425 137.765 ;
        RECT 112.795 136.625 112.965 137.765 ;
        RECT 114.455 136.965 114.740 137.765 ;
        RECT 115.860 137.075 116.190 137.765 ;
        RECT 116.860 137.385 117.280 137.765 ;
        RECT 118.560 137.385 118.890 137.765 ;
        RECT 119.410 137.385 119.790 137.765 ;
        RECT 121.435 137.265 121.765 137.765 ;
        RECT 122.375 137.265 122.705 137.765 ;
        RECT 123.745 137.005 124.075 137.765 ;
        RECT 124.685 136.675 126.355 137.765 ;
        RECT 126.525 136.675 127.735 137.765 ;
        RECT 124.685 136.155 125.435 136.675 ;
        RECT 126.525 136.135 127.045 136.675 ;
        RECT 15.435 133.585 15.955 134.125 ;
        RECT 14.745 132.495 15.955 133.585 ;
        RECT 16.185 132.495 16.395 133.635 ;
        RECT 17.065 132.495 17.295 133.635 ;
        RECT 18.255 132.495 18.425 133.255 ;
        RECT 20.795 132.495 20.965 133.635 ;
        RECT 22.455 132.495 22.740 133.295 ;
        RECT 23.860 132.495 24.190 133.185 ;
        RECT 24.860 132.495 25.280 132.875 ;
        RECT 26.560 132.495 26.890 132.875 ;
        RECT 27.410 132.495 27.790 132.875 ;
        RECT 29.435 132.495 29.765 132.995 ;
        RECT 30.375 132.495 30.705 132.995 ;
        RECT 31.745 132.495 32.075 133.255 ;
        RECT 33.895 132.495 34.065 133.255 ;
        RECT 36.435 132.495 36.605 133.635 ;
        RECT 37.285 132.495 37.575 133.660 ;
        RECT 40.505 133.585 41.025 134.125 ;
        RECT 38.225 132.495 38.505 133.295 ;
        RECT 40.505 132.495 41.715 133.585 ;
        RECT 43.715 132.495 43.995 133.295 ;
        RECT 45.155 132.495 45.325 133.635 ;
        RECT 45.595 132.495 45.845 133.295 ;
        RECT 47.120 132.495 47.450 133.295 ;
        RECT 48.835 132.495 49.005 133.635 ;
        RECT 61.665 133.585 62.185 134.125 ;
        RECT 49.275 132.495 49.525 133.295 ;
        RECT 50.800 132.495 51.130 133.295 ;
        RECT 52.815 132.495 53.100 133.295 ;
        RECT 54.220 132.495 54.550 133.185 ;
        RECT 55.220 132.495 55.640 132.875 ;
        RECT 56.920 132.495 57.250 132.875 ;
        RECT 57.770 132.495 58.150 132.875 ;
        RECT 59.795 132.495 60.125 132.995 ;
        RECT 60.735 132.495 61.065 132.995 ;
        RECT 61.665 132.495 62.875 133.585 ;
        RECT 63.045 132.495 63.335 133.660 ;
        RECT 64.015 132.495 64.185 133.635 ;
        RECT 64.455 132.495 64.705 133.295 ;
        RECT 65.980 132.495 66.310 133.295 ;
        RECT 69.700 132.930 70.050 134.180 ;
        RECT 75.220 132.930 75.570 134.180 ;
        RECT 68.110 132.495 73.455 132.930 ;
        RECT 73.630 132.495 78.975 132.930 ;
        RECT 80.975 132.495 81.255 133.295 ;
        RECT 83.500 132.930 83.850 134.180 ;
        RECT 81.910 132.495 87.255 132.930 ;
        RECT 87.485 132.495 87.695 133.635 ;
        RECT 88.365 132.495 88.595 133.635 ;
        RECT 88.805 132.495 89.095 133.660 ;
        RECT 111.805 133.585 113.015 134.105 ;
        RECT 90.075 132.495 90.360 133.295 ;
        RECT 91.480 132.495 91.810 133.185 ;
        RECT 92.480 132.495 92.900 132.875 ;
        RECT 94.180 132.495 94.510 132.875 ;
        RECT 95.030 132.495 95.410 132.875 ;
        RECT 97.055 132.495 97.385 132.995 ;
        RECT 97.995 132.495 98.325 132.995 ;
        RECT 99.735 132.495 100.020 133.295 ;
        RECT 101.140 132.495 101.470 133.185 ;
        RECT 102.140 132.495 102.560 132.875 ;
        RECT 103.840 132.495 104.170 132.875 ;
        RECT 104.690 132.495 105.070 132.875 ;
        RECT 106.715 132.495 107.045 132.995 ;
        RECT 107.655 132.495 107.985 132.995 ;
        RECT 110.415 132.495 110.695 133.295 ;
        RECT 111.805 132.495 114.395 133.585 ;
        RECT 114.565 132.495 114.855 133.660 ;
        RECT 115.485 133.585 117.175 134.105 ;
        RECT 115.485 132.495 118.995 133.585 ;
        RECT 119.605 132.495 119.935 133.255 ;
        RECT 122.600 132.930 122.950 134.180 ;
        RECT 126.525 133.585 127.045 134.125 ;
        RECT 121.010 132.495 126.355 132.930 ;
        RECT 126.525 132.495 127.735 133.585 ;
        RECT 14.660 132.325 127.820 132.495 ;
        RECT 14.745 131.235 15.955 132.325 ;
        RECT 15.435 130.695 15.955 131.235 ;
        RECT 16.585 131.235 20.095 132.325 ;
        RECT 21.015 131.565 21.185 132.325 ;
        RECT 16.585 130.715 18.275 131.235 ;
        RECT 23.555 131.185 23.725 132.325 ;
        RECT 24.405 131.160 24.695 132.325 ;
        RECT 24.870 131.890 30.215 132.325 ;
        RECT 26.460 130.640 26.810 131.890 ;
        RECT 31.195 131.525 31.480 132.325 ;
        RECT 32.600 131.635 32.930 132.325 ;
        RECT 33.600 131.945 34.020 132.325 ;
        RECT 35.300 131.945 35.630 132.325 ;
        RECT 36.150 131.945 36.530 132.325 ;
        RECT 38.175 131.825 38.505 132.325 ;
        RECT 39.115 131.825 39.445 132.325 ;
        RECT 40.485 131.565 40.815 132.325 ;
        RECT 41.425 131.235 42.635 132.325 ;
        RECT 43.005 131.655 43.285 132.325 ;
        RECT 43.955 131.605 44.285 132.325 ;
        RECT 45.305 131.655 45.585 132.325 ;
        RECT 46.255 131.605 46.585 132.325 ;
        RECT 47.405 131.235 49.995 132.325 ;
        RECT 41.425 130.695 41.945 131.235 ;
        RECT 47.405 130.715 48.615 131.235 ;
        RECT 50.165 131.160 50.455 132.325 ;
        RECT 50.625 131.235 54.135 132.325 ;
        RECT 54.310 131.890 59.655 132.325 ;
        RECT 59.830 131.890 65.175 132.325 ;
        RECT 50.625 130.715 52.315 131.235 ;
        RECT 55.900 130.640 56.250 131.890 ;
        RECT 61.420 130.640 61.770 131.890 ;
        RECT 66.095 131.565 66.265 132.325 ;
        RECT 68.635 131.185 68.805 132.325 ;
        RECT 69.950 131.900 70.285 132.325 ;
        RECT 70.845 131.545 71.175 132.325 ;
        RECT 72.435 131.605 72.765 132.325 ;
        RECT 73.435 131.655 73.715 132.325 ;
        RECT 74.525 131.545 74.855 132.325 ;
        RECT 75.415 131.900 75.750 132.325 ;
        RECT 75.925 131.160 76.215 132.325 ;
        RECT 76.845 131.235 78.515 132.325 ;
        RECT 79.335 131.605 79.665 132.325 ;
        RECT 80.335 131.655 80.615 132.325 ;
        RECT 80.985 131.235 82.195 132.325 ;
        RECT 82.370 131.890 87.715 132.325 ;
        RECT 76.845 130.715 77.595 131.235 ;
        RECT 80.985 130.695 81.505 131.235 ;
        RECT 83.960 130.640 84.310 131.890 ;
        RECT 87.925 131.185 88.155 132.325 ;
        RECT 88.825 131.185 89.035 132.325 ;
        RECT 90.015 131.565 90.185 132.325 ;
        RECT 92.555 131.185 92.725 132.325 ;
        RECT 94.305 131.565 94.635 132.325 ;
        RECT 95.685 131.565 96.015 132.325 ;
        RECT 96.625 131.235 97.835 132.325 ;
        RECT 98.485 131.525 98.765 132.325 ;
        RECT 96.625 130.695 97.145 131.235 ;
        RECT 101.685 131.160 101.975 132.325 ;
        RECT 102.145 131.235 103.815 132.325 ;
        RECT 105.815 131.525 106.095 132.325 ;
        RECT 106.745 131.235 110.255 132.325 ;
        RECT 111.075 131.605 111.405 132.325 ;
        RECT 112.075 131.655 112.355 132.325 ;
        RECT 112.725 131.235 115.315 132.325 ;
        RECT 115.490 131.890 120.835 132.325 ;
        RECT 121.010 131.890 126.355 132.325 ;
        RECT 102.145 130.715 102.895 131.235 ;
        RECT 106.745 130.715 108.435 131.235 ;
        RECT 112.725 130.715 113.935 131.235 ;
        RECT 117.080 130.640 117.430 131.890 ;
        RECT 122.600 130.640 122.950 131.890 ;
        RECT 126.525 131.235 127.735 132.325 ;
        RECT 126.525 130.695 127.045 131.235 ;
        RECT 15.435 128.145 15.955 128.685 ;
        RECT 14.745 127.055 15.955 128.145 ;
        RECT 26.705 128.145 27.225 128.685 ;
        RECT 17.855 127.055 18.140 127.855 ;
        RECT 19.260 127.055 19.590 127.745 ;
        RECT 20.260 127.055 20.680 127.435 ;
        RECT 21.960 127.055 22.290 127.435 ;
        RECT 22.810 127.055 23.190 127.435 ;
        RECT 24.835 127.055 25.165 127.555 ;
        RECT 25.775 127.055 26.105 127.555 ;
        RECT 26.705 127.055 27.915 128.145 ;
        RECT 29.680 127.490 30.030 128.740 ;
        RECT 28.090 127.055 33.435 127.490 ;
        RECT 33.645 127.055 33.875 128.195 ;
        RECT 34.545 127.055 34.755 128.195 ;
        RECT 35.185 127.055 35.465 127.725 ;
        RECT 36.135 127.055 36.465 127.775 ;
        RECT 37.285 127.055 37.575 128.220 ;
        RECT 38.205 128.145 39.415 128.665 ;
        RECT 38.205 127.055 40.795 128.145 ;
        RECT 42.560 127.490 42.910 128.740 ;
        RECT 40.970 127.055 46.315 127.490 ;
        RECT 46.685 127.055 46.965 127.725 ;
        RECT 47.635 127.055 47.965 127.775 ;
        RECT 50.840 127.490 51.190 128.740 ;
        RECT 49.250 127.055 54.595 127.490 ;
        RECT 55.515 127.055 55.685 127.815 ;
        RECT 58.055 127.055 58.225 128.195 ;
        RECT 60.285 128.145 61.495 128.665 ;
        RECT 59.345 127.055 59.675 127.815 ;
        RECT 60.285 127.055 62.875 128.145 ;
        RECT 63.045 127.055 63.335 128.220 ;
        RECT 63.505 128.145 64.025 128.685 ;
        RECT 63.505 127.055 64.715 128.145 ;
        RECT 65.695 127.055 65.980 127.855 ;
        RECT 67.100 127.055 67.430 127.745 ;
        RECT 68.100 127.055 68.520 127.435 ;
        RECT 69.800 127.055 70.130 127.435 ;
        RECT 70.650 127.055 71.030 127.435 ;
        RECT 72.675 127.055 73.005 127.555 ;
        RECT 73.615 127.055 73.945 127.555 ;
        RECT 74.745 127.055 75.025 127.725 ;
        RECT 75.695 127.055 76.025 127.775 ;
        RECT 77.045 127.055 77.325 127.725 ;
        RECT 77.995 127.055 78.325 127.775 ;
        RECT 79.895 127.055 80.065 127.815 ;
        RECT 82.435 127.055 82.605 128.195 ;
        RECT 86.045 128.145 87.255 128.665 ;
        RECT 83.935 127.055 84.265 127.775 ;
        RECT 84.935 127.055 85.215 127.725 ;
        RECT 86.045 127.055 88.635 128.145 ;
        RECT 88.805 127.055 89.095 128.220 ;
        RECT 101.685 128.145 102.895 128.665 ;
        RECT 90.535 127.055 90.820 127.855 ;
        RECT 91.940 127.055 92.270 127.745 ;
        RECT 92.940 127.055 93.360 127.435 ;
        RECT 94.640 127.055 94.970 127.435 ;
        RECT 95.490 127.055 95.870 127.435 ;
        RECT 97.515 127.055 97.845 127.555 ;
        RECT 98.455 127.055 98.785 127.555 ;
        RECT 99.585 127.055 99.865 127.725 ;
        RECT 100.535 127.055 100.865 127.775 ;
        RECT 101.685 127.055 104.275 128.145 ;
        RECT 105.095 127.055 105.425 127.775 ;
        RECT 106.095 127.055 106.375 127.725 ;
        RECT 107.395 127.055 107.725 127.775 ;
        RECT 108.395 127.055 108.675 127.725 ;
        RECT 109.695 127.055 110.025 127.775 ;
        RECT 110.695 127.055 110.975 127.725 ;
        RECT 111.860 127.055 112.145 127.925 ;
        RECT 112.750 127.055 113.005 127.515 ;
        RECT 113.605 127.055 113.915 127.855 ;
        RECT 114.565 127.055 114.855 128.220 ;
        RECT 115.675 127.055 116.005 127.775 ;
        RECT 116.675 127.055 116.955 127.725 ;
        RECT 118.285 127.055 118.515 128.195 ;
        RECT 119.185 127.055 119.395 128.195 ;
        RECT 121.465 128.145 121.985 128.685 ;
        RECT 122.845 128.145 124.535 128.665 ;
        RECT 126.525 128.145 127.045 128.685 ;
        RECT 120.525 127.055 120.855 127.815 ;
        RECT 121.465 127.055 122.675 128.145 ;
        RECT 122.845 127.055 126.355 128.145 ;
        RECT 126.525 127.055 127.735 128.145 ;
        RECT 14.660 126.885 127.820 127.055 ;
        RECT 14.745 125.795 15.955 126.885 ;
        RECT 15.435 125.255 15.955 125.795 ;
        RECT 17.045 125.795 20.555 126.885 ;
        RECT 17.045 125.275 18.735 125.795 ;
        RECT 20.785 125.745 20.995 126.885 ;
        RECT 21.665 125.745 21.895 126.885 ;
        RECT 23.465 126.125 23.795 126.885 ;
        RECT 24.405 125.720 24.695 126.885 ;
        RECT 24.865 125.795 26.075 126.885 ;
        RECT 24.865 125.255 25.385 125.795 ;
        RECT 26.755 125.745 26.925 126.885 ;
        RECT 29.295 126.125 29.465 126.885 ;
        RECT 30.385 125.795 32.975 126.885 ;
        RECT 33.895 126.125 34.065 126.885 ;
        RECT 30.385 125.275 31.595 125.795 ;
        RECT 36.435 125.745 36.605 126.885 ;
        RECT 37.485 126.215 37.765 126.885 ;
        RECT 38.435 126.165 38.765 126.885 ;
        RECT 40.705 126.215 40.985 126.885 ;
        RECT 41.655 126.165 41.985 126.885 ;
        RECT 43.005 126.215 43.285 126.885 ;
        RECT 43.955 126.165 44.285 126.885 ;
        RECT 45.755 126.165 46.085 126.885 ;
        RECT 46.755 126.215 47.035 126.885 ;
        RECT 47.460 126.015 47.745 126.885 ;
        RECT 48.350 126.425 48.605 126.885 ;
        RECT 49.205 126.085 49.515 126.885 ;
        RECT 50.165 125.720 50.455 126.885 ;
        RECT 51.095 126.075 51.390 126.885 ;
        RECT 51.990 126.075 52.250 126.885 ;
        RECT 52.850 126.880 59.125 126.885 ;
        RECT 52.850 126.085 53.110 126.880 ;
        RECT 53.710 126.155 53.970 126.880 ;
        RECT 54.570 126.155 54.830 126.880 ;
        RECT 55.430 126.155 55.690 126.880 ;
        RECT 56.290 126.155 56.535 126.880 ;
        RECT 57.150 126.155 57.395 126.880 ;
        RECT 58.010 126.155 58.255 126.880 ;
        RECT 58.870 126.155 59.125 126.880 ;
        RECT 59.755 126.140 60.025 126.885 ;
        RECT 61.035 126.125 61.205 126.885 ;
        RECT 63.575 125.745 63.745 126.885 ;
        RECT 64.885 125.795 68.395 126.885 ;
        RECT 64.885 125.275 66.575 125.795 ;
        RECT 68.625 125.745 68.835 126.885 ;
        RECT 69.505 125.745 69.735 126.885 ;
        RECT 70.385 126.125 70.715 126.885 ;
        RECT 71.325 125.795 72.535 126.885 ;
        RECT 73.185 126.085 73.495 126.885 ;
        RECT 74.095 126.425 74.350 126.885 ;
        RECT 74.955 126.015 75.240 126.885 ;
        RECT 71.325 125.255 71.845 125.795 ;
        RECT 75.925 125.720 76.215 126.885 ;
        RECT 77.195 126.085 77.480 126.885 ;
        RECT 78.600 126.195 78.930 126.885 ;
        RECT 79.600 126.505 80.020 126.885 ;
        RECT 81.300 126.505 81.630 126.885 ;
        RECT 82.150 126.505 82.530 126.885 ;
        RECT 84.175 126.385 84.505 126.885 ;
        RECT 85.115 126.385 85.445 126.885 ;
        RECT 86.155 126.085 86.325 126.885 ;
        RECT 86.995 126.085 87.165 126.885 ;
        RECT 87.835 126.085 88.005 126.885 ;
        RECT 88.675 126.085 88.845 126.885 ;
        RECT 89.515 126.085 89.685 126.885 ;
        RECT 90.355 126.085 90.525 126.885 ;
        RECT 91.195 126.085 91.365 126.885 ;
        RECT 92.035 126.085 92.205 126.885 ;
        RECT 92.875 126.085 93.045 126.885 ;
        RECT 93.715 126.085 93.885 126.885 ;
        RECT 94.555 126.085 94.725 126.885 ;
        RECT 95.395 126.035 95.565 126.885 ;
        RECT 96.235 126.035 96.405 126.885 ;
        RECT 98.005 125.795 101.515 126.885 ;
        RECT 98.005 125.275 99.695 125.795 ;
        RECT 101.685 125.720 101.975 126.885 ;
        RECT 102.145 125.795 103.355 126.885 ;
        RECT 103.525 125.795 107.035 126.885 ;
        RECT 107.955 126.125 108.125 126.885 ;
        RECT 102.145 125.255 102.665 125.795 ;
        RECT 103.525 125.275 105.215 125.795 ;
        RECT 110.495 125.745 110.665 126.885 ;
        RECT 112.095 126.125 112.265 126.885 ;
        RECT 114.635 125.745 114.805 126.885 ;
        RECT 116.295 126.085 116.580 126.885 ;
        RECT 117.700 126.195 118.030 126.885 ;
        RECT 118.700 126.505 119.120 126.885 ;
        RECT 120.400 126.505 120.730 126.885 ;
        RECT 121.250 126.505 121.630 126.885 ;
        RECT 123.275 126.385 123.605 126.885 ;
        RECT 124.215 126.385 124.545 126.885 ;
        RECT 125.145 125.795 126.355 126.885 ;
        RECT 126.525 125.795 127.735 126.885 ;
        RECT 125.145 125.255 125.665 125.795 ;
        RECT 126.525 125.255 127.045 125.795 ;
        RECT 15.435 122.705 15.955 123.245 ;
        RECT 14.745 121.615 15.955 122.705 ;
        RECT 26.245 122.705 26.995 123.225 ;
        RECT 17.055 121.615 17.350 122.425 ;
        RECT 17.950 121.615 18.210 122.425 ;
        RECT 18.810 121.620 19.070 122.415 ;
        RECT 19.670 121.620 19.930 122.345 ;
        RECT 20.530 121.620 20.790 122.345 ;
        RECT 21.390 121.620 21.650 122.345 ;
        RECT 22.250 121.620 22.495 122.345 ;
        RECT 23.110 121.620 23.355 122.345 ;
        RECT 23.970 121.620 24.215 122.345 ;
        RECT 24.830 121.620 25.085 122.345 ;
        RECT 18.810 121.615 25.085 121.620 ;
        RECT 25.715 121.615 25.985 122.360 ;
        RECT 26.245 121.615 27.915 122.705 ;
        RECT 28.175 121.615 28.445 122.360 ;
        RECT 29.075 121.620 29.330 122.345 ;
        RECT 29.945 121.620 30.190 122.345 ;
        RECT 30.805 121.620 31.050 122.345 ;
        RECT 31.665 121.620 31.910 122.345 ;
        RECT 32.510 121.620 32.770 122.345 ;
        RECT 33.370 121.620 33.630 122.345 ;
        RECT 34.230 121.620 34.490 122.345 ;
        RECT 35.090 121.620 35.350 122.415 ;
        RECT 29.075 121.615 35.350 121.620 ;
        RECT 35.950 121.615 36.210 122.425 ;
        RECT 36.810 121.615 37.105 122.425 ;
        RECT 37.285 121.615 37.575 122.780 ;
        RECT 38.495 121.615 38.665 122.375 ;
        RECT 41.035 121.615 41.205 122.755 ;
        RECT 43.480 122.050 43.830 123.300 ;
        RECT 49.000 122.050 49.350 123.300 ;
        RECT 41.890 121.615 47.235 122.050 ;
        RECT 47.410 121.615 52.755 122.050 ;
        RECT 53.735 121.615 54.020 122.415 ;
        RECT 55.140 121.615 55.470 122.305 ;
        RECT 56.140 121.615 56.560 121.995 ;
        RECT 57.840 121.615 58.170 121.995 ;
        RECT 58.690 121.615 59.070 121.995 ;
        RECT 60.715 121.615 61.045 122.115 ;
        RECT 61.655 121.615 61.985 122.115 ;
        RECT 63.045 121.615 63.335 122.780 ;
        RECT 64.255 121.615 64.425 122.375 ;
        RECT 66.795 121.615 66.965 122.755 ;
        RECT 67.645 122.705 68.855 123.225 ;
        RECT 67.645 121.615 70.235 122.705 ;
        RECT 72.000 122.050 72.350 123.300 ;
        RECT 77.520 122.050 77.870 123.300 ;
        RECT 70.410 121.615 75.755 122.050 ;
        RECT 75.930 121.615 81.275 122.050 ;
        RECT 81.505 121.615 81.715 122.755 ;
        RECT 82.385 121.615 82.615 122.755 ;
        RECT 85.125 122.705 86.815 123.225 ;
        RECT 83.725 121.615 84.055 122.375 ;
        RECT 85.125 121.615 88.635 122.705 ;
        RECT 88.805 121.615 89.095 122.780 ;
        RECT 98.465 122.705 98.985 123.245 ;
        RECT 89.275 121.615 89.570 122.425 ;
        RECT 90.170 121.615 90.430 122.425 ;
        RECT 91.030 121.620 91.290 122.415 ;
        RECT 91.890 121.620 92.150 122.345 ;
        RECT 92.750 121.620 93.010 122.345 ;
        RECT 93.610 121.620 93.870 122.345 ;
        RECT 94.470 121.620 94.715 122.345 ;
        RECT 95.330 121.620 95.575 122.345 ;
        RECT 96.190 121.620 96.435 122.345 ;
        RECT 97.050 121.620 97.305 122.345 ;
        RECT 91.030 121.615 97.305 121.620 ;
        RECT 97.935 121.615 98.205 122.360 ;
        RECT 98.465 121.615 99.675 122.705 ;
        RECT 101.440 122.050 101.790 123.300 ;
        RECT 99.850 121.615 105.195 122.050 ;
        RECT 105.375 121.615 105.670 122.425 ;
        RECT 106.270 121.615 106.530 122.425 ;
        RECT 107.130 121.620 107.390 122.415 ;
        RECT 107.990 121.620 108.250 122.345 ;
        RECT 108.850 121.620 109.110 122.345 ;
        RECT 109.710 121.620 109.970 122.345 ;
        RECT 110.570 121.620 110.815 122.345 ;
        RECT 111.430 121.620 111.675 122.345 ;
        RECT 112.290 121.620 112.535 122.345 ;
        RECT 113.150 121.620 113.405 122.345 ;
        RECT 107.130 121.615 113.405 121.620 ;
        RECT 114.035 121.615 114.305 122.360 ;
        RECT 114.565 121.615 114.855 122.780 ;
        RECT 125.145 122.705 125.665 123.245 ;
        RECT 126.525 122.705 127.045 123.245 ;
        RECT 116.295 121.615 116.580 122.415 ;
        RECT 117.700 121.615 118.030 122.305 ;
        RECT 118.700 121.615 119.120 121.995 ;
        RECT 120.400 121.615 120.730 121.995 ;
        RECT 121.250 121.615 121.630 121.995 ;
        RECT 123.275 121.615 123.605 122.115 ;
        RECT 124.215 121.615 124.545 122.115 ;
        RECT 125.145 121.615 126.355 122.705 ;
        RECT 126.525 121.615 127.735 122.705 ;
        RECT 14.660 121.445 127.820 121.615 ;
        RECT 14.745 120.355 15.955 121.445 ;
        RECT 15.435 119.815 15.955 120.355 ;
        RECT 16.585 120.355 20.095 121.445 ;
        RECT 21.015 120.685 21.185 121.445 ;
        RECT 16.585 119.835 18.275 120.355 ;
        RECT 23.555 120.305 23.725 121.445 ;
        RECT 24.405 120.280 24.695 121.445 ;
        RECT 26.225 120.685 26.555 121.445 ;
        RECT 27.625 120.355 29.295 121.445 ;
        RECT 27.625 119.835 28.375 120.355 ;
        RECT 29.505 120.305 29.735 121.445 ;
        RECT 30.405 120.305 30.615 121.445 ;
        RECT 30.885 120.305 31.115 121.445 ;
        RECT 31.785 120.305 31.995 121.445 ;
        RECT 33.035 120.645 33.320 121.445 ;
        RECT 34.440 120.755 34.770 121.445 ;
        RECT 35.440 121.065 35.860 121.445 ;
        RECT 37.140 121.065 37.470 121.445 ;
        RECT 37.990 121.065 38.370 121.445 ;
        RECT 40.015 120.945 40.345 121.445 ;
        RECT 40.955 120.945 41.285 121.445 ;
        RECT 42.635 120.685 42.805 121.445 ;
        RECT 45.175 120.305 45.345 121.445 ;
        RECT 46.775 120.685 46.945 121.445 ;
        RECT 49.315 120.305 49.485 121.445 ;
        RECT 50.165 120.280 50.455 121.445 ;
        RECT 50.665 120.305 50.895 121.445 ;
        RECT 51.565 120.305 51.775 121.445 ;
        RECT 52.005 120.355 53.215 121.445 ;
        RECT 52.005 119.815 52.525 120.355 ;
        RECT 53.535 120.295 53.865 121.445 ;
        RECT 54.375 120.645 54.705 121.445 ;
        RECT 55.225 120.645 55.465 121.445 ;
        RECT 56.735 120.275 57.065 121.445 ;
        RECT 57.795 120.275 58.125 121.445 ;
        RECT 58.855 120.305 59.185 121.445 ;
        RECT 60.175 120.645 60.460 121.445 ;
        RECT 61.580 120.755 61.910 121.445 ;
        RECT 62.580 121.065 63.000 121.445 ;
        RECT 64.280 121.065 64.610 121.445 ;
        RECT 65.130 121.065 65.510 121.445 ;
        RECT 67.155 120.945 67.485 121.445 ;
        RECT 68.095 120.945 68.425 121.445 ;
        RECT 69.465 120.685 69.795 121.445 ;
        RECT 70.865 120.355 74.375 121.445 ;
        RECT 70.865 119.835 72.555 120.355 ;
        RECT 74.585 120.305 74.815 121.445 ;
        RECT 75.485 120.305 75.695 121.445 ;
        RECT 75.925 120.280 76.215 121.445 ;
        RECT 77.595 120.685 77.765 121.445 ;
        RECT 80.135 120.305 80.305 121.445 ;
        RECT 81.425 120.685 81.755 121.445 ;
        RECT 82.425 120.305 82.635 121.445 ;
        RECT 83.305 120.305 83.535 121.445 ;
        RECT 84.645 120.685 84.975 121.445 ;
        RECT 85.585 120.355 89.095 121.445 ;
        RECT 85.585 119.835 87.275 120.355 ;
        RECT 89.305 120.305 89.535 121.445 ;
        RECT 90.205 120.305 90.415 121.445 ;
        RECT 90.685 120.305 90.915 121.445 ;
        RECT 91.585 120.305 91.795 121.445 ;
        RECT 92.835 120.645 93.120 121.445 ;
        RECT 94.240 120.755 94.570 121.445 ;
        RECT 95.240 121.065 95.660 121.445 ;
        RECT 96.940 121.065 97.270 121.445 ;
        RECT 97.790 121.065 98.170 121.445 ;
        RECT 99.815 120.945 100.145 121.445 ;
        RECT 100.755 120.945 101.085 121.445 ;
        RECT 101.685 120.280 101.975 121.445 ;
        RECT 102.585 120.685 102.915 121.445 ;
        RECT 103.565 120.305 103.795 121.445 ;
        RECT 104.465 120.305 104.675 121.445 ;
        RECT 105.655 120.685 105.825 121.445 ;
        RECT 108.195 120.305 108.365 121.445 ;
        RECT 109.855 120.645 110.140 121.445 ;
        RECT 111.260 120.755 111.590 121.445 ;
        RECT 112.260 121.065 112.680 121.445 ;
        RECT 113.960 121.065 114.290 121.445 ;
        RECT 114.810 121.065 115.190 121.445 ;
        RECT 116.835 120.945 117.165 121.445 ;
        RECT 117.775 120.945 118.105 121.445 ;
        RECT 118.745 120.305 118.975 121.445 ;
        RECT 119.645 120.305 119.855 121.445 ;
        RECT 120.985 120.685 121.315 121.445 ;
        RECT 122.845 120.355 126.355 121.445 ;
        RECT 126.525 120.355 127.735 121.445 ;
        RECT 122.845 119.835 124.535 120.355 ;
        RECT 126.525 119.815 127.045 120.355 ;
        RECT 15.435 117.265 15.955 117.805 ;
        RECT 14.745 116.175 15.955 117.265 ;
        RECT 16.125 117.265 16.875 117.785 ;
        RECT 16.125 116.175 17.795 117.265 ;
        RECT 18.775 116.175 19.060 116.975 ;
        RECT 20.180 116.175 20.510 116.865 ;
        RECT 21.180 116.175 21.600 116.555 ;
        RECT 22.880 116.175 23.210 116.555 ;
        RECT 23.730 116.175 24.110 116.555 ;
        RECT 25.755 116.175 26.085 116.675 ;
        RECT 26.695 116.175 27.025 116.675 ;
        RECT 28.435 116.175 28.720 116.975 ;
        RECT 29.840 116.175 30.170 116.865 ;
        RECT 30.840 116.175 31.260 116.555 ;
        RECT 32.540 116.175 32.870 116.555 ;
        RECT 33.390 116.175 33.770 116.555 ;
        RECT 35.415 116.175 35.745 116.675 ;
        RECT 36.355 116.175 36.685 116.675 ;
        RECT 37.285 116.175 37.575 117.340 ;
        RECT 38.555 116.175 38.840 116.975 ;
        RECT 39.960 116.175 40.290 116.865 ;
        RECT 40.960 116.175 41.380 116.555 ;
        RECT 42.660 116.175 42.990 116.555 ;
        RECT 43.510 116.175 43.890 116.555 ;
        RECT 45.535 116.175 45.865 116.675 ;
        RECT 46.475 116.175 46.805 116.675 ;
        RECT 48.215 116.175 48.500 116.975 ;
        RECT 49.620 116.175 49.950 116.865 ;
        RECT 50.620 116.175 51.040 116.555 ;
        RECT 52.320 116.175 52.650 116.555 ;
        RECT 53.170 116.175 53.550 116.555 ;
        RECT 55.195 116.175 55.525 116.675 ;
        RECT 56.135 116.175 56.465 116.675 ;
        RECT 57.125 116.175 57.335 117.315 ;
        RECT 58.005 116.175 58.235 117.315 ;
        RECT 58.905 117.265 60.115 117.785 ;
        RECT 58.905 116.175 61.495 117.265 ;
        RECT 61.705 116.175 61.935 117.315 ;
        RECT 62.605 116.175 62.815 117.315 ;
        RECT 63.045 116.175 63.335 117.340 ;
        RECT 64.315 116.175 64.600 116.975 ;
        RECT 65.720 116.175 66.050 116.865 ;
        RECT 66.720 116.175 67.140 116.555 ;
        RECT 68.420 116.175 68.750 116.555 ;
        RECT 69.270 116.175 69.650 116.555 ;
        RECT 71.295 116.175 71.625 116.675 ;
        RECT 72.235 116.175 72.565 116.675 ;
        RECT 73.975 116.175 74.260 116.975 ;
        RECT 75.380 116.175 75.710 116.865 ;
        RECT 76.380 116.175 76.800 116.555 ;
        RECT 78.080 116.175 78.410 116.555 ;
        RECT 78.930 116.175 79.310 116.555 ;
        RECT 80.955 116.175 81.285 116.675 ;
        RECT 81.895 116.175 82.225 116.675 ;
        RECT 83.335 116.175 83.505 117.315 ;
        RECT 85.875 116.175 86.045 116.935 ;
        RECT 87.465 116.175 87.695 117.315 ;
        RECT 88.365 116.175 88.575 117.315 ;
        RECT 88.805 116.175 89.095 117.340 ;
        RECT 90.075 116.175 90.360 116.975 ;
        RECT 91.480 116.175 91.810 116.865 ;
        RECT 92.480 116.175 92.900 116.555 ;
        RECT 94.180 116.175 94.510 116.555 ;
        RECT 95.030 116.175 95.410 116.555 ;
        RECT 97.055 116.175 97.385 116.675 ;
        RECT 97.995 116.175 98.325 116.675 ;
        RECT 99.365 116.175 99.695 116.935 ;
        RECT 102.035 116.175 102.320 116.975 ;
        RECT 103.440 116.175 103.770 116.865 ;
        RECT 104.440 116.175 104.860 116.555 ;
        RECT 106.140 116.175 106.470 116.555 ;
        RECT 106.990 116.175 107.370 116.555 ;
        RECT 109.015 116.175 109.345 116.675 ;
        RECT 109.955 116.175 110.285 116.675 ;
        RECT 111.325 116.175 111.655 116.935 ;
        RECT 112.785 116.175 112.995 117.315 ;
        RECT 113.665 116.175 113.895 117.315 ;
        RECT 114.565 116.175 114.855 117.340 ;
        RECT 126.525 117.265 127.045 117.805 ;
        RECT 115.925 116.175 116.255 116.935 ;
        RECT 117.335 116.175 117.630 116.985 ;
        RECT 118.230 116.175 118.490 116.985 ;
        RECT 119.090 116.180 119.350 116.975 ;
        RECT 119.950 116.180 120.210 116.905 ;
        RECT 120.810 116.180 121.070 116.905 ;
        RECT 121.670 116.180 121.930 116.905 ;
        RECT 122.530 116.180 122.775 116.905 ;
        RECT 123.390 116.180 123.635 116.905 ;
        RECT 124.250 116.180 124.495 116.905 ;
        RECT 125.110 116.180 125.365 116.905 ;
        RECT 119.090 116.175 125.365 116.180 ;
        RECT 125.995 116.175 126.265 116.920 ;
        RECT 126.525 116.175 127.735 117.265 ;
        RECT 14.660 116.005 127.820 116.175 ;
        RECT 14.745 114.915 15.955 116.005 ;
        RECT 15.435 114.375 15.955 114.915 ;
        RECT 16.585 114.915 20.095 116.005 ;
        RECT 16.585 114.395 18.275 114.915 ;
        RECT 20.305 114.865 20.535 116.005 ;
        RECT 21.205 114.865 21.415 116.005 ;
        RECT 21.705 114.865 21.915 116.005 ;
        RECT 22.585 114.865 22.815 116.005 ;
        RECT 23.465 115.245 23.795 116.005 ;
        RECT 24.405 114.840 24.695 116.005 ;
        RECT 24.875 115.195 25.170 116.005 ;
        RECT 25.770 115.195 26.030 116.005 ;
        RECT 26.630 116.000 32.905 116.005 ;
        RECT 26.630 115.205 26.890 116.000 ;
        RECT 27.490 115.275 27.750 116.000 ;
        RECT 28.350 115.275 28.610 116.000 ;
        RECT 29.210 115.275 29.470 116.000 ;
        RECT 30.070 115.275 30.315 116.000 ;
        RECT 30.930 115.275 31.175 116.000 ;
        RECT 31.790 115.275 32.035 116.000 ;
        RECT 32.650 115.275 32.905 116.000 ;
        RECT 33.535 115.260 33.805 116.005 ;
        RECT 34.155 115.260 34.425 116.005 ;
        RECT 35.055 116.000 41.330 116.005 ;
        RECT 35.055 115.275 35.310 116.000 ;
        RECT 35.925 115.275 36.170 116.000 ;
        RECT 36.785 115.275 37.030 116.000 ;
        RECT 37.645 115.275 37.890 116.000 ;
        RECT 38.490 115.275 38.750 116.000 ;
        RECT 39.350 115.275 39.610 116.000 ;
        RECT 40.210 115.275 40.470 116.000 ;
        RECT 41.070 115.205 41.330 116.000 ;
        RECT 41.930 115.195 42.190 116.005 ;
        RECT 42.790 115.195 43.085 116.005 ;
        RECT 43.705 115.245 44.035 116.005 ;
        RECT 44.705 114.865 44.915 116.005 ;
        RECT 45.585 114.865 45.815 116.005 ;
        RECT 46.025 114.915 47.695 116.005 ;
        RECT 48.305 115.245 48.635 116.005 ;
        RECT 46.025 114.395 46.775 114.915 ;
        RECT 50.165 114.840 50.455 116.005 ;
        RECT 50.625 114.915 52.295 116.005 ;
        RECT 52.905 115.245 53.235 116.005 ;
        RECT 54.770 115.570 60.115 116.005 ;
        RECT 60.290 115.570 65.635 116.005 ;
        RECT 50.625 114.395 51.375 114.915 ;
        RECT 56.360 114.320 56.710 115.570 ;
        RECT 61.880 114.320 62.230 115.570 ;
        RECT 65.845 114.865 66.075 116.005 ;
        RECT 66.745 114.865 66.955 116.005 ;
        RECT 68.545 115.245 68.875 116.005 ;
        RECT 70.410 115.570 75.755 116.005 ;
        RECT 72.000 114.320 72.350 115.570 ;
        RECT 75.925 114.840 76.215 116.005 ;
        RECT 78.115 115.205 78.400 116.005 ;
        RECT 79.520 115.315 79.850 116.005 ;
        RECT 80.520 115.625 80.940 116.005 ;
        RECT 82.220 115.625 82.550 116.005 ;
        RECT 83.070 115.625 83.450 116.005 ;
        RECT 85.095 115.505 85.425 116.005 ;
        RECT 86.035 115.505 86.365 116.005 ;
        RECT 87.425 114.915 90.935 116.005 ;
        RECT 91.855 115.245 92.025 116.005 ;
        RECT 87.425 114.395 89.115 114.915 ;
        RECT 94.395 114.865 94.565 116.005 ;
        RECT 95.705 114.915 97.375 116.005 ;
        RECT 98.295 115.245 98.465 116.005 ;
        RECT 95.705 114.395 96.455 114.915 ;
        RECT 100.835 114.865 101.005 116.005 ;
        RECT 101.685 114.840 101.975 116.005 ;
        RECT 102.145 114.915 105.655 116.005 ;
        RECT 105.830 115.570 111.175 116.005 ;
        RECT 102.145 114.395 103.835 114.915 ;
        RECT 107.420 114.320 107.770 115.570 ;
        RECT 112.095 115.245 112.265 116.005 ;
        RECT 114.635 114.865 114.805 116.005 ;
        RECT 115.485 114.915 117.155 116.005 ;
        RECT 117.755 115.505 118.085 116.005 ;
        RECT 119.090 115.545 119.340 116.005 ;
        RECT 121.230 115.575 121.560 116.005 ;
        RECT 122.195 115.545 122.565 116.005 ;
        RECT 124.180 115.545 124.430 116.005 ;
        RECT 124.950 115.625 125.280 116.005 ;
        RECT 115.485 114.395 116.235 114.915 ;
        RECT 125.620 114.865 125.925 116.005 ;
        RECT 126.525 114.915 127.735 116.005 ;
        RECT 126.525 114.375 127.045 114.915 ;
        RECT 15.435 111.825 15.955 112.365 ;
        RECT 14.745 110.735 15.955 111.825 ;
        RECT 17.855 110.735 18.140 111.535 ;
        RECT 19.260 110.735 19.590 111.425 ;
        RECT 20.260 110.735 20.680 111.115 ;
        RECT 21.960 110.735 22.290 111.115 ;
        RECT 22.810 110.735 23.190 111.115 ;
        RECT 24.835 110.735 25.165 111.235 ;
        RECT 25.775 110.735 26.105 111.235 ;
        RECT 27.135 110.735 27.465 111.235 ;
        RECT 28.470 110.735 28.720 111.195 ;
        RECT 30.610 110.735 30.940 111.165 ;
        RECT 31.575 110.735 31.945 111.195 ;
        RECT 33.560 110.735 33.810 111.195 ;
        RECT 34.330 110.735 34.660 111.115 ;
        RECT 35.000 110.735 35.305 111.875 ;
        RECT 36.345 110.735 36.675 111.495 ;
        RECT 37.285 110.735 37.575 111.900 ;
        RECT 46.945 111.825 47.465 112.365 ;
        RECT 48.325 111.825 50.015 112.345 ;
        RECT 37.755 110.735 38.050 111.545 ;
        RECT 38.650 110.735 38.910 111.545 ;
        RECT 39.510 110.740 39.770 111.535 ;
        RECT 40.370 110.740 40.630 111.465 ;
        RECT 41.230 110.740 41.490 111.465 ;
        RECT 42.090 110.740 42.350 111.465 ;
        RECT 42.950 110.740 43.195 111.465 ;
        RECT 43.810 110.740 44.055 111.465 ;
        RECT 44.670 110.740 44.915 111.465 ;
        RECT 45.530 110.740 45.785 111.465 ;
        RECT 39.510 110.735 45.785 110.740 ;
        RECT 46.415 110.735 46.685 111.480 ;
        RECT 46.945 110.735 48.155 111.825 ;
        RECT 48.325 110.735 51.835 111.825 ;
        RECT 53.600 111.170 53.950 112.420 ;
        RECT 59.120 111.170 59.470 112.420 ;
        RECT 52.010 110.735 57.355 111.170 ;
        RECT 57.530 110.735 62.875 111.170 ;
        RECT 63.045 110.735 63.335 111.900 ;
        RECT 64.425 111.825 66.115 112.345 ;
        RECT 64.425 110.735 67.935 111.825 ;
        RECT 69.700 111.170 70.050 112.420 ;
        RECT 75.220 111.170 75.570 112.420 ;
        RECT 68.110 110.735 73.455 111.170 ;
        RECT 73.630 110.735 78.975 111.170 ;
        RECT 79.185 110.735 79.415 111.875 ;
        RECT 80.085 110.735 80.295 111.875 ;
        RECT 80.675 110.735 81.005 111.885 ;
        RECT 81.515 110.735 81.845 111.535 ;
        RECT 82.365 110.735 82.605 111.535 ;
        RECT 84.880 111.170 85.230 112.420 ;
        RECT 83.290 110.735 88.635 111.170 ;
        RECT 88.805 110.735 89.095 111.900 ;
        RECT 89.725 111.825 91.415 112.345 ;
        RECT 89.725 110.735 93.235 111.825 ;
        RECT 93.465 110.735 93.675 111.875 ;
        RECT 94.345 110.735 94.575 111.875 ;
        RECT 96.840 111.170 97.190 112.420 ;
        RECT 102.360 111.170 102.710 112.420 ;
        RECT 107.665 111.825 108.185 112.365 ;
        RECT 95.250 110.735 100.595 111.170 ;
        RECT 100.770 110.735 106.115 111.170 ;
        RECT 106.725 110.735 107.055 111.495 ;
        RECT 107.665 110.735 108.875 111.825 ;
        RECT 110.640 111.170 110.990 112.420 ;
        RECT 109.050 110.735 114.395 111.170 ;
        RECT 114.565 110.735 114.855 111.900 ;
        RECT 126.525 111.825 127.045 112.365 ;
        RECT 115.115 110.735 115.385 111.480 ;
        RECT 116.015 110.740 116.270 111.465 ;
        RECT 116.885 110.740 117.130 111.465 ;
        RECT 117.745 110.740 117.990 111.465 ;
        RECT 118.605 110.740 118.850 111.465 ;
        RECT 119.450 110.740 119.710 111.465 ;
        RECT 120.310 110.740 120.570 111.465 ;
        RECT 121.170 110.740 121.430 111.465 ;
        RECT 122.030 110.740 122.290 111.535 ;
        RECT 116.015 110.735 122.290 110.740 ;
        RECT 122.890 110.735 123.150 111.545 ;
        RECT 123.750 110.735 124.045 111.545 ;
        RECT 124.665 110.735 124.995 111.495 ;
        RECT 126.525 110.735 127.735 111.825 ;
        RECT 14.660 110.565 127.820 110.735 ;
        RECT 14.745 109.475 15.955 110.565 ;
        RECT 15.435 108.935 15.955 109.475 ;
        RECT 16.125 109.475 17.335 110.565 ;
        RECT 17.510 110.130 22.855 110.565 ;
        RECT 16.125 108.935 16.645 109.475 ;
        RECT 19.100 108.880 19.450 110.130 ;
        RECT 23.065 109.425 23.295 110.565 ;
        RECT 23.965 109.425 24.175 110.565 ;
        RECT 24.405 109.400 24.695 110.565 ;
        RECT 24.865 109.475 26.075 110.565 ;
        RECT 26.685 109.805 27.015 110.565 ;
        RECT 28.065 109.805 28.395 110.565 ;
        RECT 29.015 109.755 29.310 110.565 ;
        RECT 29.910 109.755 30.170 110.565 ;
        RECT 30.770 110.560 37.045 110.565 ;
        RECT 30.770 109.765 31.030 110.560 ;
        RECT 31.630 109.835 31.890 110.560 ;
        RECT 32.490 109.835 32.750 110.560 ;
        RECT 33.350 109.835 33.610 110.560 ;
        RECT 34.210 109.835 34.455 110.560 ;
        RECT 35.070 109.835 35.315 110.560 ;
        RECT 35.930 109.835 36.175 110.560 ;
        RECT 36.790 109.835 37.045 110.560 ;
        RECT 37.675 109.820 37.945 110.565 ;
        RECT 38.635 110.065 38.965 110.565 ;
        RECT 39.970 110.105 40.220 110.565 ;
        RECT 42.110 110.135 42.440 110.565 ;
        RECT 43.075 110.105 43.445 110.565 ;
        RECT 45.060 110.105 45.310 110.565 ;
        RECT 45.830 110.185 46.160 110.565 ;
        RECT 24.865 108.935 25.385 109.475 ;
        RECT 46.500 109.425 46.805 110.565 ;
        RECT 47.845 109.805 48.175 110.565 ;
        RECT 48.785 109.475 49.995 110.565 ;
        RECT 48.785 108.935 49.305 109.475 ;
        RECT 50.165 109.400 50.455 110.565 ;
        RECT 51.525 109.805 51.855 110.565 ;
        RECT 53.385 109.475 56.895 110.565 ;
        RECT 57.505 109.805 57.835 110.565 ;
        RECT 58.445 109.475 60.115 110.565 ;
        RECT 60.795 109.765 61.035 110.565 ;
        RECT 61.555 109.765 61.885 110.565 ;
        RECT 53.385 108.955 55.075 109.475 ;
        RECT 58.445 108.955 59.195 109.475 ;
        RECT 62.395 109.415 62.725 110.565 ;
        RECT 63.945 109.805 64.275 110.565 ;
        RECT 64.975 109.820 65.245 110.565 ;
        RECT 65.875 110.560 72.150 110.565 ;
        RECT 65.875 109.835 66.130 110.560 ;
        RECT 66.745 109.835 66.990 110.560 ;
        RECT 67.605 109.835 67.850 110.560 ;
        RECT 68.465 109.835 68.710 110.560 ;
        RECT 69.310 109.835 69.570 110.560 ;
        RECT 70.170 109.835 70.430 110.560 ;
        RECT 71.030 109.835 71.290 110.560 ;
        RECT 71.890 109.765 72.150 110.560 ;
        RECT 72.750 109.755 73.010 110.565 ;
        RECT 73.610 109.755 73.905 110.565 ;
        RECT 74.605 109.425 74.815 110.565 ;
        RECT 75.485 109.425 75.715 110.565 ;
        RECT 75.925 109.400 76.215 110.565 ;
        RECT 76.935 109.820 77.205 110.565 ;
        RECT 77.835 110.560 84.110 110.565 ;
        RECT 77.835 109.835 78.090 110.560 ;
        RECT 78.705 109.835 78.950 110.560 ;
        RECT 79.565 109.835 79.810 110.560 ;
        RECT 80.425 109.835 80.670 110.560 ;
        RECT 81.270 109.835 81.530 110.560 ;
        RECT 82.130 109.835 82.390 110.560 ;
        RECT 82.990 109.835 83.250 110.560 ;
        RECT 83.850 109.765 84.110 110.560 ;
        RECT 84.710 109.755 84.970 110.565 ;
        RECT 85.570 109.755 85.865 110.565 ;
        RECT 86.085 109.425 86.315 110.565 ;
        RECT 86.985 109.425 87.195 110.565 ;
        RECT 87.865 109.805 88.195 110.565 ;
        RECT 88.895 109.820 89.165 110.565 ;
        RECT 89.795 110.560 96.070 110.565 ;
        RECT 89.795 109.835 90.050 110.560 ;
        RECT 90.665 109.835 90.910 110.560 ;
        RECT 91.525 109.835 91.770 110.560 ;
        RECT 92.385 109.835 92.630 110.560 ;
        RECT 93.230 109.835 93.490 110.560 ;
        RECT 94.090 109.835 94.350 110.560 ;
        RECT 94.950 109.835 95.210 110.560 ;
        RECT 95.810 109.765 96.070 110.560 ;
        RECT 96.670 109.755 96.930 110.565 ;
        RECT 97.530 109.755 97.825 110.565 ;
        RECT 98.965 109.425 99.195 110.565 ;
        RECT 99.865 109.425 100.075 110.565 ;
        RECT 100.745 109.805 101.075 110.565 ;
        RECT 101.685 109.400 101.975 110.565 ;
        RECT 102.235 109.820 102.505 110.565 ;
        RECT 103.135 110.560 109.410 110.565 ;
        RECT 103.135 109.835 103.390 110.560 ;
        RECT 104.005 109.835 104.250 110.560 ;
        RECT 104.865 109.835 105.110 110.560 ;
        RECT 105.725 109.835 105.970 110.560 ;
        RECT 106.570 109.835 106.830 110.560 ;
        RECT 107.430 109.835 107.690 110.560 ;
        RECT 108.290 109.835 108.550 110.560 ;
        RECT 109.150 109.765 109.410 110.560 ;
        RECT 110.010 109.755 110.270 110.565 ;
        RECT 110.870 109.755 111.165 110.565 ;
        RECT 111.785 109.805 112.115 110.565 ;
        RECT 113.165 109.805 113.495 110.565 ;
        RECT 115.005 109.805 115.335 110.565 ;
        RECT 115.985 109.425 116.215 110.565 ;
        RECT 116.885 109.425 117.095 110.565 ;
        RECT 117.755 109.425 118.060 110.565 ;
        RECT 118.400 110.185 118.730 110.565 ;
        RECT 119.250 110.105 119.500 110.565 ;
        RECT 121.115 110.105 121.485 110.565 ;
        RECT 122.120 110.135 122.450 110.565 ;
        RECT 124.340 110.105 124.590 110.565 ;
        RECT 125.595 110.065 125.925 110.565 ;
        RECT 126.525 109.475 127.735 110.565 ;
        RECT 126.525 108.935 127.045 109.475 ;
        RECT 15.435 106.385 15.955 106.925 ;
        RECT 14.745 105.295 15.955 106.385 ;
        RECT 16.125 106.385 16.645 106.925 ;
        RECT 16.125 105.295 17.335 106.385 ;
        RECT 17.565 105.295 17.775 106.435 ;
        RECT 18.445 105.295 18.675 106.435 ;
        RECT 19.315 105.295 19.620 106.435 ;
        RECT 19.960 105.295 20.290 105.675 ;
        RECT 20.810 105.295 21.060 105.755 ;
        RECT 22.675 105.295 23.045 105.755 ;
        RECT 23.680 105.295 24.010 105.725 ;
        RECT 25.900 105.295 26.150 105.755 ;
        RECT 27.155 105.295 27.485 105.795 ;
        RECT 28.515 105.295 28.820 106.435 ;
        RECT 29.160 105.295 29.490 105.675 ;
        RECT 30.010 105.295 30.260 105.755 ;
        RECT 31.875 105.295 32.245 105.755 ;
        RECT 32.880 105.295 33.210 105.725 ;
        RECT 35.100 105.295 35.350 105.755 ;
        RECT 36.355 105.295 36.685 105.795 ;
        RECT 37.285 105.295 37.575 106.460 ;
        RECT 37.785 105.295 38.015 106.435 ;
        RECT 38.685 105.295 38.895 106.435 ;
        RECT 39.215 105.295 39.485 106.040 ;
        RECT 40.115 105.300 40.370 106.025 ;
        RECT 40.985 105.300 41.230 106.025 ;
        RECT 41.845 105.300 42.090 106.025 ;
        RECT 42.705 105.300 42.950 106.025 ;
        RECT 43.550 105.300 43.810 106.025 ;
        RECT 44.410 105.300 44.670 106.025 ;
        RECT 45.270 105.300 45.530 106.025 ;
        RECT 46.130 105.300 46.390 106.095 ;
        RECT 40.115 105.295 46.390 105.300 ;
        RECT 46.990 105.295 47.250 106.105 ;
        RECT 47.850 105.295 48.145 106.105 ;
        RECT 48.755 105.295 49.060 106.435 ;
        RECT 49.400 105.295 49.730 105.675 ;
        RECT 50.250 105.295 50.500 105.755 ;
        RECT 52.115 105.295 52.485 105.755 ;
        RECT 53.120 105.295 53.450 105.725 ;
        RECT 55.340 105.295 55.590 105.755 ;
        RECT 56.595 105.295 56.925 105.795 ;
        RECT 57.585 105.295 57.795 106.435 ;
        RECT 58.465 105.295 58.695 106.435 ;
        RECT 58.905 106.385 59.425 106.925 ;
        RECT 58.905 105.295 60.115 106.385 ;
        RECT 60.325 105.295 60.555 106.435 ;
        RECT 61.225 105.295 61.435 106.435 ;
        RECT 62.105 105.295 62.435 106.055 ;
        RECT 63.045 105.295 63.335 106.460 ;
        RECT 63.545 105.295 63.775 106.435 ;
        RECT 64.445 105.295 64.655 106.435 ;
        RECT 65.315 105.295 65.620 106.435 ;
        RECT 65.960 105.295 66.290 105.675 ;
        RECT 66.810 105.295 67.060 105.755 ;
        RECT 68.675 105.295 69.045 105.755 ;
        RECT 69.680 105.295 70.010 105.725 ;
        RECT 71.900 105.295 72.150 105.755 ;
        RECT 73.155 105.295 73.485 105.795 ;
        RECT 75.065 105.295 75.275 106.435 ;
        RECT 75.945 105.295 76.175 106.435 ;
        RECT 76.825 105.295 77.155 106.055 ;
        RECT 78.195 105.295 78.500 106.435 ;
        RECT 78.840 105.295 79.170 105.675 ;
        RECT 79.690 105.295 79.940 105.755 ;
        RECT 81.555 105.295 81.925 105.755 ;
        RECT 82.560 105.295 82.890 105.725 ;
        RECT 84.780 105.295 85.030 105.755 ;
        RECT 86.035 105.295 86.365 105.795 ;
        RECT 87.405 105.295 87.735 106.055 ;
        RECT 88.805 105.295 89.095 106.460 ;
        RECT 90.615 105.295 90.920 106.435 ;
        RECT 91.260 105.295 91.590 105.675 ;
        RECT 92.110 105.295 92.360 105.755 ;
        RECT 93.975 105.295 94.345 105.755 ;
        RECT 94.980 105.295 95.310 105.725 ;
        RECT 97.200 105.295 97.450 105.755 ;
        RECT 98.455 105.295 98.785 105.795 ;
        RECT 99.815 105.295 100.120 106.435 ;
        RECT 100.460 105.295 100.790 105.675 ;
        RECT 101.310 105.295 101.560 105.755 ;
        RECT 103.175 105.295 103.545 105.755 ;
        RECT 104.180 105.295 104.510 105.725 ;
        RECT 106.400 105.295 106.650 105.755 ;
        RECT 107.655 105.295 107.985 105.795 ;
        RECT 108.645 105.295 108.855 106.435 ;
        RECT 109.525 105.295 109.755 106.435 ;
        RECT 110.005 105.295 110.235 106.435 ;
        RECT 110.905 105.295 111.115 106.435 ;
        RECT 111.345 106.385 112.095 106.905 ;
        RECT 111.345 105.295 113.015 106.385 ;
        RECT 113.225 105.295 113.455 106.435 ;
        RECT 114.125 105.295 114.335 106.435 ;
        RECT 114.565 105.295 114.855 106.460 ;
        RECT 115.455 105.295 115.760 106.435 ;
        RECT 116.100 105.295 116.430 105.675 ;
        RECT 116.950 105.295 117.200 105.755 ;
        RECT 118.815 105.295 119.185 105.755 ;
        RECT 119.820 105.295 120.150 105.725 ;
        RECT 122.040 105.295 122.290 105.755 ;
        RECT 123.295 105.295 123.625 105.795 ;
        RECT 124.265 105.295 124.495 106.435 ;
        RECT 125.165 105.295 125.375 106.435 ;
        RECT 126.525 106.385 127.045 106.925 ;
        RECT 126.525 105.295 127.735 106.385 ;
        RECT 14.660 105.125 127.820 105.295 ;
        RECT 14.745 104.035 15.955 105.125 ;
        RECT 15.435 103.495 15.955 104.035 ;
        RECT 16.125 104.035 18.715 105.125 ;
        RECT 18.890 104.690 24.235 105.125 ;
        RECT 16.125 103.515 17.335 104.035 ;
        RECT 20.480 103.440 20.830 104.690 ;
        RECT 24.405 103.960 24.695 105.125 ;
        RECT 24.865 104.035 26.075 105.125 ;
        RECT 24.865 103.495 25.385 104.035 ;
        RECT 26.305 103.985 26.515 105.125 ;
        RECT 27.185 103.985 27.415 105.125 ;
        RECT 27.665 103.985 27.895 105.125 ;
        RECT 28.565 103.985 28.775 105.125 ;
        RECT 29.445 104.365 29.775 105.125 ;
        RECT 30.825 104.365 31.155 105.125 ;
        RECT 32.195 103.985 32.500 105.125 ;
        RECT 32.840 104.745 33.170 105.125 ;
        RECT 33.690 104.665 33.940 105.125 ;
        RECT 35.555 104.665 35.925 105.125 ;
        RECT 36.560 104.695 36.890 105.125 ;
        RECT 38.780 104.665 39.030 105.125 ;
        RECT 40.035 104.625 40.365 105.125 ;
        RECT 41.395 103.985 41.700 105.125 ;
        RECT 42.040 104.745 42.370 105.125 ;
        RECT 42.890 104.665 43.140 105.125 ;
        RECT 44.755 104.665 45.125 105.125 ;
        RECT 45.760 104.695 46.090 105.125 ;
        RECT 47.980 104.665 48.230 105.125 ;
        RECT 49.235 104.625 49.565 105.125 ;
        RECT 50.165 103.960 50.455 105.125 ;
        RECT 51.605 103.985 51.815 105.125 ;
        RECT 52.485 103.985 52.715 105.125 ;
        RECT 52.925 104.035 54.135 105.125 ;
        RECT 52.925 103.495 53.445 104.035 ;
        RECT 54.735 103.985 55.040 105.125 ;
        RECT 55.380 104.745 55.710 105.125 ;
        RECT 56.230 104.665 56.480 105.125 ;
        RECT 58.095 104.665 58.465 105.125 ;
        RECT 59.100 104.695 59.430 105.125 ;
        RECT 61.320 104.665 61.570 105.125 ;
        RECT 62.575 104.625 62.905 105.125 ;
        RECT 63.935 103.985 64.240 105.125 ;
        RECT 64.580 104.745 64.910 105.125 ;
        RECT 65.430 104.665 65.680 105.125 ;
        RECT 67.295 104.665 67.665 105.125 ;
        RECT 68.300 104.695 68.630 105.125 ;
        RECT 70.520 104.665 70.770 105.125 ;
        RECT 71.775 104.625 72.105 105.125 ;
        RECT 73.165 104.035 75.755 105.125 ;
        RECT 73.165 103.515 74.375 104.035 ;
        RECT 75.925 103.960 76.215 105.125 ;
        RECT 76.815 103.985 77.120 105.125 ;
        RECT 77.460 104.745 77.790 105.125 ;
        RECT 78.310 104.665 78.560 105.125 ;
        RECT 80.175 104.665 80.545 105.125 ;
        RECT 81.180 104.695 81.510 105.125 ;
        RECT 83.400 104.665 83.650 105.125 ;
        RECT 84.655 104.625 84.985 105.125 ;
        RECT 86.015 103.985 86.320 105.125 ;
        RECT 86.660 104.745 86.990 105.125 ;
        RECT 87.510 104.665 87.760 105.125 ;
        RECT 89.375 104.665 89.745 105.125 ;
        RECT 90.380 104.695 90.710 105.125 ;
        RECT 92.600 104.665 92.850 105.125 ;
        RECT 93.855 104.625 94.185 105.125 ;
        RECT 95.225 104.365 95.555 105.125 ;
        RECT 96.170 104.690 101.515 105.125 ;
        RECT 97.760 103.440 98.110 104.690 ;
        RECT 101.685 103.960 101.975 105.125 ;
        RECT 102.575 104.625 102.905 105.125 ;
        RECT 103.910 104.665 104.160 105.125 ;
        RECT 106.050 104.695 106.380 105.125 ;
        RECT 107.015 104.665 107.385 105.125 ;
        RECT 109.000 104.665 109.250 105.125 ;
        RECT 109.770 104.745 110.100 105.125 ;
        RECT 110.440 103.985 110.745 105.125 ;
        RECT 111.775 103.985 112.080 105.125 ;
        RECT 112.420 104.745 112.750 105.125 ;
        RECT 113.270 104.665 113.520 105.125 ;
        RECT 115.135 104.665 115.505 105.125 ;
        RECT 116.140 104.695 116.470 105.125 ;
        RECT 118.360 104.665 118.610 105.125 ;
        RECT 119.615 104.625 119.945 105.125 ;
        RECT 121.465 104.035 124.975 105.125 ;
        RECT 125.585 104.365 125.915 105.125 ;
        RECT 126.525 104.035 127.735 105.125 ;
        RECT 121.465 103.515 123.155 104.035 ;
        RECT 126.525 103.495 127.045 104.035 ;
        RECT 15.435 100.945 15.955 101.485 ;
        RECT 14.745 99.855 15.955 100.945 ;
        RECT 16.125 100.945 17.335 101.465 ;
        RECT 16.125 99.855 18.715 100.945 ;
        RECT 20.480 100.290 20.830 101.540 ;
        RECT 18.890 99.855 24.235 100.290 ;
        RECT 24.405 99.855 24.695 101.020 ;
        RECT 25.325 100.945 26.535 101.465 ;
        RECT 25.325 99.855 27.915 100.945 ;
        RECT 28.175 99.855 28.445 100.600 ;
        RECT 29.075 99.860 29.330 100.585 ;
        RECT 29.945 99.860 30.190 100.585 ;
        RECT 30.805 99.860 31.050 100.585 ;
        RECT 31.665 99.860 31.910 100.585 ;
        RECT 32.510 99.860 32.770 100.585 ;
        RECT 33.370 99.860 33.630 100.585 ;
        RECT 34.230 99.860 34.490 100.585 ;
        RECT 35.090 99.860 35.350 100.655 ;
        RECT 29.075 99.855 35.350 99.860 ;
        RECT 35.950 99.855 36.210 100.665 ;
        RECT 36.810 99.855 37.105 100.665 ;
        RECT 37.285 99.855 37.575 101.020 ;
        RECT 38.265 99.855 38.475 100.995 ;
        RECT 39.145 99.855 39.375 100.995 ;
        RECT 40.025 99.855 40.355 100.615 ;
        RECT 41.055 99.855 41.325 100.600 ;
        RECT 41.955 99.860 42.210 100.585 ;
        RECT 42.825 99.860 43.070 100.585 ;
        RECT 43.685 99.860 43.930 100.585 ;
        RECT 44.545 99.860 44.790 100.585 ;
        RECT 45.390 99.860 45.650 100.585 ;
        RECT 46.250 99.860 46.510 100.585 ;
        RECT 47.110 99.860 47.370 100.585 ;
        RECT 47.970 99.860 48.230 100.655 ;
        RECT 41.955 99.855 48.230 99.860 ;
        RECT 48.830 99.855 49.090 100.665 ;
        RECT 49.690 99.855 49.985 100.665 ;
        RECT 50.165 99.855 50.455 101.020 ;
        RECT 51.085 100.945 51.835 101.465 ;
        RECT 51.085 99.855 52.755 100.945 ;
        RECT 53.015 99.855 53.285 100.600 ;
        RECT 53.915 99.860 54.170 100.585 ;
        RECT 54.785 99.860 55.030 100.585 ;
        RECT 55.645 99.860 55.890 100.585 ;
        RECT 56.505 99.860 56.750 100.585 ;
        RECT 57.350 99.860 57.610 100.585 ;
        RECT 58.210 99.860 58.470 100.585 ;
        RECT 59.070 99.860 59.330 100.585 ;
        RECT 59.930 99.860 60.190 100.655 ;
        RECT 53.915 99.855 60.190 99.860 ;
        RECT 60.790 99.855 61.050 100.665 ;
        RECT 61.650 99.855 61.945 100.665 ;
        RECT 63.045 99.855 63.335 101.020 ;
        RECT 73.165 100.945 74.375 101.465 ;
        RECT 63.515 99.855 63.810 100.665 ;
        RECT 64.410 99.855 64.670 100.665 ;
        RECT 65.270 99.860 65.530 100.655 ;
        RECT 66.130 99.860 66.390 100.585 ;
        RECT 66.990 99.860 67.250 100.585 ;
        RECT 67.850 99.860 68.110 100.585 ;
        RECT 68.710 99.860 68.955 100.585 ;
        RECT 69.570 99.860 69.815 100.585 ;
        RECT 70.430 99.860 70.675 100.585 ;
        RECT 71.290 99.860 71.545 100.585 ;
        RECT 65.270 99.855 71.545 99.860 ;
        RECT 72.175 99.855 72.445 100.600 ;
        RECT 73.165 99.855 75.755 100.945 ;
        RECT 75.925 99.855 76.215 101.020 ;
        RECT 86.045 100.945 87.255 101.465 ;
        RECT 76.395 99.855 76.690 100.665 ;
        RECT 77.290 99.855 77.550 100.665 ;
        RECT 78.150 99.860 78.410 100.655 ;
        RECT 79.010 99.860 79.270 100.585 ;
        RECT 79.870 99.860 80.130 100.585 ;
        RECT 80.730 99.860 80.990 100.585 ;
        RECT 81.590 99.860 81.835 100.585 ;
        RECT 82.450 99.860 82.695 100.585 ;
        RECT 83.310 99.860 83.555 100.585 ;
        RECT 84.170 99.860 84.425 100.585 ;
        RECT 78.150 99.855 84.425 99.860 ;
        RECT 85.055 99.855 85.325 100.600 ;
        RECT 86.045 99.855 88.635 100.945 ;
        RECT 88.805 99.855 89.095 101.020 ;
        RECT 98.925 100.945 100.135 101.465 ;
        RECT 89.275 99.855 89.570 100.665 ;
        RECT 90.170 99.855 90.430 100.665 ;
        RECT 91.030 99.860 91.290 100.655 ;
        RECT 91.890 99.860 92.150 100.585 ;
        RECT 92.750 99.860 93.010 100.585 ;
        RECT 93.610 99.860 93.870 100.585 ;
        RECT 94.470 99.860 94.715 100.585 ;
        RECT 95.330 99.860 95.575 100.585 ;
        RECT 96.190 99.860 96.435 100.585 ;
        RECT 97.050 99.860 97.305 100.585 ;
        RECT 91.030 99.855 97.305 99.860 ;
        RECT 97.935 99.855 98.205 100.600 ;
        RECT 98.925 99.855 101.515 100.945 ;
        RECT 101.685 99.855 101.975 101.020 ;
        RECT 111.805 100.945 113.015 101.465 ;
        RECT 102.235 99.855 102.505 100.600 ;
        RECT 103.135 99.860 103.390 100.585 ;
        RECT 104.005 99.860 104.250 100.585 ;
        RECT 104.865 99.860 105.110 100.585 ;
        RECT 105.725 99.860 105.970 100.585 ;
        RECT 106.570 99.860 106.830 100.585 ;
        RECT 107.430 99.860 107.690 100.585 ;
        RECT 108.290 99.860 108.550 100.585 ;
        RECT 109.150 99.860 109.410 100.655 ;
        RECT 103.135 99.855 109.410 99.860 ;
        RECT 110.010 99.855 110.270 100.665 ;
        RECT 110.870 99.855 111.165 100.665 ;
        RECT 111.805 99.855 114.395 100.945 ;
        RECT 114.565 99.855 114.855 101.020 ;
        RECT 124.685 100.945 125.435 101.465 ;
        RECT 126.525 100.945 127.045 101.485 ;
        RECT 115.035 99.855 115.330 100.665 ;
        RECT 115.930 99.855 116.190 100.665 ;
        RECT 116.790 99.860 117.050 100.655 ;
        RECT 117.650 99.860 117.910 100.585 ;
        RECT 118.510 99.860 118.770 100.585 ;
        RECT 119.370 99.860 119.630 100.585 ;
        RECT 120.230 99.860 120.475 100.585 ;
        RECT 121.090 99.860 121.335 100.585 ;
        RECT 121.950 99.860 122.195 100.585 ;
        RECT 122.810 99.860 123.065 100.585 ;
        RECT 116.790 99.855 123.065 99.860 ;
        RECT 123.695 99.855 123.965 100.600 ;
        RECT 124.685 99.855 126.355 100.945 ;
        RECT 126.525 99.855 127.735 100.945 ;
        RECT 14.660 99.685 127.820 99.855 ;
        RECT 19.165 66.070 30.165 66.940 ;
        RECT 19.165 54.930 20.835 66.070 ;
        RECT 21.235 55.300 21.405 65.340 ;
        RECT 27.095 54.930 27.265 66.070 ;
        RECT 29.525 54.930 30.165 66.070 ;
        RECT 19.165 52.860 30.165 54.930 ;
        RECT 19.165 49.370 21.005 52.860 ;
        RECT 22.765 52.780 30.165 52.860 ;
        RECT 21.405 50.095 21.575 52.135 ;
        RECT 22.765 49.370 25.085 52.780 ;
        RECT 19.165 48.650 25.085 49.370 ;
        RECT 24.025 46.290 25.085 48.650 ;
        RECT 26.845 46.290 27.015 52.780 ;
        RECT 28.775 46.290 30.165 52.780 ;
        RECT 30.365 66.080 41.365 66.950 ;
        RECT 30.365 54.940 32.035 66.080 ;
        RECT 32.435 55.310 32.605 65.350 ;
        RECT 38.295 54.940 38.465 66.080 ;
        RECT 40.725 54.940 41.365 66.080 ;
        RECT 30.365 52.870 41.365 54.940 ;
        RECT 30.365 49.380 32.205 52.870 ;
        RECT 33.965 52.790 41.365 52.870 ;
        RECT 32.605 50.105 32.775 52.145 ;
        RECT 33.965 49.380 36.285 52.790 ;
        RECT 30.365 48.660 36.285 49.380 ;
        RECT 24.025 45.800 30.165 46.290 ;
        RECT 35.225 46.300 36.285 48.660 ;
        RECT 38.045 46.300 38.215 52.790 ;
        RECT 39.975 46.300 41.365 52.790 ;
        RECT 41.585 66.050 52.585 66.920 ;
        RECT 41.585 54.910 43.255 66.050 ;
        RECT 43.655 55.280 43.825 65.320 ;
        RECT 49.515 54.910 49.685 66.050 ;
        RECT 51.945 54.910 52.585 66.050 ;
        RECT 41.585 52.840 52.585 54.910 ;
        RECT 41.585 49.350 43.425 52.840 ;
        RECT 45.185 52.760 52.585 52.840 ;
        RECT 43.825 50.075 43.995 52.115 ;
        RECT 45.185 49.350 47.505 52.760 ;
        RECT 41.585 48.630 47.505 49.350 ;
        RECT 35.225 45.810 41.365 46.300 ;
        RECT 46.445 46.270 47.505 48.630 ;
        RECT 49.265 46.270 49.435 52.760 ;
        RECT 51.195 46.270 52.585 52.760 ;
        RECT 52.835 66.030 63.835 66.900 ;
        RECT 52.835 54.890 54.505 66.030 ;
        RECT 54.905 55.260 55.075 65.300 ;
        RECT 60.765 54.890 60.935 66.030 ;
        RECT 63.195 54.890 63.835 66.030 ;
        RECT 52.835 52.820 63.835 54.890 ;
        RECT 52.835 49.330 54.675 52.820 ;
        RECT 56.435 52.740 63.835 52.820 ;
        RECT 55.075 50.055 55.245 52.095 ;
        RECT 56.435 49.330 58.755 52.740 ;
        RECT 52.835 48.610 58.755 49.330 ;
        RECT 46.445 45.780 52.585 46.270 ;
        RECT 57.695 46.250 58.755 48.610 ;
        RECT 60.515 46.250 60.685 52.740 ;
        RECT 62.445 46.250 63.835 52.740 ;
        RECT 64.055 66.020 75.055 66.890 ;
        RECT 64.055 54.880 65.725 66.020 ;
        RECT 66.125 55.250 66.295 65.290 ;
        RECT 71.985 54.880 72.155 66.020 ;
        RECT 74.415 54.880 75.055 66.020 ;
        RECT 64.055 52.810 75.055 54.880 ;
        RECT 64.055 49.320 65.895 52.810 ;
        RECT 67.655 52.730 75.055 52.810 ;
        RECT 66.295 50.045 66.465 52.085 ;
        RECT 67.655 49.320 69.975 52.730 ;
        RECT 64.055 48.600 69.975 49.320 ;
        RECT 57.695 45.760 63.835 46.250 ;
        RECT 68.915 46.240 69.975 48.600 ;
        RECT 71.735 46.240 71.905 52.730 ;
        RECT 73.665 46.240 75.055 52.730 ;
        RECT 75.295 66.010 86.295 66.880 ;
        RECT 75.295 54.870 76.965 66.010 ;
        RECT 77.365 55.240 77.535 65.280 ;
        RECT 83.225 54.870 83.395 66.010 ;
        RECT 85.655 54.870 86.295 66.010 ;
        RECT 75.295 52.800 86.295 54.870 ;
        RECT 75.295 49.310 77.135 52.800 ;
        RECT 78.895 52.720 86.295 52.800 ;
        RECT 77.535 50.035 77.705 52.075 ;
        RECT 78.895 49.310 81.215 52.720 ;
        RECT 75.295 48.590 81.215 49.310 ;
        RECT 68.915 45.750 75.055 46.240 ;
        RECT 80.155 46.230 81.215 48.590 ;
        RECT 82.975 46.230 83.145 52.720 ;
        RECT 84.905 46.230 86.295 52.720 ;
        RECT 86.545 66.020 97.545 66.890 ;
        RECT 131.125 66.880 140.025 66.890 ;
        RECT 86.545 54.880 88.215 66.020 ;
        RECT 88.615 55.250 88.785 65.290 ;
        RECT 94.475 54.880 94.645 66.020 ;
        RECT 96.905 54.880 97.545 66.020 ;
        RECT 86.545 52.810 97.545 54.880 ;
        RECT 86.545 49.320 88.385 52.810 ;
        RECT 90.145 52.730 97.545 52.810 ;
        RECT 88.785 50.045 88.955 52.085 ;
        RECT 90.145 49.320 92.465 52.730 ;
        RECT 86.545 48.600 92.465 49.320 ;
        RECT 80.155 45.740 86.295 46.230 ;
        RECT 91.405 46.240 92.465 48.600 ;
        RECT 94.225 46.240 94.395 52.730 ;
        RECT 96.155 46.240 97.545 52.730 ;
        RECT 97.825 66.010 108.825 66.880 ;
        RECT 97.825 54.870 99.495 66.010 ;
        RECT 99.895 55.240 100.065 65.280 ;
        RECT 105.755 54.870 105.925 66.010 ;
        RECT 108.185 54.870 108.825 66.010 ;
        RECT 97.825 52.800 108.825 54.870 ;
        RECT 97.825 49.310 99.665 52.800 ;
        RECT 101.425 52.720 108.825 52.800 ;
        RECT 100.065 50.035 100.235 52.075 ;
        RECT 101.425 49.310 103.745 52.720 ;
        RECT 97.825 48.590 103.745 49.310 ;
        RECT 91.405 45.750 97.545 46.240 ;
        RECT 102.685 46.230 103.745 48.590 ;
        RECT 105.505 46.230 105.675 52.720 ;
        RECT 107.435 46.230 108.825 52.720 ;
        RECT 109.095 66.010 120.095 66.880 ;
        RECT 109.095 54.870 110.765 66.010 ;
        RECT 111.165 55.240 111.335 65.280 ;
        RECT 117.025 54.870 117.195 66.010 ;
        RECT 119.455 54.870 120.095 66.010 ;
        RECT 109.095 52.800 120.095 54.870 ;
        RECT 109.095 49.310 110.935 52.800 ;
        RECT 112.695 52.720 120.095 52.800 ;
        RECT 111.335 50.035 111.505 52.075 ;
        RECT 112.695 49.310 115.015 52.720 ;
        RECT 109.095 48.590 115.015 49.310 ;
        RECT 102.685 45.740 108.825 46.230 ;
        RECT 113.955 46.230 115.015 48.590 ;
        RECT 116.775 46.230 116.945 52.720 ;
        RECT 118.705 46.230 120.095 52.720 ;
        RECT 120.345 66.010 140.025 66.880 ;
        RECT 120.345 54.870 122.015 66.010 ;
        RECT 122.415 55.240 122.585 65.280 ;
        RECT 128.275 54.870 128.445 66.010 ;
        RECT 130.705 65.980 140.025 66.010 ;
        RECT 130.705 54.870 132.765 65.980 ;
        RECT 133.165 55.210 133.335 65.250 ;
        RECT 120.345 54.840 132.765 54.870 ;
        RECT 139.025 54.840 140.025 65.980 ;
        RECT 120.345 54.720 140.025 54.840 ;
        RECT 120.345 53.550 140.035 54.720 ;
        RECT 120.345 52.800 131.345 53.550 ;
        RECT 120.345 49.310 122.185 52.800 ;
        RECT 123.945 52.720 131.345 52.800 ;
        RECT 122.585 50.035 122.755 52.075 ;
        RECT 123.945 49.310 126.265 52.720 ;
        RECT 120.345 48.590 126.265 49.310 ;
        RECT 113.955 45.740 120.095 46.230 ;
        RECT 125.205 46.230 126.265 48.590 ;
        RECT 128.025 46.230 128.195 52.720 ;
        RECT 129.955 46.230 131.345 52.720 ;
        RECT 125.205 45.740 131.345 46.230 ;
        RECT 18.575 39.120 24.715 39.610 ;
        RECT 18.575 32.630 19.965 39.120 ;
        RECT 21.725 32.630 21.895 39.120 ;
        RECT 23.655 36.760 24.715 39.120 ;
        RECT 29.855 39.120 35.995 39.610 ;
        RECT 23.655 36.040 29.575 36.760 ;
        RECT 23.655 32.630 25.975 36.040 ;
        RECT 27.165 33.275 27.335 35.315 ;
        RECT 18.575 32.550 25.975 32.630 ;
        RECT 27.735 32.550 29.575 36.040 ;
        RECT 18.575 30.480 29.575 32.550 ;
        RECT 18.575 19.340 19.215 30.480 ;
        RECT 21.475 19.340 21.645 30.480 ;
        RECT 27.335 20.070 27.505 30.110 ;
        RECT 27.905 19.340 29.575 30.480 ;
        RECT 18.575 18.470 29.575 19.340 ;
        RECT 29.855 32.630 31.245 39.120 ;
        RECT 33.005 32.630 33.175 39.120 ;
        RECT 34.935 36.760 35.995 39.120 ;
        RECT 41.145 39.100 47.285 39.590 ;
        RECT 34.935 36.040 40.855 36.760 ;
        RECT 34.935 32.630 37.255 36.040 ;
        RECT 38.445 33.275 38.615 35.315 ;
        RECT 29.855 32.550 37.255 32.630 ;
        RECT 39.015 32.550 40.855 36.040 ;
        RECT 29.855 30.480 40.855 32.550 ;
        RECT 29.855 19.340 30.495 30.480 ;
        RECT 32.755 19.340 32.925 30.480 ;
        RECT 38.615 20.070 38.785 30.110 ;
        RECT 39.185 19.340 40.855 30.480 ;
        RECT 29.855 18.470 40.855 19.340 ;
        RECT 41.145 32.610 42.535 39.100 ;
        RECT 44.295 32.610 44.465 39.100 ;
        RECT 46.225 36.740 47.285 39.100 ;
        RECT 52.365 39.100 58.505 39.590 ;
        RECT 46.225 36.020 52.145 36.740 ;
        RECT 46.225 32.610 48.545 36.020 ;
        RECT 49.735 33.255 49.905 35.295 ;
        RECT 41.145 32.530 48.545 32.610 ;
        RECT 50.305 32.530 52.145 36.020 ;
        RECT 41.145 30.460 52.145 32.530 ;
        RECT 41.145 19.320 41.785 30.460 ;
        RECT 44.045 19.320 44.215 30.460 ;
        RECT 49.905 20.050 50.075 30.090 ;
        RECT 50.475 19.320 52.145 30.460 ;
        RECT 41.145 18.450 52.145 19.320 ;
        RECT 52.365 32.610 53.755 39.100 ;
        RECT 55.515 32.610 55.685 39.100 ;
        RECT 57.445 36.740 58.505 39.100 ;
        RECT 63.565 39.100 69.705 39.590 ;
        RECT 57.445 36.020 63.365 36.740 ;
        RECT 57.445 32.610 59.765 36.020 ;
        RECT 60.955 33.255 61.125 35.295 ;
        RECT 52.365 32.530 59.765 32.610 ;
        RECT 61.525 32.530 63.365 36.020 ;
        RECT 52.365 30.460 63.365 32.530 ;
        RECT 52.365 19.320 53.005 30.460 ;
        RECT 55.265 19.320 55.435 30.460 ;
        RECT 61.125 20.050 61.295 30.090 ;
        RECT 61.695 19.320 63.365 30.460 ;
        RECT 52.365 18.450 63.365 19.320 ;
        RECT 63.565 32.610 64.955 39.100 ;
        RECT 66.715 32.610 66.885 39.100 ;
        RECT 68.645 36.740 69.705 39.100 ;
        RECT 74.855 39.090 80.995 39.580 ;
        RECT 68.645 36.020 74.565 36.740 ;
        RECT 68.645 32.610 70.965 36.020 ;
        RECT 72.155 33.255 72.325 35.295 ;
        RECT 63.565 32.530 70.965 32.610 ;
        RECT 72.725 32.530 74.565 36.020 ;
        RECT 63.565 30.460 74.565 32.530 ;
        RECT 63.565 19.320 64.205 30.460 ;
        RECT 66.465 19.320 66.635 30.460 ;
        RECT 72.325 20.050 72.495 30.090 ;
        RECT 72.895 19.320 74.565 30.460 ;
        RECT 63.565 18.450 74.565 19.320 ;
        RECT 74.855 32.600 76.245 39.090 ;
        RECT 78.005 32.600 78.175 39.090 ;
        RECT 79.935 36.730 80.995 39.090 ;
        RECT 86.095 39.110 92.235 39.600 ;
        RECT 79.935 36.010 85.855 36.730 ;
        RECT 79.935 32.600 82.255 36.010 ;
        RECT 83.445 33.245 83.615 35.285 ;
        RECT 74.855 32.520 82.255 32.600 ;
        RECT 84.015 32.520 85.855 36.010 ;
        RECT 74.855 30.450 85.855 32.520 ;
        RECT 74.855 19.310 75.495 30.450 ;
        RECT 77.755 19.310 77.925 30.450 ;
        RECT 83.615 20.040 83.785 30.080 ;
        RECT 84.185 19.310 85.855 30.450 ;
        RECT 74.855 18.440 85.855 19.310 ;
        RECT 86.095 32.620 87.485 39.110 ;
        RECT 89.245 32.620 89.415 39.110 ;
        RECT 91.175 36.750 92.235 39.110 ;
        RECT 97.305 39.130 103.445 39.620 ;
        RECT 91.175 36.030 97.095 36.750 ;
        RECT 91.175 32.620 93.495 36.030 ;
        RECT 94.685 33.265 94.855 35.305 ;
        RECT 86.095 32.540 93.495 32.620 ;
        RECT 95.255 32.540 97.095 36.030 ;
        RECT 86.095 30.470 97.095 32.540 ;
        RECT 86.095 19.330 86.735 30.470 ;
        RECT 88.995 19.330 89.165 30.470 ;
        RECT 94.855 20.060 95.025 30.100 ;
        RECT 95.425 19.330 97.095 30.470 ;
        RECT 86.095 18.460 97.095 19.330 ;
        RECT 97.305 32.640 98.695 39.130 ;
        RECT 100.455 32.640 100.625 39.130 ;
        RECT 102.385 36.770 103.445 39.130 ;
        RECT 108.505 39.170 114.645 39.660 ;
        RECT 102.385 36.050 108.305 36.770 ;
        RECT 102.385 32.640 104.705 36.050 ;
        RECT 105.895 33.285 106.065 35.325 ;
        RECT 97.305 32.560 104.705 32.640 ;
        RECT 106.465 32.560 108.305 36.050 ;
        RECT 97.305 30.490 108.305 32.560 ;
        RECT 97.305 19.350 97.945 30.490 ;
        RECT 100.205 19.350 100.375 30.490 ;
        RECT 106.065 20.080 106.235 30.120 ;
        RECT 106.635 19.350 108.305 30.490 ;
        RECT 97.305 18.480 108.305 19.350 ;
        RECT 108.505 32.680 109.895 39.170 ;
        RECT 111.655 32.680 111.825 39.170 ;
        RECT 113.585 36.810 114.645 39.170 ;
        RECT 119.715 39.190 125.855 39.680 ;
        RECT 113.585 36.090 119.505 36.810 ;
        RECT 113.585 32.680 115.905 36.090 ;
        RECT 117.095 33.325 117.265 35.365 ;
        RECT 108.505 32.600 115.905 32.680 ;
        RECT 117.665 32.600 119.505 36.090 ;
        RECT 108.505 30.530 119.505 32.600 ;
        RECT 108.505 19.390 109.145 30.530 ;
        RECT 111.405 19.390 111.575 30.530 ;
        RECT 117.265 20.120 117.435 30.160 ;
        RECT 117.835 19.390 119.505 30.530 ;
        RECT 108.505 18.520 119.505 19.390 ;
        RECT 119.715 32.700 121.105 39.190 ;
        RECT 122.865 32.700 123.035 39.190 ;
        RECT 124.795 36.830 125.855 39.190 ;
        RECT 124.795 36.110 130.715 36.830 ;
        RECT 124.795 32.700 127.115 36.110 ;
        RECT 128.305 33.345 128.475 35.385 ;
        RECT 119.715 32.620 127.115 32.700 ;
        RECT 128.875 32.620 130.715 36.110 ;
        RECT 119.715 31.140 130.715 32.620 ;
        RECT 119.715 30.550 139.465 31.140 ;
        RECT 119.715 19.410 120.355 30.550 ;
        RECT 122.615 19.410 122.785 30.550 ;
        RECT 129.045 30.520 139.465 30.550 ;
        RECT 128.475 20.140 128.645 30.180 ;
        RECT 129.045 19.410 132.075 30.520 ;
        RECT 132.475 20.110 132.645 30.150 ;
        RECT 119.715 19.380 132.075 19.410 ;
        RECT 138.335 19.380 139.465 30.520 ;
        RECT 119.715 18.540 139.465 19.380 ;
        RECT 131.925 18.520 139.465 18.540 ;
      LAYER met1 ;
        RECT 14.660 208.330 127.820 208.810 ;
        RECT 14.660 202.890 127.820 203.370 ;
        RECT 14.660 197.450 127.820 197.930 ;
        RECT 14.660 192.010 127.820 192.490 ;
        RECT 14.660 186.570 127.820 187.050 ;
        RECT 14.660 181.130 127.820 181.610 ;
        RECT 14.660 175.690 127.820 176.170 ;
        RECT 14.660 170.250 127.820 170.730 ;
        RECT 14.660 164.810 127.820 165.290 ;
        RECT 14.660 159.370 127.820 159.850 ;
        RECT 14.660 153.930 127.820 154.410 ;
        RECT 14.660 148.490 127.820 148.970 ;
        RECT 14.660 143.050 127.820 143.530 ;
        RECT 14.660 137.610 127.820 138.090 ;
        RECT 14.660 132.170 127.820 132.650 ;
        RECT 14.660 126.730 127.820 127.210 ;
        RECT 14.660 121.290 127.820 121.770 ;
        RECT 14.660 115.850 127.820 116.330 ;
        RECT 14.660 110.410 127.820 110.890 ;
        RECT 14.660 104.970 127.820 105.450 ;
        RECT 14.660 99.530 127.820 100.010 ;
        RECT 137.920 77.810 143.450 77.960 ;
        RECT 137.190 76.610 143.450 77.810 ;
        RECT 137.920 75.460 143.450 76.610 ;
        RECT 29.635 71.170 43.285 71.180 ;
        RECT 15.510 71.155 17.040 71.160 ;
        RECT 18.435 71.155 43.285 71.170 ;
        RECT 12.285 71.150 43.285 71.155 ;
        RECT 12.285 71.130 54.505 71.150 ;
        RECT 141.810 71.140 143.230 75.460 ;
        RECT 12.285 71.120 65.755 71.130 ;
        RECT 12.285 71.110 76.975 71.120 ;
        RECT 85.815 71.110 99.465 71.120 ;
        RECT 140.220 71.110 143.240 71.140 ;
        RECT 12.285 70.030 143.240 71.110 ;
        RECT 12.285 70.020 32.085 70.030 ;
        RECT 12.285 70.005 19.375 70.020 ;
        RECT 12.320 15.450 13.470 70.005 ;
        RECT 15.510 68.660 17.040 70.005 ;
        RECT 40.855 70.000 143.240 70.030 ;
        RECT 52.105 69.980 143.240 70.000 ;
        RECT 63.325 69.970 143.240 69.980 ;
        RECT 74.565 69.960 88.215 69.970 ;
        RECT 97.095 69.960 143.240 69.970 ;
        RECT 140.220 69.910 143.240 69.960 ;
        RECT 21.205 65.140 21.435 65.320 ;
        RECT 32.405 65.150 32.635 65.330 ;
        RECT 21.125 55.220 21.485 65.140 ;
        RECT 32.325 55.230 32.685 65.150 ;
        RECT 43.625 65.120 43.855 65.300 ;
        RECT 43.545 55.200 43.905 65.120 ;
        RECT 54.875 65.100 55.105 65.280 ;
        RECT 54.795 55.180 55.155 65.100 ;
        RECT 66.095 65.090 66.325 65.270 ;
        RECT 66.015 55.170 66.375 65.090 ;
        RECT 77.335 65.080 77.565 65.260 ;
        RECT 88.585 65.090 88.815 65.270 ;
        RECT 77.255 55.160 77.615 65.080 ;
        RECT 88.505 55.170 88.865 65.090 ;
        RECT 99.865 65.080 100.095 65.260 ;
        RECT 111.135 65.080 111.365 65.260 ;
        RECT 122.385 65.080 122.615 65.260 ;
        RECT 133.135 65.130 133.365 65.230 ;
        RECT 99.785 55.160 100.145 65.080 ;
        RECT 111.055 55.160 111.415 65.080 ;
        RECT 122.305 55.160 122.665 65.080 ;
        RECT 133.005 55.240 133.405 65.130 ;
        RECT 133.135 55.230 133.365 55.240 ;
        RECT 20.815 54.230 25.555 54.530 ;
        RECT 32.015 54.240 36.755 54.540 ;
        RECT 43.235 54.210 47.975 54.510 ;
        RECT 54.485 54.190 59.225 54.490 ;
        RECT 65.705 54.180 70.445 54.480 ;
        RECT 76.945 54.170 81.685 54.470 ;
        RECT 88.195 54.180 92.935 54.480 ;
        RECT 99.475 54.170 104.215 54.470 ;
        RECT 110.745 54.170 115.485 54.470 ;
        RECT 121.995 54.170 126.735 54.470 ;
        RECT 21.375 52.010 21.605 52.115 ;
        RECT 32.575 52.020 32.805 52.125 ;
        RECT 21.245 50.290 21.615 52.010 ;
        RECT 32.445 50.300 32.815 52.020 ;
        RECT 43.795 51.990 44.025 52.095 ;
        RECT 21.375 50.115 21.605 50.290 ;
        RECT 32.575 50.125 32.805 50.300 ;
        RECT 43.665 50.270 44.035 51.990 ;
        RECT 55.045 51.970 55.275 52.075 ;
        RECT 43.795 50.095 44.025 50.270 ;
        RECT 54.915 50.250 55.285 51.970 ;
        RECT 66.265 51.960 66.495 52.065 ;
        RECT 55.045 50.075 55.275 50.250 ;
        RECT 66.135 50.240 66.505 51.960 ;
        RECT 77.505 51.950 77.735 52.055 ;
        RECT 88.755 51.960 88.985 52.065 ;
        RECT 66.265 50.065 66.495 50.240 ;
        RECT 77.375 50.230 77.745 51.950 ;
        RECT 88.625 50.240 88.995 51.960 ;
        RECT 100.035 51.950 100.265 52.055 ;
        RECT 111.305 51.950 111.535 52.055 ;
        RECT 122.555 51.950 122.785 52.055 ;
        RECT 77.505 50.055 77.735 50.230 ;
        RECT 88.755 50.065 88.985 50.240 ;
        RECT 99.905 50.230 100.275 51.950 ;
        RECT 111.175 50.230 111.545 51.950 ;
        RECT 122.425 50.230 122.795 51.950 ;
        RECT 100.035 50.055 100.265 50.230 ;
        RECT 111.305 50.055 111.535 50.230 ;
        RECT 122.555 50.055 122.785 50.230 ;
        RECT 27.135 35.120 27.365 35.295 ;
        RECT 38.415 35.120 38.645 35.295 ;
        RECT 27.125 33.400 27.495 35.120 ;
        RECT 38.405 33.400 38.775 35.120 ;
        RECT 49.705 35.100 49.935 35.275 ;
        RECT 60.925 35.100 61.155 35.275 ;
        RECT 72.125 35.100 72.355 35.275 ;
        RECT 27.135 33.295 27.365 33.400 ;
        RECT 38.415 33.295 38.645 33.400 ;
        RECT 49.695 33.380 50.065 35.100 ;
        RECT 60.915 33.380 61.285 35.100 ;
        RECT 72.115 33.380 72.485 35.100 ;
        RECT 83.415 35.090 83.645 35.265 ;
        RECT 94.655 35.110 94.885 35.285 ;
        RECT 105.865 35.130 106.095 35.305 ;
        RECT 117.065 35.170 117.295 35.345 ;
        RECT 128.275 35.190 128.505 35.365 ;
        RECT 49.705 33.275 49.935 33.380 ;
        RECT 60.925 33.275 61.155 33.380 ;
        RECT 72.125 33.275 72.355 33.380 ;
        RECT 83.405 33.370 83.775 35.090 ;
        RECT 94.645 33.390 95.015 35.110 ;
        RECT 105.855 33.410 106.225 35.130 ;
        RECT 117.055 33.450 117.425 35.170 ;
        RECT 128.265 33.470 128.635 35.190 ;
        RECT 83.415 33.265 83.645 33.370 ;
        RECT 94.655 33.285 94.885 33.390 ;
        RECT 105.865 33.305 106.095 33.410 ;
        RECT 117.065 33.345 117.295 33.450 ;
        RECT 128.275 33.365 128.505 33.470 ;
        RECT 23.185 30.880 27.925 31.180 ;
        RECT 34.465 30.880 39.205 31.180 ;
        RECT 45.755 30.860 50.495 31.160 ;
        RECT 56.975 30.860 61.715 31.160 ;
        RECT 68.175 30.860 72.915 31.160 ;
        RECT 79.465 30.850 84.205 31.150 ;
        RECT 90.705 30.870 95.445 31.170 ;
        RECT 101.915 30.890 106.655 31.190 ;
        RECT 113.115 30.930 117.855 31.230 ;
        RECT 124.325 30.950 129.065 31.250 ;
        RECT 27.255 20.270 27.615 30.190 ;
        RECT 38.535 20.270 38.895 30.190 ;
        RECT 27.305 20.090 27.535 20.270 ;
        RECT 38.585 20.090 38.815 20.270 ;
        RECT 49.825 20.250 50.185 30.170 ;
        RECT 61.045 20.250 61.405 30.170 ;
        RECT 72.245 20.250 72.605 30.170 ;
        RECT 49.875 20.070 50.105 20.250 ;
        RECT 61.095 20.070 61.325 20.250 ;
        RECT 72.295 20.070 72.525 20.250 ;
        RECT 83.535 20.240 83.895 30.160 ;
        RECT 94.775 20.260 95.135 30.180 ;
        RECT 105.985 20.280 106.345 30.200 ;
        RECT 117.185 20.320 117.545 30.240 ;
        RECT 128.395 20.340 128.755 30.260 ;
        RECT 83.585 20.060 83.815 20.240 ;
        RECT 94.825 20.080 95.055 20.260 ;
        RECT 106.035 20.100 106.265 20.280 ;
        RECT 117.235 20.140 117.465 20.320 ;
        RECT 128.445 20.160 128.675 20.340 ;
        RECT 132.345 20.170 132.755 30.180 ;
        RECT 132.445 20.130 132.675 20.170 ;
        RECT 131.215 15.460 132.585 15.470 ;
        RECT 12.290 15.390 17.625 15.450 ;
        RECT 117.795 15.440 132.785 15.460 ;
        RECT 106.585 15.400 132.785 15.440 ;
        RECT 12.290 15.370 41.585 15.390 ;
        RECT 95.385 15.380 132.785 15.400 ;
        RECT 12.290 15.360 75.295 15.370 ;
        RECT 84.175 15.360 132.785 15.380 ;
        RECT 12.290 14.320 132.785 15.360 ;
        RECT 12.290 14.310 131.445 14.320 ;
        RECT 12.290 14.300 120.235 14.310 ;
        RECT 12.320 14.280 13.470 14.300 ;
        RECT 16.655 14.290 120.235 14.300 ;
        RECT 16.655 14.250 109.035 14.290 ;
        RECT 16.655 14.240 97.825 14.250 ;
        RECT 39.225 14.230 97.825 14.240 ;
        RECT 39.225 14.220 86.585 14.230 ;
        RECT 72.935 14.210 86.585 14.220 ;
      LAYER met2 ;
        RECT 31.880 208.385 33.760 208.755 ;
        RECT 61.880 208.385 63.760 208.755 ;
        RECT 91.880 208.385 93.760 208.755 ;
        RECT 121.880 208.385 123.760 208.755 ;
        RECT 31.880 202.945 33.760 203.315 ;
        RECT 61.880 202.945 63.760 203.315 ;
        RECT 91.880 202.945 93.760 203.315 ;
        RECT 121.880 202.945 123.760 203.315 ;
        RECT 31.880 197.505 33.760 197.875 ;
        RECT 61.880 197.505 63.760 197.875 ;
        RECT 91.880 197.505 93.760 197.875 ;
        RECT 121.880 197.505 123.760 197.875 ;
        RECT 31.880 192.065 33.760 192.435 ;
        RECT 61.880 192.065 63.760 192.435 ;
        RECT 91.880 192.065 93.760 192.435 ;
        RECT 121.880 192.065 123.760 192.435 ;
        RECT 31.880 186.625 33.760 186.995 ;
        RECT 61.880 186.625 63.760 186.995 ;
        RECT 91.880 186.625 93.760 186.995 ;
        RECT 121.880 186.625 123.760 186.995 ;
        RECT 31.880 181.185 33.760 181.555 ;
        RECT 61.880 181.185 63.760 181.555 ;
        RECT 91.880 181.185 93.760 181.555 ;
        RECT 121.880 181.185 123.760 181.555 ;
        RECT 31.880 175.745 33.760 176.115 ;
        RECT 61.880 175.745 63.760 176.115 ;
        RECT 91.880 175.745 93.760 176.115 ;
        RECT 121.880 175.745 123.760 176.115 ;
        RECT 31.880 170.305 33.760 170.675 ;
        RECT 61.880 170.305 63.760 170.675 ;
        RECT 91.880 170.305 93.760 170.675 ;
        RECT 121.880 170.305 123.760 170.675 ;
        RECT 31.880 164.865 33.760 165.235 ;
        RECT 61.880 164.865 63.760 165.235 ;
        RECT 91.880 164.865 93.760 165.235 ;
        RECT 121.880 164.865 123.760 165.235 ;
        RECT 31.880 159.425 33.760 159.795 ;
        RECT 61.880 159.425 63.760 159.795 ;
        RECT 91.880 159.425 93.760 159.795 ;
        RECT 121.880 159.425 123.760 159.795 ;
        RECT 31.880 153.985 33.760 154.355 ;
        RECT 61.880 153.985 63.760 154.355 ;
        RECT 91.880 153.985 93.760 154.355 ;
        RECT 121.880 153.985 123.760 154.355 ;
        RECT 31.880 148.545 33.760 148.915 ;
        RECT 61.880 148.545 63.760 148.915 ;
        RECT 91.880 148.545 93.760 148.915 ;
        RECT 121.880 148.545 123.760 148.915 ;
        RECT 31.880 143.105 33.760 143.475 ;
        RECT 61.880 143.105 63.760 143.475 ;
        RECT 91.880 143.105 93.760 143.475 ;
        RECT 121.880 143.105 123.760 143.475 ;
        RECT 31.880 137.665 33.760 138.035 ;
        RECT 61.880 137.665 63.760 138.035 ;
        RECT 91.880 137.665 93.760 138.035 ;
        RECT 121.880 137.665 123.760 138.035 ;
        RECT 31.880 132.225 33.760 132.595 ;
        RECT 61.880 132.225 63.760 132.595 ;
        RECT 91.880 132.225 93.760 132.595 ;
        RECT 121.880 132.225 123.760 132.595 ;
        RECT 31.880 126.785 33.760 127.155 ;
        RECT 61.880 126.785 63.760 127.155 ;
        RECT 91.880 126.785 93.760 127.155 ;
        RECT 121.880 126.785 123.760 127.155 ;
        RECT 31.880 121.345 33.760 121.715 ;
        RECT 61.880 121.345 63.760 121.715 ;
        RECT 91.880 121.345 93.760 121.715 ;
        RECT 121.880 121.345 123.760 121.715 ;
        RECT 31.880 115.905 33.760 116.275 ;
        RECT 61.880 115.905 63.760 116.275 ;
        RECT 91.880 115.905 93.760 116.275 ;
        RECT 121.880 115.905 123.760 116.275 ;
        RECT 31.880 110.465 33.760 110.835 ;
        RECT 61.880 110.465 63.760 110.835 ;
        RECT 91.880 110.465 93.760 110.835 ;
        RECT 121.880 110.465 123.760 110.835 ;
        RECT 31.880 105.025 33.760 105.395 ;
        RECT 61.880 105.025 63.760 105.395 ;
        RECT 91.880 105.025 93.760 105.395 ;
        RECT 121.880 105.025 123.760 105.395 ;
        RECT 31.880 99.585 33.760 99.955 ;
        RECT 61.880 99.585 63.760 99.955 ;
        RECT 91.880 99.585 93.760 99.955 ;
        RECT 121.880 99.585 123.760 99.955 ;
        RECT 137.240 76.560 139.870 77.860 ;
        RECT 15.560 68.610 16.990 71.210 ;
        RECT 132.925 70.810 133.225 70.900 ;
        RECT 20.955 70.010 21.845 70.740 ;
        RECT 32.155 70.020 33.045 70.750 ;
        RECT 21.055 65.190 21.315 70.010 ;
        RECT 32.255 65.200 32.515 70.020 ;
        RECT 43.375 69.990 44.265 70.720 ;
        RECT 21.055 63.640 21.435 65.190 ;
        RECT 32.255 63.650 32.635 65.200 ;
        RECT 21.175 55.800 21.435 63.640 ;
        RECT 32.375 55.810 32.635 63.650 ;
        RECT 43.475 65.170 43.735 69.990 ;
        RECT 54.625 69.970 55.515 70.700 ;
        RECT 43.475 63.620 43.855 65.170 ;
        RECT 21.085 55.290 21.445 55.800 ;
        RECT 32.285 55.300 32.645 55.810 ;
        RECT 43.595 55.780 43.855 63.620 ;
        RECT 54.725 65.150 54.985 69.970 ;
        RECT 65.845 69.960 66.735 70.690 ;
        RECT 54.725 63.600 55.105 65.150 ;
        RECT 21.065 54.860 21.445 55.290 ;
        RECT 32.265 54.870 32.645 55.300 ;
        RECT 43.505 55.270 43.865 55.780 ;
        RECT 54.845 55.760 55.105 63.600 ;
        RECT 65.945 65.140 66.205 69.960 ;
        RECT 77.085 69.950 77.975 70.680 ;
        RECT 88.335 69.960 89.225 70.690 ;
        RECT 65.945 63.590 66.325 65.140 ;
        RECT 21.065 54.580 21.315 54.860 ;
        RECT 32.265 54.590 32.515 54.870 ;
        RECT 43.485 54.840 43.865 55.270 ;
        RECT 54.755 55.250 55.115 55.760 ;
        RECT 66.065 55.750 66.325 63.590 ;
        RECT 77.185 65.130 77.445 69.950 ;
        RECT 88.435 65.140 88.695 69.960 ;
        RECT 99.615 69.950 100.505 70.680 ;
        RECT 110.885 69.950 111.775 70.680 ;
        RECT 122.135 69.950 123.025 70.680 ;
        RECT 132.615 70.040 134.265 70.810 ;
        RECT 77.185 63.580 77.565 65.130 ;
        RECT 88.435 63.590 88.815 65.140 ;
        RECT 20.865 54.180 25.505 54.580 ;
        RECT 32.065 54.190 36.705 54.590 ;
        RECT 43.485 54.560 43.735 54.840 ;
        RECT 54.735 54.820 55.115 55.250 ;
        RECT 65.975 55.240 66.335 55.750 ;
        RECT 77.305 55.740 77.565 63.580 ;
        RECT 88.555 55.750 88.815 63.590 ;
        RECT 99.715 65.130 99.975 69.950 ;
        RECT 110.985 65.130 111.245 69.950 ;
        RECT 122.235 65.130 122.495 69.950 ;
        RECT 132.925 65.180 133.225 70.040 ;
        RECT 99.715 63.580 100.095 65.130 ;
        RECT 110.985 63.580 111.365 65.130 ;
        RECT 122.235 63.580 122.615 65.130 ;
        RECT 21.065 52.060 21.315 54.180 ;
        RECT 32.265 52.070 32.515 54.190 ;
        RECT 43.285 54.160 47.925 54.560 ;
        RECT 54.735 54.540 54.985 54.820 ;
        RECT 65.955 54.810 66.335 55.240 ;
        RECT 77.215 55.230 77.575 55.740 ;
        RECT 88.465 55.240 88.825 55.750 ;
        RECT 99.835 55.740 100.095 63.580 ;
        RECT 111.105 55.740 111.365 63.580 ;
        RECT 122.355 55.740 122.615 63.580 ;
        RECT 132.925 61.010 133.355 65.180 ;
        RECT 21.065 51.970 21.565 52.060 ;
        RECT 32.265 51.980 32.765 52.070 ;
        RECT 21.055 51.240 21.565 51.970 ;
        RECT 32.255 51.250 32.765 51.980 ;
        RECT 43.485 52.040 43.735 54.160 ;
        RECT 54.535 54.140 59.175 54.540 ;
        RECT 65.955 54.530 66.205 54.810 ;
        RECT 77.195 54.800 77.575 55.230 ;
        RECT 88.445 54.810 88.825 55.240 ;
        RECT 99.745 55.230 100.105 55.740 ;
        RECT 111.015 55.230 111.375 55.740 ;
        RECT 122.265 55.230 122.625 55.740 ;
        RECT 43.485 51.950 43.985 52.040 ;
        RECT 21.295 50.240 21.565 51.240 ;
        RECT 32.495 50.250 32.765 51.250 ;
        RECT 43.475 51.220 43.985 51.950 ;
        RECT 54.735 52.020 54.985 54.140 ;
        RECT 65.755 54.130 70.395 54.530 ;
        RECT 77.195 54.520 77.445 54.800 ;
        RECT 88.445 54.530 88.695 54.810 ;
        RECT 99.725 54.800 100.105 55.230 ;
        RECT 110.995 54.800 111.375 55.230 ;
        RECT 122.245 54.800 122.625 55.230 ;
        RECT 133.055 55.190 133.355 61.010 ;
        RECT 54.735 51.930 55.235 52.020 ;
        RECT 43.715 50.220 43.985 51.220 ;
        RECT 54.725 51.200 55.235 51.930 ;
        RECT 65.955 52.010 66.205 54.130 ;
        RECT 76.995 54.120 81.635 54.520 ;
        RECT 88.245 54.130 92.885 54.530 ;
        RECT 99.725 54.520 99.975 54.800 ;
        RECT 110.995 54.520 111.245 54.800 ;
        RECT 122.245 54.520 122.495 54.800 ;
        RECT 65.955 51.920 66.455 52.010 ;
        RECT 54.965 50.200 55.235 51.200 ;
        RECT 65.945 51.190 66.455 51.920 ;
        RECT 77.195 52.000 77.445 54.120 ;
        RECT 88.445 52.010 88.695 54.130 ;
        RECT 99.525 54.120 104.165 54.520 ;
        RECT 110.795 54.120 115.435 54.520 ;
        RECT 122.045 54.120 126.685 54.520 ;
        RECT 77.195 51.910 77.695 52.000 ;
        RECT 88.445 51.920 88.945 52.010 ;
        RECT 66.185 50.190 66.455 51.190 ;
        RECT 77.185 51.180 77.695 51.910 ;
        RECT 88.435 51.190 88.945 51.920 ;
        RECT 99.725 52.000 99.975 54.120 ;
        RECT 110.995 52.000 111.245 54.120 ;
        RECT 122.245 52.000 122.495 54.120 ;
        RECT 99.725 51.910 100.225 52.000 ;
        RECT 110.995 51.910 111.495 52.000 ;
        RECT 122.245 51.910 122.745 52.000 ;
        RECT 77.425 50.180 77.695 51.180 ;
        RECT 88.675 50.190 88.945 51.190 ;
        RECT 99.715 51.180 100.225 51.910 ;
        RECT 110.985 51.180 111.495 51.910 ;
        RECT 122.235 51.180 122.745 51.910 ;
        RECT 99.955 50.180 100.225 51.180 ;
        RECT 111.225 50.180 111.495 51.180 ;
        RECT 122.475 50.180 122.745 51.180 ;
        RECT 27.175 34.170 27.445 35.170 ;
        RECT 38.455 34.170 38.725 35.170 ;
        RECT 27.175 33.440 27.685 34.170 ;
        RECT 38.455 33.440 38.965 34.170 ;
        RECT 49.745 34.150 50.015 35.150 ;
        RECT 60.965 34.150 61.235 35.150 ;
        RECT 72.165 34.150 72.435 35.150 ;
        RECT 27.175 33.350 27.675 33.440 ;
        RECT 38.455 33.350 38.955 33.440 ;
        RECT 27.425 31.230 27.675 33.350 ;
        RECT 38.705 31.230 38.955 33.350 ;
        RECT 49.745 33.420 50.255 34.150 ;
        RECT 60.965 33.420 61.475 34.150 ;
        RECT 72.165 33.420 72.675 34.150 ;
        RECT 83.455 34.140 83.725 35.140 ;
        RECT 94.695 34.160 94.965 35.160 ;
        RECT 105.905 34.180 106.175 35.180 ;
        RECT 117.105 34.220 117.375 35.220 ;
        RECT 128.315 34.240 128.585 35.240 ;
        RECT 49.745 33.330 50.245 33.420 ;
        RECT 60.965 33.330 61.465 33.420 ;
        RECT 72.165 33.330 72.665 33.420 ;
        RECT 23.235 30.830 27.875 31.230 ;
        RECT 34.515 30.830 39.155 31.230 ;
        RECT 49.995 31.210 50.245 33.330 ;
        RECT 61.215 31.210 61.465 33.330 ;
        RECT 72.415 31.210 72.665 33.330 ;
        RECT 83.455 33.410 83.965 34.140 ;
        RECT 94.695 33.430 95.205 34.160 ;
        RECT 105.905 33.450 106.415 34.180 ;
        RECT 117.105 33.490 117.615 34.220 ;
        RECT 128.315 33.510 128.825 34.240 ;
        RECT 83.455 33.320 83.955 33.410 ;
        RECT 94.695 33.340 95.195 33.430 ;
        RECT 105.905 33.360 106.405 33.450 ;
        RECT 117.105 33.400 117.605 33.490 ;
        RECT 128.315 33.420 128.815 33.510 ;
        RECT 27.425 30.550 27.675 30.830 ;
        RECT 38.705 30.550 38.955 30.830 ;
        RECT 45.805 30.810 50.445 31.210 ;
        RECT 57.025 30.810 61.665 31.210 ;
        RECT 68.225 30.810 72.865 31.210 ;
        RECT 83.705 31.200 83.955 33.320 ;
        RECT 94.945 31.220 95.195 33.340 ;
        RECT 106.155 31.240 106.405 33.360 ;
        RECT 117.355 31.280 117.605 33.400 ;
        RECT 128.565 31.300 128.815 33.420 ;
        RECT 27.295 30.120 27.675 30.550 ;
        RECT 38.575 30.120 38.955 30.550 ;
        RECT 49.995 30.530 50.245 30.810 ;
        RECT 61.215 30.530 61.465 30.810 ;
        RECT 72.415 30.530 72.665 30.810 ;
        RECT 79.515 30.800 84.155 31.200 ;
        RECT 90.755 30.820 95.395 31.220 ;
        RECT 101.965 30.840 106.605 31.240 ;
        RECT 113.165 30.880 117.805 31.280 ;
        RECT 124.375 30.900 129.015 31.300 ;
        RECT 27.295 29.610 27.655 30.120 ;
        RECT 38.575 29.610 38.935 30.120 ;
        RECT 49.865 30.100 50.245 30.530 ;
        RECT 61.085 30.100 61.465 30.530 ;
        RECT 72.285 30.100 72.665 30.530 ;
        RECT 83.705 30.520 83.955 30.800 ;
        RECT 94.945 30.540 95.195 30.820 ;
        RECT 106.155 30.560 106.405 30.840 ;
        RECT 117.355 30.600 117.605 30.880 ;
        RECT 128.565 30.620 128.815 30.900 ;
        RECT 27.305 21.770 27.565 29.610 ;
        RECT 38.585 21.770 38.845 29.610 ;
        RECT 49.865 29.590 50.225 30.100 ;
        RECT 61.085 29.590 61.445 30.100 ;
        RECT 72.285 29.590 72.645 30.100 ;
        RECT 83.575 30.090 83.955 30.520 ;
        RECT 94.815 30.110 95.195 30.540 ;
        RECT 106.025 30.130 106.405 30.560 ;
        RECT 117.225 30.170 117.605 30.600 ;
        RECT 128.435 30.190 128.815 30.620 ;
        RECT 27.305 20.220 27.685 21.770 ;
        RECT 38.585 20.220 38.965 21.770 ;
        RECT 27.425 15.400 27.685 20.220 ;
        RECT 38.705 15.400 38.965 20.220 ;
        RECT 49.875 21.750 50.135 29.590 ;
        RECT 61.095 21.750 61.355 29.590 ;
        RECT 72.295 21.750 72.555 29.590 ;
        RECT 83.575 29.580 83.935 30.090 ;
        RECT 94.815 29.600 95.175 30.110 ;
        RECT 106.025 29.620 106.385 30.130 ;
        RECT 117.225 29.660 117.585 30.170 ;
        RECT 128.435 29.680 128.795 30.190 ;
        RECT 49.875 20.200 50.255 21.750 ;
        RECT 61.095 20.200 61.475 21.750 ;
        RECT 72.295 20.200 72.675 21.750 ;
        RECT 26.895 14.670 27.785 15.400 ;
        RECT 38.175 14.670 39.065 15.400 ;
        RECT 49.995 15.380 50.255 20.200 ;
        RECT 61.215 15.380 61.475 20.200 ;
        RECT 72.415 15.380 72.675 20.200 ;
        RECT 83.585 21.740 83.845 29.580 ;
        RECT 94.825 21.760 95.085 29.600 ;
        RECT 106.035 21.780 106.295 29.620 ;
        RECT 117.235 21.820 117.495 29.660 ;
        RECT 128.445 21.840 128.705 29.680 ;
        RECT 132.395 24.340 132.705 30.230 ;
        RECT 83.585 20.190 83.965 21.740 ;
        RECT 94.825 20.210 95.205 21.760 ;
        RECT 106.035 20.230 106.415 21.780 ;
        RECT 117.235 20.270 117.615 21.820 ;
        RECT 128.445 20.290 128.825 21.840 ;
        RECT 49.465 14.650 50.355 15.380 ;
        RECT 60.685 14.650 61.575 15.380 ;
        RECT 71.885 14.650 72.775 15.380 ;
        RECT 83.705 15.370 83.965 20.190 ;
        RECT 94.945 15.390 95.205 20.210 ;
        RECT 106.155 15.410 106.415 20.230 ;
        RECT 117.355 15.450 117.615 20.270 ;
        RECT 128.565 15.470 128.825 20.290 ;
        RECT 132.195 20.120 132.705 24.340 ;
        RECT 132.195 15.510 132.505 20.120 ;
        RECT 83.175 14.640 84.065 15.370 ;
        RECT 94.415 14.660 95.305 15.390 ;
        RECT 105.625 14.680 106.515 15.410 ;
        RECT 116.825 14.720 117.715 15.450 ;
        RECT 128.035 14.740 128.925 15.470 ;
        RECT 131.975 14.270 132.735 15.510 ;
      LAYER met3 ;
        RECT 31.830 208.405 33.810 208.735 ;
        RECT 61.830 208.405 63.810 208.735 ;
        RECT 91.830 208.405 93.810 208.735 ;
        RECT 121.830 208.405 123.810 208.735 ;
        RECT 31.830 202.965 33.810 203.295 ;
        RECT 61.830 202.965 63.810 203.295 ;
        RECT 91.830 202.965 93.810 203.295 ;
        RECT 121.830 202.965 123.810 203.295 ;
        RECT 31.830 197.525 33.810 197.855 ;
        RECT 61.830 197.525 63.810 197.855 ;
        RECT 91.830 197.525 93.810 197.855 ;
        RECT 121.830 197.525 123.810 197.855 ;
        RECT 31.830 192.085 33.810 192.415 ;
        RECT 61.830 192.085 63.810 192.415 ;
        RECT 91.830 192.085 93.810 192.415 ;
        RECT 121.830 192.085 123.810 192.415 ;
        RECT 31.830 186.645 33.810 186.975 ;
        RECT 61.830 186.645 63.810 186.975 ;
        RECT 91.830 186.645 93.810 186.975 ;
        RECT 121.830 186.645 123.810 186.975 ;
        RECT 31.830 181.205 33.810 181.535 ;
        RECT 61.830 181.205 63.810 181.535 ;
        RECT 91.830 181.205 93.810 181.535 ;
        RECT 121.830 181.205 123.810 181.535 ;
        RECT 31.830 175.765 33.810 176.095 ;
        RECT 61.830 175.765 63.810 176.095 ;
        RECT 91.830 175.765 93.810 176.095 ;
        RECT 121.830 175.765 123.810 176.095 ;
        RECT 31.830 170.325 33.810 170.655 ;
        RECT 61.830 170.325 63.810 170.655 ;
        RECT 91.830 170.325 93.810 170.655 ;
        RECT 121.830 170.325 123.810 170.655 ;
        RECT 31.830 164.885 33.810 165.215 ;
        RECT 61.830 164.885 63.810 165.215 ;
        RECT 91.830 164.885 93.810 165.215 ;
        RECT 121.830 164.885 123.810 165.215 ;
        RECT 31.830 159.445 33.810 159.775 ;
        RECT 61.830 159.445 63.810 159.775 ;
        RECT 91.830 159.445 93.810 159.775 ;
        RECT 121.830 159.445 123.810 159.775 ;
        RECT 31.830 154.005 33.810 154.335 ;
        RECT 61.830 154.005 63.810 154.335 ;
        RECT 91.830 154.005 93.810 154.335 ;
        RECT 121.830 154.005 123.810 154.335 ;
        RECT 31.830 148.565 33.810 148.895 ;
        RECT 61.830 148.565 63.810 148.895 ;
        RECT 91.830 148.565 93.810 148.895 ;
        RECT 121.830 148.565 123.810 148.895 ;
        RECT 31.830 143.125 33.810 143.455 ;
        RECT 61.830 143.125 63.810 143.455 ;
        RECT 91.830 143.125 93.810 143.455 ;
        RECT 121.830 143.125 123.810 143.455 ;
        RECT 31.830 137.685 33.810 138.015 ;
        RECT 61.830 137.685 63.810 138.015 ;
        RECT 91.830 137.685 93.810 138.015 ;
        RECT 121.830 137.685 123.810 138.015 ;
        RECT 31.830 132.245 33.810 132.575 ;
        RECT 61.830 132.245 63.810 132.575 ;
        RECT 91.830 132.245 93.810 132.575 ;
        RECT 121.830 132.245 123.810 132.575 ;
        RECT 31.830 126.805 33.810 127.135 ;
        RECT 61.830 126.805 63.810 127.135 ;
        RECT 91.830 126.805 93.810 127.135 ;
        RECT 121.830 126.805 123.810 127.135 ;
        RECT 31.830 121.365 33.810 121.695 ;
        RECT 61.830 121.365 63.810 121.695 ;
        RECT 91.830 121.365 93.810 121.695 ;
        RECT 121.830 121.365 123.810 121.695 ;
        RECT 31.830 115.925 33.810 116.255 ;
        RECT 61.830 115.925 63.810 116.255 ;
        RECT 91.830 115.925 93.810 116.255 ;
        RECT 121.830 115.925 123.810 116.255 ;
        RECT 31.830 110.485 33.810 110.815 ;
        RECT 61.830 110.485 63.810 110.815 ;
        RECT 91.830 110.485 93.810 110.815 ;
        RECT 121.830 110.485 123.810 110.815 ;
        RECT 31.830 105.045 33.810 105.375 ;
        RECT 61.830 105.045 63.810 105.375 ;
        RECT 91.830 105.045 93.810 105.375 ;
        RECT 121.830 105.045 123.810 105.375 ;
        RECT 31.830 99.605 33.810 99.935 ;
        RECT 61.830 99.605 63.810 99.935 ;
        RECT 91.830 99.605 93.810 99.935 ;
        RECT 121.830 99.605 123.810 99.935 ;
        RECT 137.190 76.585 139.920 77.835 ;
        RECT 0.970 70.330 3.070 70.430 ;
        RECT 15.510 70.330 17.040 71.185 ;
        RECT 0.960 68.750 17.040 70.330 ;
        RECT 0.970 68.710 3.070 68.750 ;
        RECT 15.510 68.635 17.040 68.750 ;
      LAYER met4 ;
        RECT 1.000 70.435 3.000 220.760 ;
        RECT 31.820 99.530 33.820 211.530 ;
        RECT 61.820 99.530 63.820 211.530 ;
        RECT 91.820 99.530 93.820 211.530 ;
        RECT 121.820 99.720 123.820 211.530 ;
        RECT 121.810 97.750 123.830 99.720 ;
        RECT 121.820 96.830 123.820 97.750 ;
        RECT 121.820 94.830 139.410 96.830 ;
        RECT 137.410 77.815 139.410 94.830 ;
        RECT 137.235 76.605 139.875 77.815 ;
        RECT 1.000 68.705 3.025 70.435 ;
        RECT 1.000 5.000 3.000 68.705 ;
        RECT 15.555 68.655 16.995 71.165 ;
      LAYER met5 ;
        RECT 14.420 205.290 128.060 207.290 ;
        RECT 14.420 175.290 128.060 177.290 ;
        RECT 14.420 145.290 128.060 147.290 ;
        RECT 14.420 115.290 128.060 117.290 ;
    END
  END vdd
  PIN ua[2]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER li1 ;
        RECT 137.765 20.110 137.935 30.150 ;
        RECT 22.275 19.685 27.275 19.855 ;
        RECT 33.555 19.685 38.555 19.855 ;
        RECT 44.845 19.665 49.845 19.835 ;
        RECT 56.065 19.665 61.065 19.835 ;
        RECT 67.265 19.665 72.265 19.835 ;
        RECT 78.555 19.655 83.555 19.825 ;
        RECT 89.795 19.675 94.795 19.845 ;
        RECT 101.005 19.695 106.005 19.865 ;
        RECT 112.205 19.735 117.205 19.905 ;
        RECT 123.415 19.755 128.415 19.925 ;
        RECT 132.705 19.725 137.705 19.895 ;
      LAYER met1 ;
        RECT 137.735 30.120 137.965 30.130 ;
        RECT 137.665 20.080 138.055 30.120 ;
        RECT 22.185 19.620 27.335 19.900 ;
        RECT 33.465 19.620 38.615 19.900 ;
        RECT 44.755 19.600 49.905 19.880 ;
        RECT 55.975 19.600 61.125 19.880 ;
        RECT 67.175 19.600 72.325 19.880 ;
        RECT 78.465 19.590 83.615 19.870 ;
        RECT 89.705 19.610 94.855 19.890 ;
        RECT 100.915 19.630 106.065 19.910 ;
        RECT 112.115 19.670 117.265 19.950 ;
        RECT 123.325 19.690 128.475 19.970 ;
        RECT 132.635 19.640 138.025 19.930 ;
        RECT 141.500 16.960 148.010 16.980 ;
        RECT 117.765 16.940 148.010 16.960 ;
        RECT 106.555 16.900 148.010 16.940 ;
        RECT 16.625 16.870 41.575 16.890 ;
        RECT 95.355 16.880 148.010 16.900 ;
        RECT 16.625 16.860 75.285 16.870 ;
        RECT 84.145 16.860 148.010 16.880 ;
        RECT 16.625 15.840 148.010 16.860 ;
        RECT 16.625 15.810 142.660 15.840 ;
        RECT 16.625 15.790 120.225 15.810 ;
        RECT 16.625 15.750 109.025 15.790 ;
        RECT 16.625 15.740 97.815 15.750 ;
        RECT 39.195 15.730 97.815 15.740 ;
        RECT 39.195 15.720 86.575 15.730 ;
        RECT 72.905 15.710 86.575 15.720 ;
        RECT 146.870 4.560 148.010 15.840 ;
        RECT 113.130 3.420 148.010 4.560 ;
        RECT 113.130 1.610 114.270 3.420 ;
        RECT 112.900 0.360 114.290 1.610 ;
        RECT 113.130 0.330 114.270 0.360 ;
      LAYER met2 ;
        RECT 22.235 19.570 27.285 19.950 ;
        RECT 33.515 19.570 38.565 19.950 ;
        RECT 23.915 16.790 25.845 19.570 ;
        RECT 35.195 16.790 37.125 19.570 ;
        RECT 44.805 19.550 49.855 19.930 ;
        RECT 56.025 19.550 61.075 19.930 ;
        RECT 67.225 19.550 72.275 19.930 ;
        RECT 23.335 15.940 26.045 16.790 ;
        RECT 34.615 15.940 37.325 16.790 ;
        RECT 46.485 16.770 48.415 19.550 ;
        RECT 57.705 16.770 59.635 19.550 ;
        RECT 68.905 16.770 70.835 19.550 ;
        RECT 78.515 19.540 83.565 19.920 ;
        RECT 89.755 19.560 94.805 19.940 ;
        RECT 100.965 19.580 106.015 19.960 ;
        RECT 112.165 19.620 117.215 20.000 ;
        RECT 123.375 19.640 128.425 20.020 ;
        RECT 137.715 19.980 138.005 30.170 ;
        RECT 45.905 15.920 48.615 16.770 ;
        RECT 57.125 15.920 59.835 16.770 ;
        RECT 68.325 15.920 71.035 16.770 ;
        RECT 80.195 16.760 82.125 19.540 ;
        RECT 91.435 16.780 93.365 19.560 ;
        RECT 102.645 16.800 104.575 19.580 ;
        RECT 113.845 16.840 115.775 19.620 ;
        RECT 125.055 16.860 126.985 19.640 ;
        RECT 132.685 19.590 138.005 19.980 ;
        RECT 137.715 16.940 138.005 19.590 ;
        RECT 79.615 15.910 82.325 16.760 ;
        RECT 90.855 15.930 93.565 16.780 ;
        RECT 102.065 15.950 104.775 16.800 ;
        RECT 113.265 15.990 115.975 16.840 ;
        RECT 124.475 16.010 127.185 16.860 ;
        RECT 137.395 15.890 138.295 16.940 ;
        RECT 137.715 15.720 138.005 15.890 ;
        RECT 112.950 0.310 114.240 1.660 ;
      LAYER met3 ;
        RECT 112.900 0.335 114.290 1.635 ;
      LAYER met4 ;
        RECT 112.945 0.355 114.245 1.615 ;
        RECT 113.170 0.000 114.070 0.355 ;
    END
  END ua[2]
  PIN ion
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER li1 ;
        RECT 28.205 47.015 28.375 52.055 ;
        RECT 39.405 47.025 39.575 52.065 ;
        RECT 50.625 46.995 50.795 52.035 ;
        RECT 61.875 46.975 62.045 52.015 ;
        RECT 73.095 46.965 73.265 52.005 ;
        RECT 84.335 46.955 84.505 51.995 ;
        RECT 95.585 46.965 95.755 52.005 ;
        RECT 106.865 46.955 107.035 51.995 ;
        RECT 118.135 46.955 118.305 51.995 ;
        RECT 129.385 46.955 129.555 51.995 ;
        RECT 20.365 33.355 20.535 38.395 ;
        RECT 31.645 33.355 31.815 38.395 ;
        RECT 42.935 33.335 43.105 38.375 ;
        RECT 54.155 33.335 54.325 38.375 ;
        RECT 65.355 33.335 65.525 38.375 ;
        RECT 76.645 33.325 76.815 38.365 ;
        RECT 87.885 33.345 88.055 38.385 ;
        RECT 99.095 33.365 99.265 38.405 ;
        RECT 110.295 33.405 110.465 38.445 ;
        RECT 121.505 33.425 121.675 38.465 ;
      LAYER met1 ;
        RECT 28.175 51.940 28.405 52.035 ;
        RECT 39.375 51.950 39.605 52.045 ;
        RECT 28.115 46.970 28.545 51.940 ;
        RECT 39.315 46.980 39.745 51.950 ;
        RECT 50.595 51.920 50.825 52.015 ;
        RECT 50.535 46.950 50.965 51.920 ;
        RECT 61.845 51.900 62.075 51.995 ;
        RECT 61.785 46.930 62.215 51.900 ;
        RECT 73.065 51.890 73.295 51.985 ;
        RECT 73.005 46.920 73.435 51.890 ;
        RECT 84.305 51.880 84.535 51.975 ;
        RECT 95.555 51.890 95.785 51.985 ;
        RECT 84.245 46.910 84.675 51.880 ;
        RECT 95.495 46.920 95.925 51.890 ;
        RECT 106.835 51.880 107.065 51.975 ;
        RECT 118.105 51.880 118.335 51.975 ;
        RECT 129.355 51.880 129.585 51.975 ;
        RECT 106.775 46.910 107.205 51.880 ;
        RECT 118.045 46.910 118.475 51.880 ;
        RECT 129.295 46.910 129.725 51.880 ;
        RECT 29.015 43.330 41.185 43.340 ;
        RECT 17.815 43.310 41.185 43.330 ;
        RECT 142.830 43.320 144.150 43.340 ;
        RECT 17.815 43.290 52.405 43.310 ;
        RECT 141.630 43.300 144.150 43.320 ;
        RECT 17.815 43.280 63.655 43.290 ;
        RECT 119.895 43.280 144.150 43.300 ;
        RECT 17.815 43.270 74.875 43.280 ;
        RECT 85.195 43.270 97.365 43.280 ;
        RECT 108.685 43.270 144.150 43.280 ;
        RECT 17.815 42.180 144.150 43.270 ;
        RECT 18.755 42.150 142.250 42.180 ;
        RECT 18.755 42.120 131.165 42.150 ;
        RECT 18.755 42.090 109.655 42.120 ;
        RECT 18.755 42.080 98.445 42.090 ;
        RECT 41.325 42.070 98.445 42.080 ;
        RECT 142.830 42.070 144.150 42.180 ;
        RECT 41.325 42.060 87.205 42.070 ;
        RECT 75.035 42.050 87.205 42.060 ;
        RECT 20.195 33.470 20.625 38.440 ;
        RECT 31.475 33.470 31.905 38.440 ;
        RECT 20.335 33.375 20.565 33.470 ;
        RECT 31.615 33.375 31.845 33.470 ;
        RECT 42.765 33.450 43.195 38.420 ;
        RECT 53.985 33.450 54.415 38.420 ;
        RECT 65.185 33.450 65.615 38.420 ;
        RECT 42.905 33.355 43.135 33.450 ;
        RECT 54.125 33.355 54.355 33.450 ;
        RECT 65.325 33.355 65.555 33.450 ;
        RECT 76.475 33.440 76.905 38.410 ;
        RECT 87.715 33.460 88.145 38.430 ;
        RECT 98.925 33.480 99.355 38.450 ;
        RECT 110.125 33.520 110.555 38.490 ;
        RECT 121.335 33.540 121.765 38.510 ;
        RECT 142.850 37.630 144.170 38.900 ;
        RECT 76.615 33.345 76.845 33.440 ;
        RECT 87.855 33.365 88.085 33.460 ;
        RECT 99.065 33.385 99.295 33.480 ;
        RECT 110.265 33.425 110.495 33.520 ;
        RECT 121.475 33.445 121.705 33.540 ;
        RECT 142.940 19.110 144.080 37.630 ;
        RECT 142.890 17.990 144.140 19.110 ;
        RECT 142.905 15.040 144.045 15.050 ;
        RECT 142.850 13.920 144.100 15.040 ;
        RECT 142.905 8.580 144.045 13.920 ;
        RECT 74.420 7.440 144.045 8.580 ;
        RECT 74.420 1.410 75.560 7.440 ;
        RECT 74.290 0.160 75.680 1.410 ;
      LAYER met2 ;
        RECT 28.165 46.920 28.495 51.990 ;
        RECT 39.365 46.930 39.695 52.000 ;
        RECT 28.215 44.930 28.495 46.920 ;
        RECT 39.415 44.940 39.695 46.930 ;
        RECT 50.585 46.900 50.915 51.970 ;
        RECT 28.215 43.200 28.515 44.930 ;
        RECT 39.415 43.210 39.715 44.940 ;
        RECT 50.635 44.910 50.915 46.900 ;
        RECT 61.835 46.880 62.165 51.950 ;
        RECT 19.865 42.210 21.245 42.780 ;
        RECT 27.495 42.630 28.875 43.200 ;
        RECT 31.145 42.210 32.525 42.780 ;
        RECT 38.695 42.640 40.075 43.210 ;
        RECT 50.635 43.180 50.935 44.910 ;
        RECT 61.885 44.890 62.165 46.880 ;
        RECT 73.055 46.870 73.385 51.940 ;
        RECT 20.225 40.480 20.525 42.210 ;
        RECT 31.505 40.480 31.805 42.210 ;
        RECT 42.435 42.190 43.815 42.760 ;
        RECT 49.915 42.610 51.295 43.180 ;
        RECT 61.885 43.160 62.185 44.890 ;
        RECT 73.105 44.880 73.385 46.870 ;
        RECT 84.295 46.860 84.625 51.930 ;
        RECT 95.545 46.870 95.875 51.940 ;
        RECT 53.655 42.190 55.035 42.760 ;
        RECT 61.165 42.590 62.545 43.160 ;
        RECT 73.105 43.150 73.405 44.880 ;
        RECT 84.345 44.870 84.625 46.860 ;
        RECT 95.595 44.880 95.875 46.870 ;
        RECT 106.825 46.860 107.155 51.930 ;
        RECT 118.095 46.860 118.425 51.930 ;
        RECT 129.345 46.860 129.675 51.930 ;
        RECT 64.855 42.190 66.235 42.760 ;
        RECT 72.385 42.580 73.765 43.150 ;
        RECT 84.345 43.140 84.645 44.870 ;
        RECT 95.595 43.150 95.895 44.880 ;
        RECT 106.875 44.870 107.155 46.860 ;
        RECT 118.145 44.870 118.425 46.860 ;
        RECT 129.395 44.870 129.675 46.860 ;
        RECT 20.245 38.490 20.525 40.480 ;
        RECT 31.525 38.490 31.805 40.480 ;
        RECT 42.795 40.460 43.095 42.190 ;
        RECT 54.015 40.460 54.315 42.190 ;
        RECT 65.215 40.460 65.515 42.190 ;
        RECT 76.145 42.180 77.525 42.750 ;
        RECT 83.625 42.570 85.005 43.140 ;
        RECT 87.385 42.200 88.765 42.770 ;
        RECT 94.875 42.580 96.255 43.150 ;
        RECT 106.875 43.140 107.175 44.870 ;
        RECT 118.145 43.140 118.445 44.870 ;
        RECT 129.395 43.140 129.695 44.870 ;
        RECT 98.595 42.220 99.975 42.790 ;
        RECT 106.155 42.570 107.535 43.140 ;
        RECT 109.795 42.260 111.175 42.830 ;
        RECT 117.425 42.570 118.805 43.140 ;
        RECT 121.005 42.280 122.385 42.850 ;
        RECT 128.675 42.570 130.055 43.140 ;
        RECT 20.245 33.420 20.575 38.490 ;
        RECT 31.525 33.420 31.855 38.490 ;
        RECT 42.815 38.470 43.095 40.460 ;
        RECT 54.035 38.470 54.315 40.460 ;
        RECT 65.235 38.470 65.515 40.460 ;
        RECT 76.505 40.450 76.805 42.180 ;
        RECT 87.745 40.470 88.045 42.200 ;
        RECT 98.955 40.490 99.255 42.220 ;
        RECT 110.155 40.530 110.455 42.260 ;
        RECT 121.365 40.550 121.665 42.280 ;
        RECT 142.880 42.020 144.100 43.390 ;
        RECT 42.815 33.400 43.145 38.470 ;
        RECT 54.035 33.400 54.365 38.470 ;
        RECT 65.235 33.400 65.565 38.470 ;
        RECT 76.525 38.460 76.805 40.450 ;
        RECT 87.765 38.480 88.045 40.470 ;
        RECT 98.975 38.500 99.255 40.490 ;
        RECT 110.175 38.540 110.455 40.530 ;
        RECT 121.385 38.560 121.665 40.550 ;
        RECT 142.940 38.950 144.100 42.020 ;
        RECT 76.525 33.390 76.855 38.460 ;
        RECT 87.765 33.410 88.095 38.480 ;
        RECT 98.975 33.430 99.305 38.500 ;
        RECT 110.175 33.470 110.505 38.540 ;
        RECT 121.385 33.490 121.715 38.560 ;
        RECT 142.900 37.580 144.120 38.950 ;
        RECT 142.940 17.940 144.090 19.160 ;
        RECT 142.940 15.090 144.050 17.940 ;
        RECT 142.900 13.870 144.050 15.090 ;
        RECT 74.340 0.110 75.630 1.460 ;
      LAYER met3 ;
        RECT 74.290 0.135 75.680 1.435 ;
      LAYER met4 ;
        RECT 74.335 0.155 75.635 1.415 ;
        RECT 74.530 0.000 75.430 0.155 ;
    END
  END ion
  PIN vss
    ANTENNAGATEAREA 1225.708130 ;
    ANTENNADIFFAREA 525.223694 ;
    PORT
      LAYER pwell ;
        RECT 24.335 210.315 24.765 211.100 ;
        RECT 37.215 210.315 37.645 211.100 ;
        RECT 50.095 210.315 50.525 211.100 ;
        RECT 62.975 210.315 63.405 211.100 ;
        RECT 75.855 210.315 76.285 211.100 ;
        RECT 88.735 210.315 89.165 211.100 ;
        RECT 101.615 210.315 102.045 211.100 ;
        RECT 114.495 210.315 114.925 211.100 ;
        RECT 24.335 206.040 24.765 206.825 ;
        RECT 50.095 206.040 50.525 206.825 ;
        RECT 75.855 206.040 76.285 206.825 ;
        RECT 101.615 206.040 102.045 206.825 ;
        RECT 37.215 204.875 37.645 205.660 ;
        RECT 62.975 204.875 63.405 205.660 ;
        RECT 88.735 204.875 89.165 205.660 ;
        RECT 114.495 204.875 114.925 205.660 ;
        RECT 24.335 200.600 24.765 201.385 ;
        RECT 50.095 200.600 50.525 201.385 ;
        RECT 75.855 200.600 76.285 201.385 ;
        RECT 101.615 200.600 102.045 201.385 ;
        RECT 37.215 199.435 37.645 200.220 ;
        RECT 62.975 199.435 63.405 200.220 ;
        RECT 88.735 199.435 89.165 200.220 ;
        RECT 114.495 199.435 114.925 200.220 ;
        RECT 24.335 195.160 24.765 195.945 ;
        RECT 50.095 195.160 50.525 195.945 ;
        RECT 75.855 195.160 76.285 195.945 ;
        RECT 101.615 195.160 102.045 195.945 ;
        RECT 37.215 193.995 37.645 194.780 ;
        RECT 62.975 193.995 63.405 194.780 ;
        RECT 88.735 193.995 89.165 194.780 ;
        RECT 114.495 193.995 114.925 194.780 ;
        RECT 24.335 189.720 24.765 190.505 ;
        RECT 50.095 189.720 50.525 190.505 ;
        RECT 75.855 189.720 76.285 190.505 ;
        RECT 101.615 189.720 102.045 190.505 ;
        RECT 37.215 188.555 37.645 189.340 ;
        RECT 62.975 188.555 63.405 189.340 ;
        RECT 88.735 188.555 89.165 189.340 ;
        RECT 114.495 188.555 114.925 189.340 ;
        RECT 24.335 184.280 24.765 185.065 ;
        RECT 50.095 184.280 50.525 185.065 ;
        RECT 75.855 184.280 76.285 185.065 ;
        RECT 101.615 184.280 102.045 185.065 ;
        RECT 37.215 183.115 37.645 183.900 ;
        RECT 62.975 183.115 63.405 183.900 ;
        RECT 88.735 183.115 89.165 183.900 ;
        RECT 114.495 183.115 114.925 183.900 ;
        RECT 24.335 178.840 24.765 179.625 ;
        RECT 50.095 178.840 50.525 179.625 ;
        RECT 75.855 178.840 76.285 179.625 ;
        RECT 101.615 178.840 102.045 179.625 ;
        RECT 37.215 177.675 37.645 178.460 ;
        RECT 62.975 177.675 63.405 178.460 ;
        RECT 88.735 177.675 89.165 178.460 ;
        RECT 114.495 177.675 114.925 178.460 ;
        RECT 24.335 173.400 24.765 174.185 ;
        RECT 50.095 173.400 50.525 174.185 ;
        RECT 75.855 173.400 76.285 174.185 ;
        RECT 101.615 173.400 102.045 174.185 ;
        RECT 37.215 172.235 37.645 173.020 ;
        RECT 62.975 172.235 63.405 173.020 ;
        RECT 88.735 172.235 89.165 173.020 ;
        RECT 114.495 172.235 114.925 173.020 ;
        RECT 24.335 167.960 24.765 168.745 ;
        RECT 50.095 167.960 50.525 168.745 ;
        RECT 75.855 167.960 76.285 168.745 ;
        RECT 101.615 167.960 102.045 168.745 ;
        RECT 37.215 166.795 37.645 167.580 ;
        RECT 62.975 166.795 63.405 167.580 ;
        RECT 88.735 166.795 89.165 167.580 ;
        RECT 114.495 166.795 114.925 167.580 ;
        RECT 24.335 162.520 24.765 163.305 ;
        RECT 50.095 162.520 50.525 163.305 ;
        RECT 75.855 162.520 76.285 163.305 ;
        RECT 101.615 162.520 102.045 163.305 ;
        RECT 37.215 161.355 37.645 162.140 ;
        RECT 62.975 161.355 63.405 162.140 ;
        RECT 88.735 161.355 89.165 162.140 ;
        RECT 114.495 161.355 114.925 162.140 ;
        RECT 24.335 157.080 24.765 157.865 ;
        RECT 50.095 157.080 50.525 157.865 ;
        RECT 75.855 157.080 76.285 157.865 ;
        RECT 101.615 157.080 102.045 157.865 ;
        RECT 37.215 155.915 37.645 156.700 ;
        RECT 62.975 155.915 63.405 156.700 ;
        RECT 88.735 155.915 89.165 156.700 ;
        RECT 114.495 155.915 114.925 156.700 ;
        RECT 24.335 151.640 24.765 152.425 ;
        RECT 50.095 151.640 50.525 152.425 ;
        RECT 75.855 151.640 76.285 152.425 ;
        RECT 101.615 151.640 102.045 152.425 ;
        RECT 37.215 150.475 37.645 151.260 ;
        RECT 62.975 150.475 63.405 151.260 ;
        RECT 88.735 150.475 89.165 151.260 ;
        RECT 114.495 150.475 114.925 151.260 ;
        RECT 24.335 146.200 24.765 146.985 ;
        RECT 50.095 146.200 50.525 146.985 ;
        RECT 75.855 146.200 76.285 146.985 ;
        RECT 101.615 146.200 102.045 146.985 ;
        RECT 37.215 145.035 37.645 145.820 ;
        RECT 62.975 145.035 63.405 145.820 ;
        RECT 88.735 145.035 89.165 145.820 ;
        RECT 114.495 145.035 114.925 145.820 ;
        RECT 24.335 140.760 24.765 141.545 ;
        RECT 50.095 140.760 50.525 141.545 ;
        RECT 75.855 140.760 76.285 141.545 ;
        RECT 101.615 140.760 102.045 141.545 ;
        RECT 37.215 139.595 37.645 140.380 ;
        RECT 62.975 139.595 63.405 140.380 ;
        RECT 88.735 139.595 89.165 140.380 ;
        RECT 114.495 139.595 114.925 140.380 ;
        RECT 24.335 135.320 24.765 136.105 ;
        RECT 50.095 135.320 50.525 136.105 ;
        RECT 75.855 135.320 76.285 136.105 ;
        RECT 101.615 135.320 102.045 136.105 ;
        RECT 37.215 134.155 37.645 134.940 ;
        RECT 62.975 134.155 63.405 134.940 ;
        RECT 88.735 134.155 89.165 134.940 ;
        RECT 114.495 134.155 114.925 134.940 ;
        RECT 24.335 129.880 24.765 130.665 ;
        RECT 50.095 129.880 50.525 130.665 ;
        RECT 75.855 129.880 76.285 130.665 ;
        RECT 101.615 129.880 102.045 130.665 ;
        RECT 37.215 128.715 37.645 129.500 ;
        RECT 62.975 128.715 63.405 129.500 ;
        RECT 88.735 128.715 89.165 129.500 ;
        RECT 114.495 128.715 114.925 129.500 ;
        RECT 24.335 124.440 24.765 125.225 ;
        RECT 50.095 124.440 50.525 125.225 ;
        RECT 75.855 124.440 76.285 125.225 ;
        RECT 101.615 124.440 102.045 125.225 ;
        RECT 37.215 123.275 37.645 124.060 ;
        RECT 62.975 123.275 63.405 124.060 ;
        RECT 88.735 123.275 89.165 124.060 ;
        RECT 114.495 123.275 114.925 124.060 ;
        RECT 24.335 119.000 24.765 119.785 ;
        RECT 50.095 119.000 50.525 119.785 ;
        RECT 75.855 119.000 76.285 119.785 ;
        RECT 101.615 119.000 102.045 119.785 ;
        RECT 37.215 117.835 37.645 118.620 ;
        RECT 62.975 117.835 63.405 118.620 ;
        RECT 88.735 117.835 89.165 118.620 ;
        RECT 114.495 117.835 114.925 118.620 ;
        RECT 24.335 113.560 24.765 114.345 ;
        RECT 50.095 113.560 50.525 114.345 ;
        RECT 75.855 113.560 76.285 114.345 ;
        RECT 101.615 113.560 102.045 114.345 ;
        RECT 37.215 112.395 37.645 113.180 ;
        RECT 62.975 112.395 63.405 113.180 ;
        RECT 88.735 112.395 89.165 113.180 ;
        RECT 114.495 112.395 114.925 113.180 ;
        RECT 24.335 108.120 24.765 108.905 ;
        RECT 50.095 108.120 50.525 108.905 ;
        RECT 75.855 108.120 76.285 108.905 ;
        RECT 101.615 108.120 102.045 108.905 ;
        RECT 37.215 106.955 37.645 107.740 ;
        RECT 62.975 106.955 63.405 107.740 ;
        RECT 88.735 106.955 89.165 107.740 ;
        RECT 114.495 106.955 114.925 107.740 ;
        RECT 24.335 102.680 24.765 103.465 ;
        RECT 50.095 102.680 50.525 103.465 ;
        RECT 75.855 102.680 76.285 103.465 ;
        RECT 101.615 102.680 102.045 103.465 ;
        RECT 24.335 101.515 24.765 102.300 ;
        RECT 37.215 101.515 37.645 102.300 ;
        RECT 50.095 101.515 50.525 102.300 ;
        RECT 62.975 101.515 63.405 102.300 ;
        RECT 75.855 101.515 76.285 102.300 ;
        RECT 88.735 101.515 89.165 102.300 ;
        RECT 101.615 101.515 102.045 102.300 ;
        RECT 114.495 101.515 114.925 102.300 ;
        RECT 20.555 45.340 22.915 48.340 ;
        RECT 31.755 45.350 34.115 48.350 ;
        RECT 42.975 45.320 45.335 48.320 ;
        RECT 54.225 45.300 56.585 48.300 ;
        RECT 65.445 45.290 67.805 48.290 ;
        RECT 76.685 45.280 79.045 48.280 ;
        RECT 87.935 45.290 90.295 48.290 ;
        RECT 99.215 45.280 101.575 48.280 ;
        RECT 110.485 45.280 112.845 48.280 ;
        RECT 121.735 45.280 124.095 48.280 ;
        RECT 25.825 37.070 28.185 40.070 ;
        RECT 37.105 37.070 39.465 40.070 ;
        RECT 48.395 37.050 50.755 40.050 ;
        RECT 59.615 37.050 61.975 40.050 ;
        RECT 70.815 37.050 73.175 40.050 ;
        RECT 82.105 37.040 84.465 40.040 ;
        RECT 93.345 37.060 95.705 40.060 ;
        RECT 104.555 37.080 106.915 40.080 ;
        RECT 115.755 37.120 118.115 40.120 ;
        RECT 126.965 37.140 129.325 40.140 ;
      LAYER li1 ;
        RECT 14.660 211.205 127.820 211.375 ;
        RECT 14.745 210.455 15.955 211.205 ;
        RECT 14.745 209.915 15.265 210.455 ;
        RECT 16.125 210.435 18.715 211.205 ;
        RECT 18.890 210.660 24.235 211.205 ;
        RECT 17.505 209.915 18.715 210.435 ;
        RECT 22.310 209.830 22.650 210.660 ;
        RECT 24.405 210.480 24.695 211.205 ;
        RECT 24.865 210.455 26.075 211.205 ;
        RECT 26.250 210.660 31.595 211.205 ;
        RECT 31.770 210.660 37.115 211.205 ;
        RECT 25.555 209.915 26.075 210.455 ;
        RECT 29.670 209.830 30.010 210.660 ;
        RECT 35.190 209.830 35.530 210.660 ;
        RECT 37.285 210.480 37.575 211.205 ;
        RECT 37.745 210.455 38.955 211.205 ;
        RECT 39.130 210.660 44.475 211.205 ;
        RECT 44.650 210.660 49.995 211.205 ;
        RECT 38.435 209.915 38.955 210.455 ;
        RECT 42.550 209.830 42.890 210.660 ;
        RECT 48.070 209.830 48.410 210.660 ;
        RECT 50.165 210.480 50.455 211.205 ;
        RECT 50.625 210.455 51.835 211.205 ;
        RECT 52.010 210.660 57.355 211.205 ;
        RECT 57.530 210.660 62.875 211.205 ;
        RECT 51.315 209.915 51.835 210.455 ;
        RECT 55.430 209.830 55.770 210.660 ;
        RECT 60.950 209.830 61.290 210.660 ;
        RECT 63.045 210.480 63.335 211.205 ;
        RECT 63.505 210.455 64.715 211.205 ;
        RECT 64.890 210.660 70.235 211.205 ;
        RECT 70.410 210.660 75.755 211.205 ;
        RECT 64.195 209.915 64.715 210.455 ;
        RECT 68.310 209.830 68.650 210.660 ;
        RECT 73.830 209.830 74.170 210.660 ;
        RECT 75.925 210.480 76.215 211.205 ;
        RECT 76.385 210.455 77.595 211.205 ;
        RECT 77.770 210.660 83.115 211.205 ;
        RECT 83.290 210.660 88.635 211.205 ;
        RECT 77.075 209.915 77.595 210.455 ;
        RECT 81.190 209.830 81.530 210.660 ;
        RECT 86.710 209.830 87.050 210.660 ;
        RECT 88.805 210.480 89.095 211.205 ;
        RECT 89.265 210.455 90.475 211.205 ;
        RECT 90.650 210.660 95.995 211.205 ;
        RECT 96.170 210.660 101.515 211.205 ;
        RECT 89.955 209.915 90.475 210.455 ;
        RECT 94.070 209.830 94.410 210.660 ;
        RECT 99.590 209.830 99.930 210.660 ;
        RECT 101.685 210.480 101.975 211.205 ;
        RECT 102.145 210.455 103.355 211.205 ;
        RECT 103.530 210.660 108.875 211.205 ;
        RECT 109.050 210.660 114.395 211.205 ;
        RECT 102.835 209.915 103.355 210.455 ;
        RECT 106.950 209.830 107.290 210.660 ;
        RECT 112.470 209.830 112.810 210.660 ;
        RECT 114.565 210.480 114.855 211.205 ;
        RECT 115.490 210.660 120.835 211.205 ;
        RECT 121.010 210.660 126.355 211.205 ;
        RECT 118.910 209.830 119.250 210.660 ;
        RECT 124.430 209.830 124.770 210.660 ;
        RECT 126.525 210.455 127.735 211.205 ;
        RECT 127.215 209.915 127.735 210.455 ;
        RECT 14.745 206.685 15.265 207.225 ;
        RECT 17.505 206.705 18.715 207.225 ;
        RECT 14.745 205.935 15.955 206.685 ;
        RECT 16.125 205.935 18.715 206.705 ;
        RECT 22.310 206.480 22.650 207.310 ;
        RECT 26.705 206.705 27.915 207.225 ;
        RECT 18.890 205.935 24.235 206.480 ;
        RECT 24.405 205.935 24.695 206.660 ;
        RECT 25.325 205.935 27.915 206.705 ;
        RECT 31.510 206.480 31.850 207.310 ;
        RECT 37.030 206.480 37.370 207.310 ;
        RECT 42.550 206.480 42.890 207.310 ;
        RECT 48.070 206.480 48.410 207.310 ;
        RECT 51.545 206.705 52.295 207.225 ;
        RECT 28.090 205.935 33.435 206.480 ;
        RECT 33.610 205.935 38.955 206.480 ;
        RECT 39.130 205.935 44.475 206.480 ;
        RECT 44.650 205.935 49.995 206.480 ;
        RECT 50.165 205.935 50.455 206.660 ;
        RECT 50.625 205.935 52.295 206.705 ;
        RECT 55.890 206.480 56.230 207.310 ;
        RECT 61.410 206.480 61.750 207.310 ;
        RECT 66.930 206.480 67.270 207.310 ;
        RECT 72.450 206.480 72.790 207.310 ;
        RECT 52.470 205.935 57.815 206.480 ;
        RECT 57.990 205.935 63.335 206.480 ;
        RECT 63.510 205.935 68.855 206.480 ;
        RECT 69.030 205.935 74.375 206.480 ;
        RECT 74.585 205.935 74.815 206.755 ;
        RECT 75.485 205.935 75.695 206.755 ;
        RECT 77.075 206.685 77.595 207.225 ;
        RECT 75.925 205.935 76.215 206.660 ;
        RECT 76.385 205.935 77.595 206.685 ;
        RECT 78.655 205.935 79.005 206.325 ;
        RECT 79.675 205.935 79.845 206.755 ;
        RECT 83.305 206.705 84.955 207.225 ;
        RECT 81.445 205.935 84.955 206.705 ;
        RECT 88.550 206.480 88.890 207.310 ;
        RECT 94.070 206.480 94.410 207.310 ;
        RECT 99.590 206.480 99.930 207.310 ;
        RECT 103.525 206.705 104.275 207.225 ;
        RECT 85.130 205.935 90.475 206.480 ;
        RECT 90.650 205.935 95.995 206.480 ;
        RECT 96.170 205.935 101.515 206.480 ;
        RECT 101.685 205.935 101.975 206.660 ;
        RECT 102.605 205.935 104.275 206.705 ;
        RECT 107.870 206.480 108.210 207.310 ;
        RECT 113.390 206.480 113.730 207.310 ;
        RECT 118.910 206.480 119.250 207.310 ;
        RECT 124.430 206.480 124.770 207.310 ;
        RECT 127.215 206.685 127.735 207.225 ;
        RECT 104.450 205.935 109.795 206.480 ;
        RECT 109.970 205.935 115.315 206.480 ;
        RECT 115.490 205.935 120.835 206.480 ;
        RECT 121.010 205.935 126.355 206.480 ;
        RECT 126.525 205.935 127.735 206.685 ;
        RECT 14.660 205.765 127.820 205.935 ;
        RECT 14.745 205.015 15.955 205.765 ;
        RECT 14.745 204.475 15.265 205.015 ;
        RECT 17.045 204.995 20.555 205.765 ;
        RECT 20.730 205.220 26.075 205.765 ;
        RECT 26.250 205.220 31.595 205.765 ;
        RECT 31.770 205.220 37.115 205.765 ;
        RECT 18.905 204.475 20.555 204.995 ;
        RECT 24.150 204.390 24.490 205.220 ;
        RECT 29.670 204.390 30.010 205.220 ;
        RECT 35.190 204.390 35.530 205.220 ;
        RECT 37.285 205.040 37.575 205.765 ;
        RECT 38.205 204.995 40.795 205.765 ;
        RECT 40.970 205.220 46.315 205.765 ;
        RECT 46.490 205.220 51.835 205.765 ;
        RECT 52.010 205.220 57.355 205.765 ;
        RECT 57.530 205.220 62.875 205.765 ;
        RECT 39.585 204.475 40.795 204.995 ;
        RECT 44.390 204.390 44.730 205.220 ;
        RECT 49.910 204.390 50.250 205.220 ;
        RECT 55.430 204.390 55.770 205.220 ;
        RECT 60.950 204.390 61.290 205.220 ;
        RECT 63.045 205.040 63.335 205.765 ;
        RECT 63.505 204.995 65.175 205.765 ;
        RECT 64.425 204.475 65.175 204.995 ;
        RECT 65.405 204.945 65.615 205.765 ;
        RECT 66.285 204.945 66.515 205.765 ;
        RECT 67.225 204.945 67.455 205.765 ;
        RECT 68.125 204.945 68.335 205.765 ;
        RECT 68.995 205.305 69.300 205.765 ;
        RECT 70.785 205.325 70.975 205.765 ;
        RECT 72.875 205.305 73.205 205.765 ;
        RECT 75.805 205.405 76.135 205.765 ;
        RECT 76.835 205.385 77.165 205.765 ;
        RECT 78.195 205.305 78.500 205.765 ;
        RECT 79.985 205.325 80.175 205.765 ;
        RECT 82.075 205.305 82.405 205.765 ;
        RECT 85.005 205.405 85.335 205.765 ;
        RECT 86.035 205.385 86.365 205.765 ;
        RECT 86.965 204.995 88.635 205.765 ;
        RECT 88.805 205.040 89.095 205.765 ;
        RECT 89.725 204.995 92.315 205.765 ;
        RECT 92.490 205.220 97.835 205.765 ;
        RECT 98.010 205.220 103.355 205.765 ;
        RECT 103.530 205.220 108.875 205.765 ;
        RECT 109.050 205.220 114.395 205.765 ;
        RECT 87.885 204.475 88.635 204.995 ;
        RECT 91.105 204.475 92.315 204.995 ;
        RECT 95.910 204.390 96.250 205.220 ;
        RECT 101.430 204.390 101.770 205.220 ;
        RECT 106.950 204.390 107.290 205.220 ;
        RECT 112.470 204.390 112.810 205.220 ;
        RECT 114.565 205.040 114.855 205.765 ;
        RECT 115.490 205.220 120.835 205.765 ;
        RECT 121.010 205.220 126.355 205.765 ;
        RECT 118.910 204.390 119.250 205.220 ;
        RECT 124.430 204.390 124.770 205.220 ;
        RECT 126.525 205.015 127.735 205.765 ;
        RECT 127.215 204.475 127.735 205.015 ;
        RECT 14.745 201.245 15.265 201.785 ;
        RECT 17.505 201.265 18.715 201.785 ;
        RECT 14.745 200.495 15.955 201.245 ;
        RECT 16.125 200.495 18.715 201.265 ;
        RECT 22.310 201.040 22.650 201.870 ;
        RECT 26.705 201.265 27.915 201.785 ;
        RECT 18.890 200.495 24.235 201.040 ;
        RECT 24.405 200.495 24.695 201.220 ;
        RECT 25.325 200.495 27.915 201.265 ;
        RECT 31.510 201.040 31.850 201.870 ;
        RECT 37.030 201.040 37.370 201.870 ;
        RECT 42.550 201.040 42.890 201.870 ;
        RECT 48.070 201.040 48.410 201.870 ;
        RECT 52.945 201.265 54.595 201.785 ;
        RECT 28.090 200.495 33.435 201.040 ;
        RECT 33.610 200.495 38.955 201.040 ;
        RECT 39.130 200.495 44.475 201.040 ;
        RECT 44.650 200.495 49.995 201.040 ;
        RECT 50.165 200.495 50.455 201.220 ;
        RECT 51.085 200.495 54.595 201.265 ;
        RECT 58.190 201.040 58.530 201.870 ;
        RECT 54.770 200.495 60.115 201.040 ;
        RECT 60.715 200.495 61.045 200.875 ;
        RECT 61.745 200.495 62.075 200.855 ;
        RECT 64.675 200.495 65.005 200.955 ;
        RECT 66.905 200.495 67.095 200.935 ;
        RECT 68.535 200.495 68.705 201.305 ;
        RECT 69.375 200.495 69.545 200.965 ;
        RECT 70.215 200.495 70.385 200.965 ;
        RECT 71.335 200.495 71.610 200.975 ;
        RECT 72.195 200.495 72.530 200.895 ;
        RECT 73.180 200.495 73.510 200.875 ;
        RECT 74.110 200.495 74.370 201.335 ;
        RECT 75.235 201.245 75.755 201.785 ;
        RECT 89.725 201.265 90.475 201.785 ;
        RECT 74.545 200.495 75.755 201.245 ;
        RECT 75.925 200.495 76.215 201.220 ;
        RECT 76.855 200.495 77.130 200.975 ;
        RECT 77.715 200.495 78.050 200.895 ;
        RECT 78.665 200.495 78.995 200.875 ;
        RECT 80.035 200.495 80.340 200.955 ;
        RECT 81.825 200.495 82.015 200.935 ;
        RECT 83.915 200.495 84.245 200.955 ;
        RECT 86.845 200.495 87.175 200.855 ;
        RECT 87.875 200.495 88.205 200.875 ;
        RECT 88.805 200.495 90.475 201.265 ;
        RECT 94.070 201.040 94.410 201.870 ;
        RECT 99.590 201.040 99.930 201.870 ;
        RECT 103.525 201.265 104.275 201.785 ;
        RECT 90.650 200.495 95.995 201.040 ;
        RECT 96.170 200.495 101.515 201.040 ;
        RECT 101.685 200.495 101.975 201.220 ;
        RECT 102.605 200.495 104.275 201.265 ;
        RECT 107.870 201.040 108.210 201.870 ;
        RECT 113.390 201.040 113.730 201.870 ;
        RECT 118.910 201.040 119.250 201.870 ;
        RECT 124.430 201.040 124.770 201.870 ;
        RECT 127.215 201.245 127.735 201.785 ;
        RECT 104.450 200.495 109.795 201.040 ;
        RECT 109.970 200.495 115.315 201.040 ;
        RECT 115.490 200.495 120.835 201.040 ;
        RECT 121.010 200.495 126.355 201.040 ;
        RECT 126.525 200.495 127.735 201.245 ;
        RECT 14.660 200.325 127.820 200.495 ;
        RECT 14.745 199.575 15.955 200.325 ;
        RECT 14.745 199.035 15.265 199.575 ;
        RECT 17.045 199.555 20.555 200.325 ;
        RECT 20.730 199.780 26.075 200.325 ;
        RECT 26.250 199.780 31.595 200.325 ;
        RECT 31.770 199.780 37.115 200.325 ;
        RECT 18.905 199.035 20.555 199.555 ;
        RECT 24.150 198.950 24.490 199.780 ;
        RECT 29.670 198.950 30.010 199.780 ;
        RECT 35.190 198.950 35.530 199.780 ;
        RECT 37.285 199.600 37.575 200.325 ;
        RECT 38.205 199.555 40.795 200.325 ;
        RECT 40.970 199.780 46.315 200.325 ;
        RECT 46.490 199.780 51.835 200.325 ;
        RECT 52.010 199.780 57.355 200.325 ;
        RECT 57.530 199.780 62.875 200.325 ;
        RECT 39.585 199.035 40.795 199.555 ;
        RECT 44.390 198.950 44.730 199.780 ;
        RECT 49.910 198.950 50.250 199.780 ;
        RECT 55.430 198.950 55.770 199.780 ;
        RECT 60.950 198.950 61.290 199.780 ;
        RECT 63.045 199.600 63.335 200.325 ;
        RECT 63.965 199.555 65.635 200.325 ;
        RECT 66.245 199.945 66.575 200.325 ;
        RECT 67.695 199.945 68.025 200.325 ;
        RECT 69.935 199.945 70.265 200.325 ;
        RECT 71.295 199.945 71.625 200.325 ;
        RECT 74.395 199.945 74.725 200.325 ;
        RECT 76.020 199.865 76.345 200.325 ;
        RECT 78.135 199.865 78.405 200.325 ;
        RECT 79.575 199.785 79.825 200.325 ;
        RECT 64.885 199.035 65.635 199.555 ;
        RECT 82.345 199.525 82.655 200.325 ;
        RECT 82.885 199.505 83.095 200.325 ;
        RECT 83.765 199.505 83.995 200.325 ;
        RECT 84.245 199.505 84.475 200.325 ;
        RECT 85.145 199.505 85.355 200.325 ;
        RECT 86.045 199.555 88.635 200.325 ;
        RECT 88.805 199.600 89.095 200.325 ;
        RECT 89.725 199.555 92.315 200.325 ;
        RECT 92.490 199.780 97.835 200.325 ;
        RECT 98.010 199.780 103.355 200.325 ;
        RECT 103.530 199.780 108.875 200.325 ;
        RECT 109.050 199.780 114.395 200.325 ;
        RECT 87.425 199.035 88.635 199.555 ;
        RECT 91.105 199.035 92.315 199.555 ;
        RECT 95.910 198.950 96.250 199.780 ;
        RECT 101.430 198.950 101.770 199.780 ;
        RECT 106.950 198.950 107.290 199.780 ;
        RECT 112.470 198.950 112.810 199.780 ;
        RECT 114.565 199.600 114.855 200.325 ;
        RECT 115.490 199.780 120.835 200.325 ;
        RECT 121.010 199.780 126.355 200.325 ;
        RECT 118.910 198.950 119.250 199.780 ;
        RECT 124.430 198.950 124.770 199.780 ;
        RECT 126.525 199.575 127.735 200.325 ;
        RECT 127.215 199.035 127.735 199.575 ;
        RECT 14.745 195.805 15.265 196.345 ;
        RECT 17.505 195.825 18.715 196.345 ;
        RECT 14.745 195.055 15.955 195.805 ;
        RECT 16.125 195.055 18.715 195.825 ;
        RECT 22.310 195.600 22.650 196.430 ;
        RECT 26.705 195.825 27.915 196.345 ;
        RECT 18.890 195.055 24.235 195.600 ;
        RECT 24.405 195.055 24.695 195.780 ;
        RECT 25.325 195.055 27.915 195.825 ;
        RECT 31.510 195.600 31.850 196.430 ;
        RECT 37.030 195.600 37.370 196.430 ;
        RECT 42.550 195.600 42.890 196.430 ;
        RECT 48.070 195.600 48.410 196.430 ;
        RECT 51.545 195.825 52.295 196.345 ;
        RECT 28.090 195.055 33.435 195.600 ;
        RECT 33.610 195.055 38.955 195.600 ;
        RECT 39.130 195.055 44.475 195.600 ;
        RECT 44.650 195.055 49.995 195.600 ;
        RECT 50.165 195.055 50.455 195.780 ;
        RECT 50.625 195.055 52.295 195.825 ;
        RECT 52.525 195.055 52.735 195.875 ;
        RECT 53.405 195.055 53.635 195.875 ;
        RECT 54.765 195.825 55.515 196.345 ;
        RECT 53.845 195.055 55.515 195.825 ;
        RECT 55.745 195.055 55.955 195.875 ;
        RECT 56.625 195.055 56.855 195.875 ;
        RECT 57.755 195.805 58.275 196.345 ;
        RECT 57.065 195.055 58.275 195.805 ;
        RECT 61.870 195.600 62.210 196.430 ;
        RECT 67.390 195.600 67.730 196.430 ;
        RECT 58.450 195.055 63.795 195.600 ;
        RECT 63.970 195.055 69.315 195.600 ;
        RECT 69.915 195.055 70.165 195.595 ;
        RECT 72.295 195.055 72.625 195.455 ;
        RECT 74.175 195.055 74.505 195.455 ;
        RECT 75.925 195.055 76.215 195.780 ;
        RECT 83.030 195.600 83.370 196.430 ;
        RECT 88.550 195.600 88.890 196.430 ;
        RECT 94.070 195.600 94.410 196.430 ;
        RECT 99.590 195.600 99.930 196.430 ;
        RECT 77.470 195.055 77.710 195.565 ;
        RECT 78.400 195.055 78.615 195.565 ;
        RECT 79.610 195.055 84.955 195.600 ;
        RECT 85.130 195.055 90.475 195.600 ;
        RECT 90.650 195.055 95.995 195.600 ;
        RECT 96.170 195.055 101.515 195.600 ;
        RECT 101.685 195.055 101.975 195.780 ;
        RECT 105.570 195.600 105.910 196.430 ;
        RECT 102.150 195.055 107.495 195.600 ;
        RECT 107.705 195.055 107.935 195.875 ;
        RECT 108.605 195.055 108.815 195.875 ;
        RECT 119.625 195.825 120.835 196.345 ;
        RECT 109.475 195.055 109.780 195.515 ;
        RECT 111.265 195.055 111.455 195.495 ;
        RECT 113.355 195.055 113.685 195.515 ;
        RECT 116.285 195.055 116.615 195.415 ;
        RECT 117.315 195.055 117.645 195.435 ;
        RECT 118.245 195.055 120.835 195.825 ;
        RECT 124.430 195.600 124.770 196.430 ;
        RECT 127.215 195.805 127.735 196.345 ;
        RECT 121.010 195.055 126.355 195.600 ;
        RECT 126.525 195.055 127.735 195.805 ;
        RECT 14.660 194.885 127.820 195.055 ;
        RECT 14.745 194.135 15.955 194.885 ;
        RECT 14.745 193.595 15.265 194.135 ;
        RECT 17.045 194.115 20.555 194.885 ;
        RECT 20.730 194.340 26.075 194.885 ;
        RECT 26.250 194.340 31.595 194.885 ;
        RECT 31.770 194.340 37.115 194.885 ;
        RECT 18.905 193.595 20.555 194.115 ;
        RECT 24.150 193.510 24.490 194.340 ;
        RECT 29.670 193.510 30.010 194.340 ;
        RECT 35.190 193.510 35.530 194.340 ;
        RECT 37.285 194.160 37.575 194.885 ;
        RECT 38.210 194.340 43.555 194.885 ;
        RECT 44.155 194.505 44.485 194.885 ;
        RECT 45.185 194.525 45.515 194.885 ;
        RECT 48.115 194.425 48.445 194.885 ;
        RECT 50.345 194.445 50.535 194.885 ;
        RECT 52.020 194.425 52.325 194.885 ;
        RECT 53.355 194.425 53.660 194.885 ;
        RECT 55.145 194.445 55.335 194.885 ;
        RECT 57.235 194.425 57.565 194.885 ;
        RECT 60.165 194.525 60.495 194.885 ;
        RECT 61.195 194.505 61.525 194.885 ;
        RECT 41.630 193.510 41.970 194.340 ;
        RECT 63.045 194.160 63.335 194.885 ;
        RECT 63.965 194.115 65.635 194.885 ;
        RECT 64.885 193.595 65.635 194.115 ;
        RECT 65.865 194.065 66.075 194.885 ;
        RECT 66.745 194.065 66.975 194.885 ;
        RECT 67.185 194.135 68.395 194.885 ;
        RECT 67.875 193.595 68.395 194.135 ;
        RECT 68.565 194.115 72.075 194.885 ;
        RECT 70.425 193.595 72.075 194.115 ;
        RECT 72.245 194.065 72.505 194.885 ;
        RECT 73.615 194.485 73.945 194.885 ;
        RECT 74.455 194.485 74.830 194.885 ;
        RECT 75.930 194.485 76.305 194.885 ;
        RECT 76.815 194.485 77.145 194.885 ;
        RECT 78.255 194.065 78.515 194.885 ;
        RECT 79.150 194.340 84.495 194.885 ;
        RECT 85.405 194.350 85.915 194.885 ;
        RECT 87.875 194.485 88.205 194.885 ;
        RECT 82.570 193.510 82.910 194.340 ;
        RECT 88.805 194.160 89.095 194.885 ;
        RECT 89.785 194.065 89.995 194.885 ;
        RECT 90.665 194.065 90.895 194.885 ;
        RECT 92.005 194.505 92.335 194.885 ;
        RECT 93.405 194.115 95.995 194.885 ;
        RECT 94.785 193.595 95.995 194.115 ;
        RECT 96.205 194.065 96.435 194.885 ;
        RECT 97.105 194.065 97.315 194.885 ;
        RECT 97.975 194.425 98.280 194.885 ;
        RECT 99.765 194.445 99.955 194.885 ;
        RECT 101.855 194.425 102.185 194.885 ;
        RECT 104.785 194.525 105.115 194.885 ;
        RECT 105.815 194.505 106.145 194.885 ;
        RECT 107.300 194.425 107.625 194.885 ;
        RECT 109.415 194.425 109.685 194.885 ;
        RECT 111.165 194.350 111.675 194.885 ;
        RECT 113.635 194.485 113.965 194.885 ;
        RECT 114.565 194.160 114.855 194.885 ;
        RECT 115.085 194.065 115.295 194.885 ;
        RECT 115.965 194.065 116.195 194.885 ;
        RECT 117.325 194.115 120.835 194.885 ;
        RECT 121.010 194.340 126.355 194.885 ;
        RECT 119.185 193.595 120.835 194.115 ;
        RECT 124.430 193.510 124.770 194.340 ;
        RECT 126.525 194.135 127.735 194.885 ;
        RECT 127.215 193.595 127.735 194.135 ;
        RECT 14.745 190.365 15.265 190.905 ;
        RECT 17.505 190.385 18.715 190.905 ;
        RECT 14.745 189.615 15.955 190.365 ;
        RECT 16.125 189.615 18.715 190.385 ;
        RECT 22.310 190.160 22.650 190.990 ;
        RECT 25.785 190.385 26.535 190.905 ;
        RECT 18.890 189.615 24.235 190.160 ;
        RECT 24.405 189.615 24.695 190.340 ;
        RECT 24.865 189.615 26.535 190.385 ;
        RECT 30.130 190.160 30.470 190.990 ;
        RECT 35.650 190.160 35.990 190.990 ;
        RECT 48.785 190.385 49.995 190.905 ;
        RECT 60.745 190.385 61.955 190.905 ;
        RECT 26.710 189.615 32.055 190.160 ;
        RECT 32.230 189.615 37.575 190.160 ;
        RECT 38.175 189.615 38.480 190.075 ;
        RECT 39.965 189.615 40.155 190.055 ;
        RECT 42.055 189.615 42.385 190.075 ;
        RECT 44.985 189.615 45.315 189.975 ;
        RECT 46.015 189.615 46.345 189.995 ;
        RECT 47.405 189.615 49.995 190.385 ;
        RECT 50.165 189.615 50.455 190.340 ;
        RECT 51.985 189.615 52.315 189.995 ;
        RECT 53.665 189.615 54.175 190.150 ;
        RECT 56.135 189.615 56.465 190.015 ;
        RECT 58.425 189.615 58.755 189.995 ;
        RECT 59.365 189.615 61.955 190.385 ;
        RECT 62.555 189.615 62.885 189.995 ;
        RECT 63.585 189.615 63.915 189.975 ;
        RECT 66.515 189.615 66.845 190.075 ;
        RECT 68.745 189.615 68.935 190.055 ;
        RECT 70.420 189.615 70.725 190.075 ;
        RECT 72.215 189.615 72.565 190.005 ;
        RECT 73.235 189.615 73.405 190.435 ;
        RECT 75.235 190.365 75.755 190.905 ;
        RECT 79.605 190.385 80.355 190.905 ;
        RECT 74.545 189.615 75.755 190.365 ;
        RECT 75.925 189.615 76.215 190.340 ;
        RECT 78.175 189.615 78.510 190.355 ;
        RECT 78.685 189.615 80.355 190.385 ;
        RECT 83.950 190.160 84.290 190.990 ;
        RECT 96.625 190.385 97.375 190.905 ;
        RECT 105.365 190.385 106.115 190.905 ;
        RECT 80.530 189.615 85.875 190.160 ;
        RECT 86.855 189.615 87.140 190.075 ;
        RECT 88.270 189.615 88.930 190.095 ;
        RECT 90.540 189.615 90.860 190.075 ;
        RECT 91.600 189.615 92.010 190.055 ;
        RECT 93.835 189.615 94.165 189.995 ;
        RECT 94.775 189.615 95.105 189.995 ;
        RECT 95.705 189.615 97.375 190.385 ;
        RECT 98.285 189.615 98.795 190.150 ;
        RECT 100.755 189.615 101.085 190.015 ;
        RECT 101.685 189.615 101.975 190.340 ;
        RECT 103.045 189.615 103.375 189.995 ;
        RECT 104.445 189.615 106.115 190.385 ;
        RECT 120.315 190.365 120.835 190.905 ;
        RECT 107.025 189.615 107.535 190.150 ;
        RECT 109.495 189.615 109.825 190.015 ;
        RECT 110.855 189.615 111.160 190.075 ;
        RECT 112.645 189.615 112.835 190.055 ;
        RECT 114.735 189.615 115.065 190.075 ;
        RECT 117.665 189.615 117.995 189.975 ;
        RECT 118.695 189.615 119.025 189.995 ;
        RECT 119.625 189.615 120.835 190.365 ;
        RECT 124.430 190.160 124.770 190.990 ;
        RECT 127.215 190.365 127.735 190.905 ;
        RECT 121.010 189.615 126.355 190.160 ;
        RECT 126.525 189.615 127.735 190.365 ;
        RECT 14.660 189.445 127.820 189.615 ;
        RECT 14.745 188.695 15.955 189.445 ;
        RECT 14.745 188.155 15.265 188.695 ;
        RECT 16.125 188.675 17.795 189.445 ;
        RECT 17.970 188.900 23.315 189.445 ;
        RECT 23.490 188.900 28.835 189.445 ;
        RECT 17.045 188.155 17.795 188.675 ;
        RECT 21.390 188.070 21.730 188.900 ;
        RECT 26.910 188.070 27.250 188.900 ;
        RECT 29.065 188.625 29.275 189.445 ;
        RECT 29.945 188.625 30.175 189.445 ;
        RECT 30.845 188.675 34.355 189.445 ;
        RECT 32.705 188.155 34.355 188.675 ;
        RECT 34.565 188.625 34.795 189.445 ;
        RECT 35.465 188.625 35.675 189.445 ;
        RECT 36.345 189.065 36.675 189.445 ;
        RECT 37.285 188.720 37.575 189.445 ;
        RECT 38.175 189.065 38.505 189.445 ;
        RECT 39.115 189.065 39.445 189.445 ;
        RECT 41.270 189.005 41.680 189.445 ;
        RECT 42.420 188.985 42.740 189.445 ;
        RECT 44.350 188.965 45.010 189.445 ;
        RECT 46.140 188.985 46.425 189.445 ;
        RECT 48.145 188.910 48.655 189.445 ;
        RECT 50.615 189.045 50.945 189.445 ;
        RECT 52.115 188.985 52.385 189.445 ;
        RECT 54.175 188.985 54.500 189.445 ;
        RECT 55.685 188.675 57.355 189.445 ;
        RECT 57.530 188.900 62.875 189.445 ;
        RECT 56.605 188.155 57.355 188.675 ;
        RECT 60.950 188.070 61.290 188.900 ;
        RECT 63.045 188.720 63.335 189.445 ;
        RECT 63.505 188.695 64.715 189.445 ;
        RECT 64.195 188.155 64.715 188.695 ;
        RECT 64.885 188.675 68.395 189.445 ;
        RECT 69.135 188.985 69.405 189.445 ;
        RECT 71.195 188.985 71.520 189.445 ;
        RECT 72.245 188.695 73.455 189.445 ;
        RECT 73.630 188.900 78.975 189.445 ;
        RECT 79.955 188.985 80.240 189.445 ;
        RECT 81.370 188.965 82.030 189.445 ;
        RECT 83.640 188.985 83.960 189.445 ;
        RECT 84.700 189.005 85.110 189.445 ;
        RECT 86.935 189.065 87.265 189.445 ;
        RECT 87.875 189.065 88.205 189.445 ;
        RECT 66.745 188.155 68.395 188.675 ;
        RECT 72.935 188.155 73.455 188.695 ;
        RECT 77.050 188.070 77.390 188.900 ;
        RECT 88.805 188.720 89.095 189.445 ;
        RECT 89.325 188.625 89.535 189.445 ;
        RECT 90.205 188.625 90.435 189.445 ;
        RECT 91.085 189.065 91.415 189.445 ;
        RECT 92.025 188.675 94.615 189.445 ;
        RECT 95.355 188.985 95.625 189.445 ;
        RECT 97.415 188.985 97.740 189.445 ;
        RECT 98.895 188.985 99.200 189.445 ;
        RECT 100.685 189.005 100.875 189.445 ;
        RECT 102.775 188.985 103.105 189.445 ;
        RECT 105.705 189.085 106.035 189.445 ;
        RECT 106.735 189.065 107.065 189.445 ;
        RECT 107.670 188.900 113.015 189.445 ;
        RECT 113.625 189.065 113.955 189.445 ;
        RECT 93.405 188.155 94.615 188.675 ;
        RECT 111.090 188.070 111.430 188.900 ;
        RECT 114.565 188.720 114.855 189.445 ;
        RECT 116.385 189.065 116.715 189.445 ;
        RECT 117.325 188.675 120.835 189.445 ;
        RECT 121.010 188.900 126.355 189.445 ;
        RECT 119.185 188.155 120.835 188.675 ;
        RECT 124.430 188.070 124.770 188.900 ;
        RECT 126.525 188.695 127.735 189.445 ;
        RECT 127.215 188.155 127.735 188.695 ;
        RECT 14.745 184.925 15.265 185.465 ;
        RECT 17.505 184.945 18.715 185.465 ;
        RECT 14.745 184.175 15.955 184.925 ;
        RECT 16.125 184.175 18.715 184.945 ;
        RECT 22.310 184.720 22.650 185.550 ;
        RECT 36.365 184.945 37.575 185.465 ;
        RECT 18.890 184.175 24.235 184.720 ;
        RECT 24.405 184.175 24.695 184.900 ;
        RECT 26.215 184.175 26.545 184.555 ;
        RECT 27.245 184.175 27.575 184.535 ;
        RECT 30.175 184.175 30.505 184.635 ;
        RECT 32.405 184.175 32.595 184.615 ;
        RECT 34.080 184.175 34.385 184.635 ;
        RECT 34.985 184.175 37.575 184.945 ;
        RECT 37.785 184.175 38.015 184.995 ;
        RECT 38.685 184.175 38.895 184.995 ;
        RECT 39.555 184.175 39.885 184.575 ;
        RECT 41.845 184.175 42.355 184.710 ;
        RECT 44.615 184.175 44.945 184.575 ;
        RECT 46.905 184.175 47.415 184.710 ;
        RECT 48.845 184.175 49.055 184.995 ;
        RECT 49.725 184.175 49.955 184.995 ;
        RECT 60.515 184.925 61.035 185.465 ;
        RECT 63.065 184.945 64.715 185.465 ;
        RECT 50.165 184.175 50.455 184.900 ;
        RECT 51.055 184.175 51.360 184.635 ;
        RECT 52.845 184.175 53.035 184.615 ;
        RECT 54.935 184.175 55.265 184.635 ;
        RECT 57.865 184.175 58.195 184.535 ;
        RECT 58.895 184.175 59.225 184.555 ;
        RECT 59.825 184.175 61.035 184.925 ;
        RECT 61.205 184.175 64.715 184.945 ;
        RECT 68.310 184.720 68.650 185.550 ;
        RECT 73.830 184.720 74.170 185.550 ;
        RECT 78.225 184.945 79.435 185.465 ;
        RECT 84.205 184.945 84.955 185.465 ;
        RECT 64.890 184.175 70.235 184.720 ;
        RECT 70.410 184.175 75.755 184.720 ;
        RECT 75.925 184.175 76.215 184.900 ;
        RECT 76.845 184.175 79.435 184.945 ;
        RECT 80.175 184.175 80.445 184.635 ;
        RECT 82.235 184.175 82.560 184.635 ;
        RECT 83.285 184.175 84.955 184.945 ;
        RECT 85.865 184.175 86.375 184.710 ;
        RECT 88.335 184.175 88.665 184.575 ;
        RECT 89.325 184.175 89.535 184.995 ;
        RECT 90.205 184.175 90.435 184.995 ;
        RECT 91.565 184.945 92.315 185.465 ;
        RECT 90.645 184.175 92.315 184.945 ;
        RECT 93.055 184.175 93.325 184.635 ;
        RECT 95.115 184.175 95.440 184.635 ;
        RECT 96.905 184.175 97.415 184.710 ;
        RECT 99.375 184.175 99.705 184.575 ;
        RECT 100.745 184.175 101.075 184.555 ;
        RECT 101.685 184.175 101.975 184.900 ;
        RECT 102.205 184.175 102.415 184.995 ;
        RECT 103.085 184.175 103.315 184.995 ;
        RECT 105.845 184.945 107.495 185.465 ;
        RECT 113.665 184.945 115.315 185.465 ;
        RECT 103.985 184.175 107.495 184.945 ;
        RECT 108.235 184.175 108.505 184.635 ;
        RECT 110.295 184.175 110.620 184.635 ;
        RECT 111.805 184.175 115.315 184.945 ;
        RECT 118.910 184.720 119.250 185.550 ;
        RECT 124.430 184.720 124.770 185.550 ;
        RECT 127.215 184.925 127.735 185.465 ;
        RECT 115.490 184.175 120.835 184.720 ;
        RECT 121.010 184.175 126.355 184.720 ;
        RECT 126.525 184.175 127.735 184.925 ;
        RECT 14.660 184.005 127.820 184.175 ;
        RECT 14.745 183.255 15.955 184.005 ;
        RECT 16.590 183.460 21.935 184.005 ;
        RECT 22.545 183.625 22.875 184.005 ;
        RECT 24.040 183.545 24.365 184.005 ;
        RECT 26.155 183.545 26.425 184.005 ;
        RECT 27.735 183.545 28.005 184.005 ;
        RECT 29.795 183.545 30.120 184.005 ;
        RECT 31.275 183.605 31.605 184.005 ;
        RECT 33.565 183.470 34.075 184.005 ;
        RECT 14.745 182.715 15.265 183.255 ;
        RECT 20.010 182.630 20.350 183.460 ;
        RECT 35.445 183.235 37.115 184.005 ;
        RECT 37.285 183.280 37.575 184.005 ;
        RECT 38.315 183.545 38.585 184.005 ;
        RECT 40.375 183.545 40.700 184.005 ;
        RECT 42.325 183.625 42.655 184.005 ;
        RECT 43.835 183.545 44.105 184.005 ;
        RECT 45.895 183.545 46.220 184.005 ;
        RECT 47.515 183.545 47.785 184.005 ;
        RECT 49.575 183.545 49.900 184.005 ;
        RECT 51.055 183.605 51.385 184.005 ;
        RECT 53.345 183.470 53.855 184.005 ;
        RECT 36.365 182.715 37.115 183.235 ;
        RECT 55.265 183.185 55.495 184.005 ;
        RECT 56.165 183.185 56.375 184.005 ;
        RECT 57.175 183.545 57.445 184.005 ;
        RECT 59.235 183.545 59.560 184.005 ;
        RECT 60.725 183.625 61.055 184.005 ;
        RECT 62.105 183.625 62.435 184.005 ;
        RECT 63.045 183.280 63.335 184.005 ;
        RECT 63.965 183.235 66.555 184.005 ;
        RECT 66.730 183.460 72.075 184.005 ;
        RECT 72.515 183.610 72.845 184.005 ;
        RECT 73.385 183.605 73.715 184.005 ;
        RECT 65.345 182.715 66.555 183.235 ;
        RECT 70.150 182.630 70.490 183.460 ;
        RECT 74.255 183.265 74.585 184.005 ;
        RECT 77.760 183.545 77.985 184.005 ;
        RECT 78.675 183.205 78.925 184.005 ;
        RECT 80.035 183.545 80.340 184.005 ;
        RECT 81.825 183.565 82.015 184.005 ;
        RECT 83.915 183.545 84.245 184.005 ;
        RECT 86.845 183.645 87.175 184.005 ;
        RECT 87.875 183.625 88.205 184.005 ;
        RECT 88.805 183.280 89.095 184.005 ;
        RECT 90.625 183.625 90.955 184.005 ;
        RECT 92.915 183.545 93.220 184.005 ;
        RECT 94.705 183.565 94.895 184.005 ;
        RECT 96.795 183.545 97.125 184.005 ;
        RECT 99.725 183.645 100.055 184.005 ;
        RECT 100.755 183.625 101.085 184.005 ;
        RECT 103.035 183.605 103.365 184.005 ;
        RECT 105.325 183.470 105.835 184.005 ;
        RECT 107.300 183.545 107.625 184.005 ;
        RECT 109.415 183.545 109.685 184.005 ;
        RECT 111.165 183.470 111.675 184.005 ;
        RECT 113.635 183.605 113.965 184.005 ;
        RECT 114.565 183.280 114.855 184.005 ;
        RECT 115.915 183.545 116.220 184.005 ;
        RECT 117.705 183.565 117.895 184.005 ;
        RECT 119.795 183.545 120.125 184.005 ;
        RECT 122.725 183.645 123.055 184.005 ;
        RECT 123.755 183.625 124.085 184.005 ;
        RECT 124.685 183.235 126.355 184.005 ;
        RECT 126.525 183.255 127.735 184.005 ;
        RECT 125.605 182.715 126.355 183.235 ;
        RECT 127.215 182.715 127.735 183.255 ;
        RECT 14.745 179.485 15.265 180.025 ;
        RECT 17.505 179.505 18.715 180.025 ;
        RECT 14.745 178.735 15.955 179.485 ;
        RECT 16.125 178.735 18.715 179.505 ;
        RECT 22.310 179.280 22.650 180.110 ;
        RECT 18.890 178.735 24.235 179.280 ;
        RECT 24.405 178.735 24.695 179.460 ;
        RECT 44.390 179.280 44.730 180.110 ;
        RECT 25.295 178.735 25.625 179.115 ;
        RECT 26.325 178.735 26.655 179.095 ;
        RECT 29.255 178.735 29.585 179.195 ;
        RECT 31.485 178.735 31.675 179.175 ;
        RECT 33.160 178.735 33.465 179.195 ;
        RECT 35.095 178.735 35.365 179.195 ;
        RECT 37.155 178.735 37.480 179.195 ;
        RECT 39.105 178.735 39.435 179.115 ;
        RECT 40.970 178.735 46.315 179.280 ;
        RECT 47.055 178.735 47.325 179.195 ;
        RECT 49.115 178.735 49.440 179.195 ;
        RECT 50.165 178.735 50.455 179.460 ;
        RECT 52.115 178.735 52.385 179.195 ;
        RECT 54.175 178.735 54.500 179.195 ;
        RECT 55.655 178.735 55.960 179.195 ;
        RECT 57.445 178.735 57.635 179.175 ;
        RECT 59.535 178.735 59.865 179.195 ;
        RECT 62.465 178.735 62.795 179.095 ;
        RECT 63.495 178.735 63.825 179.115 ;
        RECT 64.945 178.735 65.155 179.555 ;
        RECT 65.825 178.735 66.055 179.555 ;
        RECT 66.270 178.735 66.530 179.575 ;
        RECT 93.635 179.485 94.155 180.025 ;
        RECT 67.130 178.735 67.460 179.115 ;
        RECT 68.375 178.735 68.705 179.130 ;
        RECT 69.245 178.735 69.575 179.135 ;
        RECT 70.115 178.735 70.445 179.475 ;
        RECT 71.755 178.735 72.085 179.115 ;
        RECT 74.855 178.735 75.185 179.115 ;
        RECT 75.925 178.735 76.215 179.460 ;
        RECT 76.655 178.735 76.985 179.130 ;
        RECT 77.525 178.735 77.855 179.135 ;
        RECT 78.395 178.735 78.725 179.475 ;
        RECT 80.345 178.735 80.855 179.270 ;
        RECT 82.815 178.735 83.145 179.135 ;
        RECT 83.745 178.735 84.050 179.245 ;
        RECT 84.650 178.735 84.910 179.260 ;
        RECT 85.510 178.735 85.770 179.295 ;
        RECT 86.370 178.735 86.630 179.215 ;
        RECT 87.230 178.735 87.490 179.215 ;
        RECT 88.090 178.735 88.335 179.215 ;
        RECT 88.950 178.735 89.195 179.215 ;
        RECT 89.805 178.735 90.055 179.215 ;
        RECT 90.665 178.735 90.915 179.215 ;
        RECT 91.525 178.735 91.785 179.215 ;
        RECT 92.385 178.735 92.685 179.215 ;
        RECT 92.945 178.735 94.155 179.485 ;
        RECT 94.895 178.735 95.165 179.195 ;
        RECT 96.955 178.735 97.280 179.195 ;
        RECT 98.575 178.735 98.845 179.195 ;
        RECT 100.635 178.735 100.960 179.195 ;
        RECT 101.685 178.735 101.975 179.460 ;
        RECT 102.585 178.735 102.915 179.115 ;
        RECT 104.495 178.735 104.745 179.535 ;
        RECT 125.145 179.505 126.355 180.025 ;
        RECT 105.435 178.735 105.660 179.195 ;
        RECT 108.405 178.735 108.915 179.270 ;
        RECT 110.875 178.735 111.205 179.135 ;
        RECT 112.235 178.735 112.540 179.195 ;
        RECT 114.025 178.735 114.215 179.175 ;
        RECT 116.115 178.735 116.445 179.195 ;
        RECT 119.045 178.735 119.375 179.095 ;
        RECT 120.075 178.735 120.405 179.115 ;
        RECT 121.445 178.735 121.775 179.115 ;
        RECT 122.825 178.735 123.155 179.115 ;
        RECT 123.765 178.735 126.355 179.505 ;
        RECT 127.215 179.485 127.735 180.025 ;
        RECT 126.525 178.735 127.735 179.485 ;
        RECT 14.660 178.565 127.820 178.735 ;
        RECT 14.745 177.815 15.955 178.565 ;
        RECT 14.745 177.275 15.265 177.815 ;
        RECT 16.125 177.795 19.635 178.565 ;
        RECT 19.810 178.020 25.155 178.565 ;
        RECT 17.985 177.275 19.635 177.795 ;
        RECT 23.230 177.190 23.570 178.020 ;
        RECT 25.385 177.745 25.595 178.565 ;
        RECT 26.265 177.745 26.495 178.565 ;
        RECT 27.145 178.185 27.475 178.565 ;
        RECT 28.515 178.105 28.820 178.565 ;
        RECT 30.305 178.125 30.495 178.565 ;
        RECT 32.395 178.105 32.725 178.565 ;
        RECT 35.325 178.205 35.655 178.565 ;
        RECT 36.355 178.185 36.685 178.565 ;
        RECT 37.285 177.840 37.575 178.565 ;
        RECT 38.175 178.165 38.505 178.565 ;
        RECT 40.465 178.030 40.975 178.565 ;
        RECT 41.885 177.795 43.555 178.565 ;
        RECT 45.560 178.105 45.785 178.565 ;
        RECT 42.805 177.275 43.555 177.795 ;
        RECT 46.475 177.765 46.725 178.565 ;
        RECT 48.375 177.765 48.625 178.565 ;
        RECT 49.315 178.105 49.540 178.565 ;
        RECT 52.055 177.765 52.305 178.565 ;
        RECT 52.995 178.105 53.220 178.565 ;
        RECT 56.425 178.030 56.935 178.565 ;
        RECT 58.895 178.165 59.225 178.565 ;
        RECT 60.345 178.085 60.625 178.565 ;
        RECT 61.230 178.085 61.485 178.565 ;
        RECT 62.130 178.085 62.405 178.565 ;
        RECT 63.045 177.840 63.335 178.565 ;
        RECT 63.970 177.725 64.230 178.565 ;
        RECT 64.830 178.185 65.160 178.565 ;
        RECT 65.810 177.725 66.070 178.565 ;
        RECT 66.670 178.185 67.000 178.565 ;
        RECT 68.615 178.205 68.945 178.565 ;
        RECT 71.135 178.170 71.465 178.565 ;
        RECT 72.005 178.165 72.335 178.565 ;
        RECT 72.875 177.825 73.205 178.565 ;
        RECT 75.920 178.105 76.145 178.565 ;
        RECT 76.835 177.765 77.085 178.565 ;
        RECT 77.875 178.085 78.045 178.565 ;
        RECT 78.715 178.085 78.885 178.565 ;
        RECT 79.555 178.085 79.725 178.565 ;
        RECT 80.395 178.085 80.565 178.565 ;
        RECT 81.235 178.085 81.405 178.565 ;
        RECT 82.075 178.085 82.245 178.565 ;
        RECT 82.915 178.085 83.085 178.565 ;
        RECT 83.755 178.085 83.925 178.565 ;
        RECT 84.595 178.085 84.765 178.565 ;
        RECT 85.435 178.085 85.605 178.565 ;
        RECT 86.275 178.085 86.445 178.565 ;
        RECT 87.115 178.085 87.285 178.565 ;
        RECT 87.955 178.085 88.125 178.565 ;
        RECT 88.805 177.840 89.095 178.565 ;
        RECT 90.190 178.020 95.535 178.565 ;
        RECT 93.610 177.190 93.950 178.020 ;
        RECT 95.765 177.745 95.975 178.565 ;
        RECT 96.645 177.745 96.875 178.565 ;
        RECT 97.085 177.795 98.755 178.565 ;
        RECT 98.005 177.275 98.755 177.795 ;
        RECT 99.435 177.765 99.685 178.565 ;
        RECT 100.375 178.105 100.600 178.565 ;
        RECT 102.605 177.795 105.195 178.565 ;
        RECT 103.985 177.275 105.195 177.795 ;
        RECT 105.875 177.765 106.125 178.565 ;
        RECT 106.815 178.105 107.040 178.565 ;
        RECT 109.600 178.105 109.925 178.565 ;
        RECT 111.715 178.105 111.985 178.565 ;
        RECT 113.225 177.745 113.455 178.565 ;
        RECT 114.125 177.745 114.335 178.565 ;
        RECT 114.565 177.840 114.855 178.565 ;
        RECT 115.025 177.795 116.695 178.565 ;
        RECT 115.945 177.275 116.695 177.795 ;
        RECT 116.905 177.745 117.135 178.565 ;
        RECT 117.805 177.745 118.015 178.565 ;
        RECT 118.245 177.795 120.835 178.565 ;
        RECT 121.010 178.020 126.355 178.565 ;
        RECT 119.625 177.275 120.835 177.795 ;
        RECT 124.430 177.190 124.770 178.020 ;
        RECT 126.525 177.815 127.735 178.565 ;
        RECT 127.215 177.275 127.735 177.815 ;
        RECT 14.745 174.045 15.265 174.585 ;
        RECT 17.505 174.065 18.715 174.585 ;
        RECT 14.745 173.295 15.955 174.045 ;
        RECT 16.125 173.295 18.715 174.065 ;
        RECT 22.310 173.840 22.650 174.670 ;
        RECT 18.890 173.295 24.235 173.840 ;
        RECT 24.405 173.295 24.695 174.020 ;
        RECT 25.845 173.295 26.055 174.115 ;
        RECT 26.725 173.295 26.955 174.115 ;
        RECT 27.735 173.295 28.005 173.755 ;
        RECT 29.795 173.295 30.120 173.755 ;
        RECT 31.735 173.295 32.065 173.695 ;
        RECT 34.025 173.295 34.535 173.830 ;
        RECT 37.280 173.295 37.505 173.755 ;
        RECT 38.195 173.295 38.445 174.095 ;
        RECT 39.635 173.295 39.885 174.095 ;
        RECT 40.575 173.295 40.800 173.755 ;
        RECT 44.640 173.295 44.865 173.755 ;
        RECT 45.555 173.295 45.805 174.095 ;
        RECT 46.995 173.295 47.245 174.095 ;
        RECT 51.315 174.045 51.835 174.585 ;
        RECT 61.665 174.065 62.415 174.585 ;
        RECT 66.285 174.065 67.935 174.585 ;
        RECT 47.935 173.295 48.160 173.755 ;
        RECT 50.165 173.295 50.455 174.020 ;
        RECT 50.625 173.295 51.835 174.045 ;
        RECT 52.575 173.295 52.845 173.755 ;
        RECT 54.635 173.295 54.960 173.755 ;
        RECT 57.345 173.295 57.855 173.830 ;
        RECT 59.815 173.295 60.145 173.695 ;
        RECT 60.745 173.295 62.415 174.065 ;
        RECT 63.025 173.295 63.355 173.675 ;
        RECT 64.425 173.295 67.935 174.065 ;
        RECT 68.545 173.295 68.785 173.775 ;
        RECT 69.375 173.295 69.705 173.775 ;
        RECT 70.215 173.295 70.545 174.095 ;
        RECT 71.330 173.295 71.590 174.135 ;
        RECT 72.190 173.295 72.520 173.675 ;
        RECT 73.640 173.295 73.970 173.675 ;
        RECT 74.570 173.295 74.830 174.135 ;
        RECT 75.925 173.295 76.215 174.020 ;
        RECT 79.140 173.295 79.365 173.755 ;
        RECT 80.055 173.295 80.305 174.095 ;
        RECT 81.495 173.295 81.745 174.095 ;
        RECT 91.795 174.045 92.315 174.585 ;
        RECT 94.345 174.065 95.995 174.585 ;
        RECT 82.435 173.295 82.660 173.755 ;
        RECT 85.220 173.295 85.545 173.755 ;
        RECT 87.335 173.295 87.605 173.755 ;
        RECT 88.815 173.295 89.090 173.775 ;
        RECT 89.735 173.295 89.990 173.775 ;
        RECT 90.595 173.295 90.875 173.775 ;
        RECT 91.105 173.295 92.315 174.045 ;
        RECT 92.485 173.295 95.995 174.065 ;
        RECT 99.590 173.840 99.930 174.670 ;
        RECT 96.170 173.295 101.515 173.840 ;
        RECT 101.685 173.295 101.975 174.020 ;
        RECT 102.145 173.295 102.450 173.805 ;
        RECT 103.050 173.295 103.310 173.820 ;
        RECT 103.910 173.295 104.170 173.855 ;
        RECT 104.770 173.295 105.030 173.775 ;
        RECT 105.630 173.295 105.890 173.775 ;
        RECT 106.490 173.295 106.735 173.775 ;
        RECT 107.350 173.295 107.595 173.775 ;
        RECT 108.205 173.295 108.455 173.775 ;
        RECT 109.065 173.295 109.315 173.775 ;
        RECT 109.925 173.295 110.185 173.775 ;
        RECT 110.785 173.295 111.085 173.775 ;
        RECT 111.855 173.295 112.105 174.095 ;
        RECT 112.795 173.295 113.020 173.755 ;
        RECT 116.860 173.295 117.085 173.755 ;
        RECT 117.775 173.295 118.025 174.095 ;
        RECT 118.765 173.295 118.975 174.115 ;
        RECT 119.645 173.295 119.875 174.115 ;
        RECT 124.430 173.840 124.770 174.670 ;
        RECT 127.215 174.045 127.735 174.585 ;
        RECT 121.010 173.295 126.355 173.840 ;
        RECT 126.525 173.295 127.735 174.045 ;
        RECT 14.660 173.125 127.820 173.295 ;
        RECT 14.745 172.375 15.955 173.125 ;
        RECT 17.050 172.580 22.395 173.125 ;
        RECT 22.570 172.580 27.915 173.125 ;
        RECT 28.090 172.580 33.435 173.125 ;
        RECT 35.440 172.665 35.665 173.125 ;
        RECT 14.745 171.835 15.265 172.375 ;
        RECT 20.470 171.750 20.810 172.580 ;
        RECT 25.990 171.750 26.330 172.580 ;
        RECT 31.510 171.750 31.850 172.580 ;
        RECT 36.355 172.325 36.605 173.125 ;
        RECT 37.285 172.400 37.575 173.125 ;
        RECT 38.715 172.325 38.965 173.125 ;
        RECT 39.655 172.665 39.880 173.125 ;
        RECT 41.885 172.355 44.475 173.125 ;
        RECT 44.735 172.645 45.035 173.125 ;
        RECT 45.635 172.645 45.895 173.125 ;
        RECT 46.505 172.645 46.755 173.125 ;
        RECT 47.365 172.645 47.615 173.125 ;
        RECT 48.225 172.645 48.470 173.125 ;
        RECT 49.085 172.645 49.330 173.125 ;
        RECT 49.930 172.645 50.190 173.125 ;
        RECT 50.790 172.645 51.050 173.125 ;
        RECT 51.650 172.565 51.910 173.125 ;
        RECT 52.510 172.600 52.770 173.125 ;
        RECT 53.370 172.615 53.675 173.125 ;
        RECT 54.275 172.665 54.580 173.125 ;
        RECT 56.065 172.685 56.255 173.125 ;
        RECT 58.155 172.665 58.485 173.125 ;
        RECT 61.085 172.765 61.415 173.125 ;
        RECT 62.115 172.745 62.445 173.125 ;
        RECT 63.045 172.400 63.335 173.125 ;
        RECT 43.265 171.835 44.475 172.355 ;
        RECT 63.565 172.305 63.775 173.125 ;
        RECT 64.445 172.305 64.675 173.125 ;
        RECT 65.810 172.580 71.155 173.125 ;
        RECT 71.330 172.580 76.675 173.125 ;
        RECT 76.850 172.580 82.195 173.125 ;
        RECT 82.805 172.645 83.045 173.125 ;
        RECT 83.635 172.645 83.965 173.125 ;
        RECT 69.230 171.750 69.570 172.580 ;
        RECT 74.750 171.750 75.090 172.580 ;
        RECT 80.270 171.750 80.610 172.580 ;
        RECT 84.475 172.325 84.805 173.125 ;
        RECT 85.695 172.665 85.965 173.125 ;
        RECT 87.755 172.665 88.080 173.125 ;
        RECT 88.805 172.400 89.095 173.125 ;
        RECT 89.765 172.305 89.995 173.125 ;
        RECT 90.665 172.305 90.875 173.125 ;
        RECT 91.535 172.665 91.840 173.125 ;
        RECT 93.325 172.685 93.515 173.125 ;
        RECT 95.415 172.665 95.745 173.125 ;
        RECT 98.345 172.765 98.675 173.125 ;
        RECT 99.375 172.745 99.705 173.125 ;
        RECT 101.225 172.355 104.735 173.125 ;
        RECT 105.425 172.655 105.725 173.125 ;
        RECT 106.320 172.655 106.580 173.125 ;
        RECT 107.180 172.655 107.475 173.125 ;
        RECT 103.085 171.835 104.735 172.355 ;
        RECT 108.635 172.325 108.885 173.125 ;
        RECT 109.575 172.665 109.800 173.125 ;
        RECT 111.805 172.375 113.015 173.125 ;
        RECT 112.495 171.835 113.015 172.375 ;
        RECT 113.225 172.305 113.455 173.125 ;
        RECT 114.125 172.305 114.335 173.125 ;
        RECT 114.565 172.400 114.855 173.125 ;
        RECT 116.375 172.665 116.680 173.125 ;
        RECT 118.165 172.685 118.355 173.125 ;
        RECT 120.255 172.665 120.585 173.125 ;
        RECT 123.185 172.765 123.515 173.125 ;
        RECT 124.215 172.745 124.545 173.125 ;
        RECT 125.145 172.375 126.355 173.125 ;
        RECT 126.525 172.375 127.735 173.125 ;
        RECT 125.835 171.835 126.355 172.375 ;
        RECT 127.215 171.835 127.735 172.375 ;
        RECT 14.745 168.605 15.265 169.145 ;
        RECT 17.505 168.625 18.715 169.145 ;
        RECT 14.745 167.855 15.955 168.605 ;
        RECT 16.125 167.855 18.715 168.625 ;
        RECT 22.310 168.400 22.650 169.230 ;
        RECT 26.245 168.625 26.995 169.145 ;
        RECT 18.890 167.855 24.235 168.400 ;
        RECT 24.405 167.855 24.695 168.580 ;
        RECT 25.325 167.855 26.995 168.625 ;
        RECT 27.225 167.855 27.435 168.675 ;
        RECT 28.105 167.855 28.335 168.675 ;
        RECT 29.465 168.625 30.215 169.145 ;
        RECT 28.545 167.855 30.215 168.625 ;
        RECT 30.445 167.855 30.655 168.675 ;
        RECT 31.325 167.855 31.555 168.675 ;
        RECT 39.125 168.625 39.875 169.145 ;
        RECT 32.335 167.855 32.605 168.315 ;
        RECT 34.395 167.855 34.720 168.315 ;
        RECT 36.115 167.855 36.445 168.545 ;
        RECT 37.695 167.855 38.025 168.345 ;
        RECT 38.205 167.855 39.875 168.625 ;
        RECT 43.470 168.400 43.810 169.230 ;
        RECT 40.050 167.855 45.395 168.400 ;
        RECT 46.075 167.855 46.325 168.655 ;
        RECT 51.545 168.625 52.295 169.145 ;
        RECT 56.605 168.625 57.355 169.145 ;
        RECT 47.015 167.855 47.240 168.315 ;
        RECT 50.165 167.855 50.455 168.580 ;
        RECT 50.625 167.855 52.295 168.625 ;
        RECT 52.985 167.855 53.285 168.325 ;
        RECT 53.880 167.855 54.140 168.325 ;
        RECT 54.740 167.855 55.035 168.325 ;
        RECT 55.685 167.855 57.355 168.625 ;
        RECT 60.950 168.400 61.290 169.230 ;
        RECT 66.470 168.400 66.810 169.230 ;
        RECT 57.530 167.855 62.875 168.400 ;
        RECT 63.050 167.855 68.395 168.400 ;
        RECT 69.040 167.855 69.370 168.235 ;
        RECT 69.970 167.855 70.230 168.695 ;
        RECT 70.410 167.855 70.670 168.695 ;
        RECT 99.865 168.625 101.515 169.145 ;
        RECT 71.270 167.855 71.600 168.235 ;
        RECT 73.175 167.855 73.450 168.335 ;
        RECT 74.095 167.855 74.350 168.335 ;
        RECT 74.955 167.855 75.235 168.335 ;
        RECT 75.925 167.855 76.215 168.580 ;
        RECT 77.125 167.855 77.635 168.390 ;
        RECT 79.595 167.855 79.925 168.255 ;
        RECT 81.335 167.855 81.620 168.315 ;
        RECT 82.750 167.855 83.410 168.335 ;
        RECT 85.020 167.855 85.340 168.315 ;
        RECT 86.080 167.855 86.490 168.295 ;
        RECT 88.315 167.855 88.645 168.235 ;
        RECT 89.255 167.855 89.585 168.235 ;
        RECT 91.845 167.855 92.355 168.390 ;
        RECT 94.315 167.855 94.645 168.255 ;
        RECT 96.605 167.855 96.935 168.235 ;
        RECT 98.005 167.855 101.515 168.625 ;
        RECT 101.685 167.855 101.975 168.580 ;
        RECT 103.035 167.855 103.340 168.315 ;
        RECT 104.825 167.855 105.015 168.295 ;
        RECT 106.915 167.855 107.245 168.315 ;
        RECT 109.845 167.855 110.175 168.215 ;
        RECT 110.875 167.855 111.205 168.235 ;
        RECT 113.155 167.855 113.485 168.255 ;
        RECT 115.445 167.855 115.955 168.390 ;
        RECT 117.420 167.855 117.745 168.315 ;
        RECT 119.535 167.855 119.805 168.315 ;
        RECT 120.585 167.855 120.815 168.675 ;
        RECT 121.485 167.855 121.695 168.675 ;
        RECT 125.835 168.605 126.355 169.145 ;
        RECT 127.215 168.605 127.735 169.145 ;
        RECT 121.930 167.855 122.265 168.255 ;
        RECT 122.850 167.855 123.125 168.335 ;
        RECT 124.205 167.855 124.535 168.235 ;
        RECT 125.145 167.855 126.355 168.605 ;
        RECT 126.525 167.855 127.735 168.605 ;
        RECT 14.660 167.685 127.820 167.855 ;
        RECT 14.745 166.935 15.955 167.685 ;
        RECT 14.745 166.395 15.265 166.935 ;
        RECT 16.585 166.915 18.255 167.685 ;
        RECT 18.855 167.225 19.160 167.685 ;
        RECT 20.645 167.245 20.835 167.685 ;
        RECT 22.735 167.225 23.065 167.685 ;
        RECT 25.665 167.325 25.995 167.685 ;
        RECT 26.695 167.305 27.025 167.685 ;
        RECT 27.715 167.205 28.015 167.685 ;
        RECT 28.615 167.205 28.875 167.685 ;
        RECT 29.485 167.205 29.735 167.685 ;
        RECT 30.345 167.205 30.595 167.685 ;
        RECT 31.205 167.205 31.450 167.685 ;
        RECT 32.065 167.205 32.310 167.685 ;
        RECT 32.910 167.205 33.170 167.685 ;
        RECT 33.770 167.205 34.030 167.685 ;
        RECT 34.630 167.125 34.890 167.685 ;
        RECT 35.490 167.160 35.750 167.685 ;
        RECT 36.350 167.175 36.655 167.685 ;
        RECT 37.285 166.960 37.575 167.685 ;
        RECT 38.185 167.305 38.515 167.685 ;
        RECT 17.505 166.395 18.255 166.915 ;
        RECT 39.185 166.865 39.395 167.685 ;
        RECT 40.065 166.865 40.295 167.685 ;
        RECT 41.405 167.305 41.735 167.685 ;
        RECT 42.385 166.865 42.615 167.685 ;
        RECT 43.285 166.865 43.495 167.685 ;
        RECT 44.295 167.225 44.565 167.685 ;
        RECT 46.355 167.225 46.680 167.685 ;
        RECT 47.835 167.225 48.140 167.685 ;
        RECT 49.625 167.245 49.815 167.685 ;
        RECT 51.715 167.225 52.045 167.685 ;
        RECT 54.645 167.325 54.975 167.685 ;
        RECT 55.675 167.305 56.005 167.685 ;
        RECT 57.585 166.865 57.795 167.685 ;
        RECT 58.465 166.865 58.695 167.685 ;
        RECT 59.975 166.885 60.305 167.685 ;
        RECT 60.815 167.205 61.145 167.685 ;
        RECT 61.735 167.205 61.975 167.685 ;
        RECT 63.045 166.960 63.335 167.685 ;
        RECT 64.575 166.885 64.905 167.685 ;
        RECT 65.415 167.205 65.745 167.685 ;
        RECT 66.335 167.205 66.575 167.685 ;
        RECT 67.245 167.205 67.525 167.685 ;
        RECT 68.130 167.205 68.385 167.685 ;
        RECT 69.030 167.205 69.305 167.685 ;
        RECT 69.945 166.935 71.155 167.685 ;
        RECT 71.835 167.325 72.165 167.685 ;
        RECT 74.085 166.935 75.295 167.685 ;
        RECT 76.275 167.225 76.560 167.685 ;
        RECT 77.690 167.205 78.350 167.685 ;
        RECT 79.960 167.225 80.280 167.685 ;
        RECT 81.020 167.245 81.430 167.685 ;
        RECT 83.255 167.305 83.585 167.685 ;
        RECT 84.195 167.305 84.525 167.685 ;
        RECT 70.635 166.395 71.155 166.935 ;
        RECT 74.775 166.395 75.295 166.935 ;
        RECT 85.185 166.865 85.395 167.685 ;
        RECT 86.065 166.865 86.295 167.685 ;
        RECT 86.565 166.865 86.775 167.685 ;
        RECT 87.445 166.865 87.675 167.685 ;
        RECT 88.805 166.960 89.095 167.685 ;
        RECT 89.725 166.915 91.395 167.685 ;
        RECT 91.570 167.140 96.915 167.685 ;
        RECT 97.895 167.225 98.180 167.685 ;
        RECT 99.310 167.205 99.970 167.685 ;
        RECT 101.580 167.225 101.900 167.685 ;
        RECT 102.640 167.245 103.050 167.685 ;
        RECT 104.875 167.305 105.205 167.685 ;
        RECT 105.815 167.305 106.145 167.685 ;
        RECT 107.775 167.225 108.045 167.685 ;
        RECT 109.835 167.225 110.160 167.685 ;
        RECT 111.440 167.225 111.765 167.685 ;
        RECT 113.555 167.225 113.825 167.685 ;
        RECT 90.645 166.395 91.395 166.915 ;
        RECT 94.990 166.310 95.330 167.140 ;
        RECT 114.565 166.960 114.855 167.685 ;
        RECT 116.375 167.225 116.680 167.685 ;
        RECT 118.165 167.245 118.355 167.685 ;
        RECT 120.255 167.225 120.585 167.685 ;
        RECT 123.185 167.325 123.515 167.685 ;
        RECT 124.215 167.305 124.545 167.685 ;
        RECT 125.145 166.935 126.355 167.685 ;
        RECT 126.525 166.935 127.735 167.685 ;
        RECT 125.835 166.395 126.355 166.935 ;
        RECT 127.215 166.395 127.735 166.935 ;
        RECT 14.745 163.165 15.265 163.705 ;
        RECT 17.505 163.185 18.715 163.705 ;
        RECT 14.745 162.415 15.955 163.165 ;
        RECT 16.125 162.415 18.715 163.185 ;
        RECT 22.310 162.960 22.650 163.790 ;
        RECT 65.805 163.185 67.015 163.705 ;
        RECT 18.890 162.415 24.235 162.960 ;
        RECT 24.405 162.415 24.695 163.140 ;
        RECT 26.225 162.415 26.555 162.795 ;
        RECT 27.595 162.415 27.900 162.875 ;
        RECT 29.385 162.415 29.575 162.855 ;
        RECT 31.475 162.415 31.805 162.875 ;
        RECT 34.405 162.415 34.735 162.775 ;
        RECT 35.435 162.415 35.765 162.795 ;
        RECT 36.795 162.415 37.100 162.875 ;
        RECT 38.585 162.415 38.775 162.855 ;
        RECT 40.675 162.415 41.005 162.875 ;
        RECT 43.605 162.415 43.935 162.775 ;
        RECT 44.635 162.415 44.965 162.795 ;
        RECT 45.995 162.415 46.325 162.815 ;
        RECT 48.285 162.415 48.795 162.950 ;
        RECT 50.165 162.415 50.455 163.140 ;
        RECT 51.365 162.415 51.875 162.950 ;
        RECT 53.835 162.415 54.165 162.815 ;
        RECT 55.195 162.415 55.500 162.875 ;
        RECT 56.985 162.415 57.175 162.855 ;
        RECT 59.075 162.415 59.405 162.875 ;
        RECT 62.005 162.415 62.335 162.775 ;
        RECT 63.035 162.415 63.365 162.795 ;
        RECT 64.425 162.415 67.015 163.185 ;
        RECT 73.830 162.960 74.170 163.790 ;
        RECT 77.305 163.185 78.055 163.705 ;
        RECT 84.665 163.185 85.415 163.705 ;
        RECT 67.245 162.415 67.525 162.895 ;
        RECT 68.130 162.415 68.385 162.895 ;
        RECT 69.030 162.415 69.305 162.895 ;
        RECT 70.410 162.415 75.755 162.960 ;
        RECT 75.925 162.415 76.215 163.140 ;
        RECT 76.385 162.415 78.055 163.185 ;
        RECT 78.965 162.415 79.475 162.950 ;
        RECT 81.435 162.415 81.765 162.815 ;
        RECT 82.805 162.415 83.135 162.795 ;
        RECT 83.745 162.415 85.415 163.185 ;
        RECT 91.310 162.960 91.650 163.790 ;
        RECT 86.025 162.415 86.355 162.795 ;
        RECT 87.890 162.415 93.235 162.960 ;
        RECT 94.145 162.415 94.655 162.950 ;
        RECT 96.615 162.415 96.945 162.815 ;
        RECT 98.285 162.415 98.795 162.950 ;
        RECT 100.755 162.415 101.085 162.815 ;
        RECT 101.685 162.415 101.975 163.140 ;
        RECT 102.700 162.415 103.025 162.875 ;
        RECT 104.815 162.415 105.085 162.875 ;
        RECT 107.175 162.415 107.505 162.815 ;
        RECT 109.465 162.415 109.975 162.950 ;
        RECT 110.945 162.415 111.155 163.235 ;
        RECT 111.825 162.415 112.055 163.235 ;
        RECT 125.145 163.185 126.355 163.705 ;
        RECT 113.615 162.415 113.920 162.875 ;
        RECT 115.405 162.415 115.595 162.855 ;
        RECT 117.495 162.415 117.825 162.875 ;
        RECT 120.425 162.415 120.755 162.775 ;
        RECT 121.455 162.415 121.785 162.795 ;
        RECT 122.825 162.415 123.155 162.795 ;
        RECT 123.765 162.415 126.355 163.185 ;
        RECT 127.215 163.165 127.735 163.705 ;
        RECT 126.525 162.415 127.735 163.165 ;
        RECT 14.660 162.245 127.820 162.415 ;
        RECT 14.745 161.495 15.955 162.245 ;
        RECT 14.745 160.955 15.265 161.495 ;
        RECT 16.125 161.475 17.795 162.245 ;
        RECT 18.775 161.785 19.060 162.245 ;
        RECT 20.190 161.765 20.850 162.245 ;
        RECT 22.460 161.785 22.780 162.245 ;
        RECT 23.520 161.805 23.930 162.245 ;
        RECT 25.755 161.865 26.085 162.245 ;
        RECT 26.695 161.865 27.025 162.245 ;
        RECT 28.055 161.845 28.385 162.245 ;
        RECT 30.345 161.710 30.855 162.245 ;
        RECT 31.765 161.495 32.975 162.245 ;
        RECT 33.885 161.710 34.395 162.245 ;
        RECT 36.355 161.845 36.685 162.245 ;
        RECT 37.285 161.520 37.575 162.245 ;
        RECT 17.045 160.955 17.795 161.475 ;
        RECT 32.455 160.955 32.975 161.495 ;
        RECT 38.205 161.475 41.715 162.245 ;
        RECT 42.440 161.785 42.765 162.245 ;
        RECT 44.555 161.785 44.825 162.245 ;
        RECT 45.565 161.495 46.775 162.245 ;
        RECT 47.515 161.785 47.785 162.245 ;
        RECT 49.575 161.785 49.900 162.245 ;
        RECT 51.365 161.710 51.875 162.245 ;
        RECT 53.835 161.845 54.165 162.245 ;
        RECT 55.335 161.785 55.605 162.245 ;
        RECT 57.395 161.785 57.720 162.245 ;
        RECT 59.345 161.865 59.675 162.245 ;
        RECT 40.065 160.955 41.715 161.475 ;
        RECT 46.255 160.955 46.775 161.495 ;
        RECT 60.285 161.475 62.875 162.245 ;
        RECT 63.045 161.520 63.335 162.245 ;
        RECT 63.505 161.495 64.715 162.245 ;
        RECT 61.665 160.955 62.875 161.475 ;
        RECT 64.195 160.955 64.715 161.495 ;
        RECT 64.890 161.405 65.150 162.245 ;
        RECT 65.750 161.865 66.080 162.245 ;
        RECT 66.730 161.405 66.990 162.245 ;
        RECT 67.590 161.865 67.920 162.245 ;
        RECT 69.040 161.865 69.370 162.245 ;
        RECT 69.970 161.405 70.230 162.245 ;
        RECT 70.880 161.865 71.210 162.245 ;
        RECT 71.810 161.405 72.070 162.245 ;
        RECT 72.245 161.475 74.835 162.245 ;
        RECT 75.010 161.700 80.355 162.245 ;
        RECT 73.625 160.955 74.835 161.475 ;
        RECT 78.430 160.870 78.770 161.700 ;
        RECT 80.585 161.425 80.795 162.245 ;
        RECT 81.465 161.425 81.695 162.245 ;
        RECT 82.645 161.710 83.155 162.245 ;
        RECT 85.115 161.845 85.445 162.245 ;
        RECT 86.945 161.865 87.275 162.245 ;
        RECT 88.805 161.520 89.095 162.245 ;
        RECT 90.075 161.785 90.360 162.245 ;
        RECT 91.490 161.765 92.150 162.245 ;
        RECT 93.760 161.785 94.080 162.245 ;
        RECT 94.820 161.805 95.230 162.245 ;
        RECT 97.055 161.865 97.385 162.245 ;
        RECT 97.995 161.865 98.325 162.245 ;
        RECT 100.285 161.865 100.615 162.245 ;
        RECT 101.285 161.425 101.495 162.245 ;
        RECT 102.165 161.425 102.395 162.245 ;
        RECT 103.160 161.785 103.485 162.245 ;
        RECT 105.275 161.785 105.545 162.245 ;
        RECT 107.315 161.785 107.585 162.245 ;
        RECT 109.375 161.785 109.700 162.245 ;
        RECT 111.165 161.710 111.675 162.245 ;
        RECT 113.635 161.845 113.965 162.245 ;
        RECT 114.565 161.520 114.855 162.245 ;
        RECT 115.765 161.710 116.275 162.245 ;
        RECT 118.235 161.845 118.565 162.245 ;
        RECT 119.735 161.785 120.005 162.245 ;
        RECT 121.795 161.785 122.120 162.245 ;
        RECT 123.285 161.865 123.615 162.245 ;
        RECT 124.685 161.475 126.355 162.245 ;
        RECT 126.525 161.495 127.735 162.245 ;
        RECT 125.605 160.955 126.355 161.475 ;
        RECT 127.215 160.955 127.735 161.495 ;
        RECT 14.745 157.725 15.265 158.265 ;
        RECT 16.815 157.725 17.335 158.265 ;
        RECT 14.745 156.975 15.955 157.725 ;
        RECT 16.125 156.975 17.335 157.725 ;
        RECT 17.565 156.975 17.775 157.795 ;
        RECT 18.445 156.975 18.675 157.795 ;
        RECT 18.925 156.975 19.155 157.795 ;
        RECT 19.825 156.975 20.035 157.795 ;
        RECT 21.005 156.975 21.515 157.510 ;
        RECT 23.475 156.975 23.805 157.375 ;
        RECT 24.405 156.975 24.695 157.700 ;
        RECT 30.130 157.520 30.470 158.350 ;
        RECT 36.595 157.725 37.115 158.265 ;
        RECT 25.305 156.975 25.635 157.355 ;
        RECT 26.710 156.975 32.055 157.520 ;
        RECT 32.780 156.975 33.105 157.435 ;
        RECT 34.895 156.975 35.165 157.435 ;
        RECT 35.905 156.975 37.115 157.725 ;
        RECT 40.710 157.520 41.050 158.350 ;
        RECT 37.290 156.975 42.635 157.520 ;
        RECT 44.640 156.975 44.865 157.435 ;
        RECT 45.555 156.975 45.805 157.775 ;
        RECT 46.995 156.975 47.245 157.775 ;
        RECT 47.935 156.975 48.160 157.435 ;
        RECT 50.165 156.975 50.455 157.700 ;
        RECT 51.135 156.975 51.385 157.775 ;
        RECT 59.570 157.520 59.910 158.350 ;
        RECT 52.075 156.975 52.300 157.435 ;
        RECT 55.205 156.975 55.535 157.355 ;
        RECT 56.150 156.975 61.495 157.520 ;
        RECT 61.815 156.975 62.145 157.775 ;
        RECT 66.745 157.745 68.395 158.265 ;
        RECT 62.655 156.975 62.985 157.455 ;
        RECT 63.575 156.975 63.815 157.455 ;
        RECT 64.885 156.975 68.395 157.745 ;
        RECT 69.040 156.975 69.370 157.355 ;
        RECT 69.970 156.975 70.230 157.815 ;
        RECT 70.880 156.975 71.210 157.355 ;
        RECT 71.810 156.975 72.070 157.815 ;
        RECT 74.080 156.975 74.305 157.435 ;
        RECT 74.995 156.975 75.245 157.775 ;
        RECT 75.925 156.975 76.215 157.700 ;
        RECT 77.355 156.975 77.605 157.775 ;
        RECT 91.565 157.745 92.775 158.265 ;
        RECT 78.295 156.975 78.520 157.435 ;
        RECT 81.335 156.975 81.620 157.435 ;
        RECT 82.750 156.975 83.410 157.455 ;
        RECT 85.020 156.975 85.340 157.435 ;
        RECT 86.080 156.975 86.490 157.415 ;
        RECT 88.315 156.975 88.645 157.355 ;
        RECT 89.255 156.975 89.585 157.355 ;
        RECT 90.185 156.975 92.775 157.745 ;
        RECT 93.005 156.975 93.215 157.795 ;
        RECT 93.885 156.975 94.115 157.795 ;
        RECT 95.245 157.745 95.995 158.265 ;
        RECT 99.865 157.745 101.515 158.265 ;
        RECT 103.985 157.745 105.195 158.265 ;
        RECT 94.325 156.975 95.995 157.745 ;
        RECT 96.605 156.975 96.935 157.355 ;
        RECT 98.005 156.975 101.515 157.745 ;
        RECT 101.685 156.975 101.975 157.700 ;
        RECT 102.605 156.975 105.195 157.745 ;
        RECT 107.435 157.725 107.955 158.265 ;
        RECT 105.805 156.975 106.135 157.355 ;
        RECT 106.745 156.975 107.955 157.725 ;
        RECT 111.550 157.520 111.890 158.350 ;
        RECT 117.070 157.520 117.410 158.350 ;
        RECT 108.130 156.975 113.475 157.520 ;
        RECT 113.650 156.975 118.995 157.520 ;
        RECT 119.315 156.975 119.645 157.775 ;
        RECT 124.705 157.745 126.355 158.265 ;
        RECT 120.155 156.975 120.485 157.455 ;
        RECT 121.075 156.975 121.315 157.455 ;
        RECT 122.845 156.975 126.355 157.745 ;
        RECT 127.215 157.725 127.735 158.265 ;
        RECT 126.525 156.975 127.735 157.725 ;
        RECT 14.660 156.805 127.820 156.975 ;
        RECT 14.745 156.055 15.955 156.805 ;
        RECT 17.395 156.345 17.680 156.805 ;
        RECT 18.810 156.325 19.470 156.805 ;
        RECT 21.080 156.345 21.400 156.805 ;
        RECT 22.140 156.365 22.550 156.805 ;
        RECT 24.375 156.425 24.705 156.805 ;
        RECT 25.315 156.425 25.645 156.805 ;
        RECT 26.685 156.425 27.015 156.805 ;
        RECT 14.745 155.515 15.265 156.055 ;
        RECT 28.545 156.035 32.055 156.805 ;
        RECT 32.795 156.345 33.065 156.805 ;
        RECT 34.855 156.345 35.180 156.805 ;
        RECT 35.905 156.055 37.115 156.805 ;
        RECT 37.285 156.080 37.575 156.805 ;
        RECT 30.405 155.515 32.055 156.035 ;
        RECT 36.595 155.515 37.115 156.055 ;
        RECT 38.205 156.035 39.875 156.805 ;
        RECT 39.125 155.515 39.875 156.035 ;
        RECT 40.555 156.005 40.805 156.805 ;
        RECT 41.495 156.345 41.720 156.805 ;
        RECT 44.235 156.005 44.485 156.805 ;
        RECT 45.175 156.345 45.400 156.805 ;
        RECT 49.240 156.345 49.465 156.805 ;
        RECT 50.155 156.005 50.405 156.805 ;
        RECT 51.545 156.035 53.215 156.805 ;
        RECT 54.195 156.345 54.480 156.805 ;
        RECT 55.610 156.325 56.270 156.805 ;
        RECT 57.880 156.345 58.200 156.805 ;
        RECT 58.940 156.365 59.350 156.805 ;
        RECT 61.175 156.425 61.505 156.805 ;
        RECT 62.115 156.425 62.445 156.805 ;
        RECT 63.045 156.080 63.335 156.805 ;
        RECT 52.465 155.515 53.215 156.035 ;
        RECT 63.545 155.985 63.775 156.805 ;
        RECT 64.445 155.985 64.655 156.805 ;
        RECT 64.885 156.035 66.555 156.805 ;
        RECT 66.815 156.325 67.115 156.805 ;
        RECT 67.715 156.325 67.975 156.805 ;
        RECT 68.585 156.325 68.835 156.805 ;
        RECT 69.445 156.325 69.695 156.805 ;
        RECT 70.305 156.325 70.550 156.805 ;
        RECT 71.165 156.325 71.410 156.805 ;
        RECT 72.010 156.325 72.270 156.805 ;
        RECT 72.870 156.325 73.130 156.805 ;
        RECT 73.730 156.245 73.990 156.805 ;
        RECT 74.590 156.280 74.850 156.805 ;
        RECT 75.450 156.295 75.755 156.805 ;
        RECT 77.760 156.345 77.985 156.805 ;
        RECT 65.805 155.515 66.555 156.035 ;
        RECT 78.675 156.005 78.925 156.805 ;
        RECT 81.035 156.005 81.285 156.805 ;
        RECT 81.975 156.345 82.200 156.805 ;
        RECT 85.125 156.035 88.635 156.805 ;
        RECT 88.805 156.080 89.095 156.805 ;
        RECT 89.265 156.035 91.855 156.805 ;
        RECT 92.030 156.260 97.375 156.805 ;
        RECT 86.985 155.515 88.635 156.035 ;
        RECT 90.645 155.515 91.855 156.035 ;
        RECT 95.450 155.430 95.790 156.260 ;
        RECT 98.055 156.005 98.305 156.805 ;
        RECT 98.995 156.345 99.220 156.805 ;
        RECT 101.685 156.035 103.355 156.805 ;
        RECT 105.360 156.345 105.585 156.805 ;
        RECT 102.605 155.515 103.355 156.035 ;
        RECT 106.275 156.005 106.525 156.805 ;
        RECT 109.040 156.345 109.265 156.805 ;
        RECT 109.955 156.005 110.205 156.805 ;
        RECT 111.395 156.005 111.645 156.805 ;
        RECT 112.335 156.345 112.560 156.805 ;
        RECT 114.565 156.080 114.855 156.805 ;
        RECT 115.025 156.055 116.235 156.805 ;
        RECT 116.845 156.325 117.085 156.805 ;
        RECT 117.675 156.325 118.005 156.805 ;
        RECT 115.715 155.515 116.235 156.055 ;
        RECT 118.515 156.005 118.845 156.805 ;
        RECT 119.165 156.035 120.835 156.805 ;
        RECT 121.010 156.260 126.355 156.805 ;
        RECT 120.085 155.515 120.835 156.035 ;
        RECT 124.430 155.430 124.770 156.260 ;
        RECT 126.525 156.055 127.735 156.805 ;
        RECT 127.215 155.515 127.735 156.055 ;
        RECT 14.745 152.285 15.265 152.825 ;
        RECT 18.445 152.305 20.095 152.825 ;
        RECT 14.745 151.535 15.955 152.285 ;
        RECT 16.585 151.535 20.095 152.305 ;
        RECT 21.005 151.535 21.515 152.070 ;
        RECT 23.475 151.535 23.805 151.935 ;
        RECT 24.405 151.535 24.695 152.260 ;
        RECT 28.750 152.080 29.090 152.910 ;
        RECT 25.330 151.535 30.675 152.080 ;
        RECT 30.885 151.535 31.115 152.355 ;
        RECT 31.785 151.535 31.995 152.355 ;
        RECT 32.665 151.535 32.995 151.915 ;
        RECT 34.035 151.535 34.365 151.935 ;
        RECT 36.325 151.535 36.835 152.070 ;
        RECT 38.255 151.535 38.505 152.335 ;
        RECT 43.265 152.305 44.475 152.825 ;
        RECT 39.195 151.535 39.420 151.995 ;
        RECT 41.885 151.535 44.475 152.305 ;
        RECT 48.070 152.080 48.410 152.910 ;
        RECT 44.650 151.535 49.995 152.080 ;
        RECT 50.165 151.535 50.455 152.260 ;
        RECT 54.970 152.080 55.310 152.910 ;
        RECT 51.550 151.535 56.895 152.080 ;
        RECT 57.105 151.535 57.335 152.355 ;
        RECT 58.005 151.535 58.215 152.355 ;
        RECT 69.945 152.305 71.155 152.825 ;
        RECT 59.255 151.535 59.540 151.995 ;
        RECT 60.670 151.535 61.330 152.015 ;
        RECT 62.940 151.535 63.260 151.995 ;
        RECT 64.000 151.535 64.410 151.975 ;
        RECT 66.235 151.535 66.565 151.915 ;
        RECT 67.175 151.535 67.505 151.915 ;
        RECT 68.565 151.535 71.155 152.305 ;
        RECT 71.800 151.535 72.130 151.915 ;
        RECT 72.730 151.535 72.990 152.375 ;
        RECT 78.225 152.305 79.435 152.825 ;
        RECT 73.675 151.535 74.005 151.895 ;
        RECT 75.925 151.535 76.215 152.260 ;
        RECT 76.845 151.535 79.435 152.305 ;
        RECT 83.030 152.080 83.370 152.910 ;
        RECT 88.550 152.080 88.890 152.910 ;
        RECT 79.610 151.535 84.955 152.080 ;
        RECT 85.130 151.535 90.475 152.080 ;
        RECT 90.685 151.535 90.915 152.355 ;
        RECT 91.585 151.535 91.795 152.355 ;
        RECT 94.345 152.305 95.995 152.825 ;
        RECT 92.485 151.535 95.995 152.305 ;
        RECT 99.590 152.080 99.930 152.910 ;
        RECT 103.985 152.305 105.195 152.825 ;
        RECT 96.170 151.535 101.515 152.080 ;
        RECT 101.685 151.535 101.975 152.260 ;
        RECT 102.605 151.535 105.195 152.305 ;
        RECT 105.875 151.535 106.125 152.335 ;
        RECT 106.815 151.535 107.040 151.995 ;
        RECT 109.555 151.535 109.805 152.335 ;
        RECT 116.610 152.080 116.950 152.910 ;
        RECT 110.495 151.535 110.720 151.995 ;
        RECT 113.190 151.535 118.535 152.080 ;
        RECT 118.765 151.535 118.975 152.355 ;
        RECT 119.645 151.535 119.875 152.355 ;
        RECT 124.705 152.305 126.355 152.825 ;
        RECT 120.985 151.535 121.315 151.915 ;
        RECT 122.845 151.535 126.355 152.305 ;
        RECT 127.215 152.285 127.735 152.825 ;
        RECT 126.525 151.535 127.735 152.285 ;
        RECT 14.660 151.365 127.820 151.535 ;
        RECT 14.745 150.615 15.955 151.365 ;
        RECT 16.935 150.905 17.220 151.365 ;
        RECT 18.350 150.885 19.010 151.365 ;
        RECT 20.620 150.905 20.940 151.365 ;
        RECT 21.680 150.925 22.090 151.365 ;
        RECT 23.915 150.985 24.245 151.365 ;
        RECT 24.855 150.985 25.185 151.365 ;
        RECT 14.745 150.075 15.265 150.615 ;
        RECT 25.785 150.595 27.455 151.365 ;
        RECT 28.435 150.905 28.720 151.365 ;
        RECT 29.850 150.885 30.510 151.365 ;
        RECT 32.120 150.905 32.440 151.365 ;
        RECT 33.180 150.925 33.590 151.365 ;
        RECT 35.415 150.985 35.745 151.365 ;
        RECT 36.355 150.985 36.685 151.365 ;
        RECT 37.285 150.640 37.575 151.365 ;
        RECT 38.205 150.595 40.795 151.365 ;
        RECT 42.800 150.905 43.025 151.365 ;
        RECT 26.705 150.075 27.455 150.595 ;
        RECT 39.585 150.075 40.795 150.595 ;
        RECT 43.715 150.565 43.965 151.365 ;
        RECT 44.645 150.615 45.855 151.365 ;
        RECT 46.035 150.865 46.365 151.365 ;
        RECT 46.935 150.965 47.265 151.365 ;
        RECT 47.775 150.965 48.155 151.365 ;
        RECT 48.795 150.865 49.125 151.365 ;
        RECT 49.695 150.965 50.025 151.365 ;
        RECT 50.535 150.965 50.915 151.365 ;
        RECT 45.335 150.075 45.855 150.615 ;
        RECT 52.055 150.565 52.305 151.365 ;
        RECT 52.995 150.905 53.220 151.365 ;
        RECT 55.685 150.595 57.355 151.365 ;
        RECT 58.265 150.830 58.775 151.365 ;
        RECT 60.735 150.965 61.065 151.365 ;
        RECT 62.105 150.985 62.435 151.365 ;
        RECT 63.045 150.640 63.335 151.365 ;
        RECT 64.405 150.985 64.735 151.365 ;
        RECT 65.805 150.595 67.475 151.365 ;
        RECT 68.120 150.985 68.450 151.365 ;
        RECT 56.605 150.075 57.355 150.595 ;
        RECT 66.725 150.075 67.475 150.595 ;
        RECT 69.050 150.525 69.310 151.365 ;
        RECT 69.490 150.525 69.750 151.365 ;
        RECT 70.350 150.985 70.680 151.365 ;
        RECT 71.385 150.885 71.665 151.365 ;
        RECT 72.270 150.885 72.525 151.365 ;
        RECT 73.170 150.885 73.445 151.365 ;
        RECT 75.475 150.885 75.750 151.365 ;
        RECT 76.395 150.885 76.650 151.365 ;
        RECT 77.255 150.885 77.535 151.365 ;
        RECT 77.775 150.865 78.105 151.365 ;
        RECT 78.675 150.965 79.005 151.365 ;
        RECT 79.515 150.965 79.895 151.365 ;
        RECT 80.985 150.595 84.495 151.365 ;
        RECT 85.405 150.830 85.915 151.365 ;
        RECT 87.875 150.965 88.205 151.365 ;
        RECT 88.805 150.640 89.095 151.365 ;
        RECT 89.695 150.985 90.025 151.365 ;
        RECT 90.635 150.985 90.965 151.365 ;
        RECT 92.790 150.925 93.200 151.365 ;
        RECT 93.940 150.905 94.260 151.365 ;
        RECT 95.870 150.885 96.530 151.365 ;
        RECT 97.660 150.905 97.945 151.365 ;
        RECT 98.930 150.820 104.275 151.365 ;
        RECT 104.905 150.965 105.285 151.365 ;
        RECT 105.795 150.965 106.125 151.365 ;
        RECT 106.695 150.865 107.025 151.365 ;
        RECT 82.845 150.075 84.495 150.595 ;
        RECT 102.350 149.990 102.690 150.820 ;
        RECT 107.715 150.565 107.965 151.365 ;
        RECT 108.655 150.905 108.880 151.365 ;
        RECT 111.455 150.905 111.725 151.365 ;
        RECT 113.515 150.905 113.840 151.365 ;
        RECT 114.565 150.640 114.855 151.365 ;
        RECT 116.375 150.905 116.680 151.365 ;
        RECT 118.165 150.925 118.355 151.365 ;
        RECT 120.255 150.905 120.585 151.365 ;
        RECT 123.185 151.005 123.515 151.365 ;
        RECT 124.215 150.985 124.545 151.365 ;
        RECT 125.145 150.615 126.355 151.365 ;
        RECT 126.525 150.615 127.735 151.365 ;
        RECT 125.835 150.075 126.355 150.615 ;
        RECT 127.215 150.075 127.735 150.615 ;
        RECT 14.745 146.845 15.265 147.385 ;
        RECT 18.445 146.865 20.095 147.385 ;
        RECT 14.745 146.095 15.955 146.845 ;
        RECT 16.585 146.095 20.095 146.865 ;
        RECT 21.005 146.095 21.515 146.630 ;
        RECT 23.475 146.095 23.805 146.495 ;
        RECT 24.405 146.095 24.695 146.820 ;
        RECT 25.365 146.095 25.595 146.915 ;
        RECT 26.265 146.095 26.475 146.915 ;
        RECT 34.985 146.865 35.735 147.385 ;
        RECT 27.145 146.095 27.475 146.475 ;
        RECT 28.525 146.095 28.855 146.475 ;
        RECT 29.895 146.095 30.225 146.495 ;
        RECT 32.185 146.095 32.695 146.630 ;
        RECT 34.065 146.095 35.735 146.865 ;
        RECT 37.740 146.095 37.965 146.555 ;
        RECT 38.655 146.095 38.905 146.895 ;
        RECT 40.095 146.095 40.345 146.895 ;
        RECT 43.955 146.845 44.475 147.385 ;
        RECT 41.035 146.095 41.260 146.555 ;
        RECT 43.265 146.095 44.475 146.845 ;
        RECT 48.070 146.640 48.410 147.470 ;
        RECT 44.650 146.095 49.995 146.640 ;
        RECT 50.165 146.095 50.455 146.820 ;
        RECT 51.975 146.095 52.305 146.495 ;
        RECT 54.265 146.095 54.775 146.630 ;
        RECT 56.195 146.095 56.445 146.895 ;
        RECT 64.655 146.845 65.175 147.385 ;
        RECT 57.135 146.095 57.360 146.555 ;
        RECT 60.565 146.095 61.075 146.630 ;
        RECT 63.035 146.095 63.365 146.495 ;
        RECT 63.965 146.095 65.175 146.845 ;
        RECT 68.770 146.640 69.110 147.470 ;
        RECT 65.350 146.095 70.695 146.640 ;
        RECT 70.870 146.095 71.130 146.935 ;
        RECT 71.730 146.095 72.060 146.475 ;
        RECT 73.180 146.095 73.510 146.475 ;
        RECT 74.110 146.095 74.370 146.935 ;
        RECT 75.235 146.845 75.755 147.385 ;
        RECT 74.545 146.095 75.755 146.845 ;
        RECT 75.925 146.095 76.215 146.820 ;
        RECT 78.220 146.095 78.445 146.555 ;
        RECT 79.135 146.095 79.385 146.895 ;
        RECT 80.575 146.095 80.825 146.895 ;
        RECT 81.515 146.095 81.740 146.555 ;
        RECT 83.805 146.095 84.015 146.915 ;
        RECT 84.685 146.095 84.915 146.915 ;
        RECT 85.935 146.095 86.220 146.555 ;
        RECT 87.350 146.095 88.010 146.575 ;
        RECT 89.620 146.095 89.940 146.555 ;
        RECT 90.680 146.095 91.090 146.535 ;
        RECT 92.915 146.095 93.245 146.475 ;
        RECT 93.855 146.095 94.185 146.475 ;
        RECT 95.745 146.095 95.975 146.915 ;
        RECT 96.645 146.095 96.855 146.915 ;
        RECT 97.825 146.095 98.335 146.630 ;
        RECT 100.295 146.095 100.625 146.495 ;
        RECT 101.685 146.095 101.975 146.820 ;
        RECT 102.585 146.095 102.915 146.475 ;
        RECT 104.445 146.095 104.825 146.495 ;
        RECT 105.335 146.095 105.665 146.495 ;
        RECT 106.235 146.095 106.565 146.595 ;
        RECT 107.255 146.095 107.505 146.895 ;
        RECT 111.345 146.865 112.095 147.385 ;
        RECT 108.195 146.095 108.420 146.555 ;
        RECT 110.425 146.095 112.095 146.865 ;
        RECT 127.215 146.845 127.735 147.385 ;
        RECT 113.005 146.095 113.515 146.630 ;
        RECT 115.475 146.095 115.805 146.495 ;
        RECT 117.215 146.095 117.500 146.555 ;
        RECT 118.630 146.095 119.290 146.575 ;
        RECT 120.900 146.095 121.220 146.555 ;
        RECT 121.960 146.095 122.370 146.535 ;
        RECT 124.195 146.095 124.525 146.475 ;
        RECT 125.135 146.095 125.465 146.475 ;
        RECT 126.525 146.095 127.735 146.845 ;
        RECT 14.660 145.925 127.820 146.095 ;
        RECT 14.745 145.175 15.955 145.925 ;
        RECT 14.745 144.635 15.265 145.175 ;
        RECT 16.585 145.155 20.095 145.925 ;
        RECT 18.445 144.635 20.095 145.155 ;
        RECT 20.325 145.105 20.535 145.925 ;
        RECT 21.205 145.105 21.435 145.925 ;
        RECT 22.915 145.465 23.200 145.925 ;
        RECT 24.330 145.445 24.990 145.925 ;
        RECT 26.600 145.465 26.920 145.925 ;
        RECT 27.660 145.485 28.070 145.925 ;
        RECT 29.895 145.545 30.225 145.925 ;
        RECT 30.835 145.545 31.165 145.925 ;
        RECT 31.770 145.380 37.115 145.925 ;
        RECT 35.190 144.550 35.530 145.380 ;
        RECT 37.285 145.200 37.575 145.925 ;
        RECT 38.205 145.155 40.795 145.925 ;
        RECT 39.585 144.635 40.795 145.155 ;
        RECT 41.005 145.105 41.235 145.925 ;
        RECT 41.905 145.105 42.115 145.925 ;
        RECT 42.775 145.545 43.105 145.925 ;
        RECT 43.715 145.545 44.045 145.925 ;
        RECT 45.870 145.485 46.280 145.925 ;
        RECT 47.020 145.465 47.340 145.925 ;
        RECT 48.950 145.445 49.610 145.925 ;
        RECT 50.740 145.465 51.025 145.925 ;
        RECT 52.445 145.545 52.775 145.925 ;
        RECT 53.385 145.175 54.595 145.925 ;
        RECT 54.075 144.635 54.595 145.175 ;
        RECT 54.765 145.155 58.275 145.925 ;
        RECT 56.625 144.635 58.275 145.155 ;
        RECT 58.485 145.105 58.715 145.925 ;
        RECT 59.385 145.105 59.595 145.925 ;
        RECT 60.285 145.155 62.875 145.925 ;
        RECT 63.045 145.200 63.335 145.925 ;
        RECT 64.705 145.390 65.215 145.925 ;
        RECT 67.175 145.525 67.505 145.925 ;
        RECT 68.570 145.380 73.915 145.925 ;
        RECT 74.090 145.380 79.435 145.925 ;
        RECT 79.615 145.425 79.945 145.925 ;
        RECT 80.515 145.525 80.845 145.925 ;
        RECT 81.355 145.525 81.735 145.925 ;
        RECT 61.665 144.635 62.875 145.155 ;
        RECT 71.990 144.550 72.330 145.380 ;
        RECT 77.510 144.550 77.850 145.380 ;
        RECT 82.825 145.155 84.495 145.925 ;
        RECT 85.405 145.390 85.915 145.925 ;
        RECT 87.875 145.525 88.205 145.925 ;
        RECT 88.805 145.200 89.095 145.925 ;
        RECT 90.625 145.545 90.955 145.925 ;
        RECT 92.005 145.545 92.335 145.925 ;
        RECT 93.515 145.465 93.785 145.925 ;
        RECT 95.575 145.465 95.900 145.925 ;
        RECT 97.055 145.465 97.360 145.925 ;
        RECT 98.845 145.485 99.035 145.925 ;
        RECT 100.935 145.465 101.265 145.925 ;
        RECT 103.865 145.565 104.195 145.925 ;
        RECT 104.895 145.545 105.225 145.925 ;
        RECT 106.285 145.155 109.795 145.925 ;
        RECT 111.800 145.465 112.025 145.925 ;
        RECT 83.745 144.635 84.495 145.155 ;
        RECT 108.145 144.635 109.795 145.155 ;
        RECT 112.715 145.125 112.965 145.925 ;
        RECT 114.565 145.200 114.855 145.925 ;
        RECT 116.225 145.390 116.735 145.925 ;
        RECT 118.695 145.525 119.025 145.925 ;
        RECT 119.665 145.105 119.895 145.925 ;
        RECT 120.565 145.105 120.775 145.925 ;
        RECT 121.905 145.545 122.235 145.925 ;
        RECT 122.845 145.155 126.355 145.925 ;
        RECT 126.525 145.175 127.735 145.925 ;
        RECT 124.705 144.635 126.355 145.155 ;
        RECT 127.215 144.635 127.735 145.175 ;
        RECT 14.745 141.405 15.265 141.945 ;
        RECT 17.505 141.425 18.715 141.945 ;
        RECT 14.745 140.655 15.955 141.405 ;
        RECT 16.125 140.655 18.715 141.425 ;
        RECT 22.310 141.200 22.650 142.030 ;
        RECT 27.185 141.425 28.835 141.945 ;
        RECT 18.890 140.655 24.235 141.200 ;
        RECT 24.405 140.655 24.695 141.380 ;
        RECT 25.325 140.655 28.835 141.425 ;
        RECT 32.430 141.200 32.770 142.030 ;
        RECT 40.065 141.425 41.715 141.945 ;
        RECT 29.010 140.655 34.355 141.200 ;
        RECT 34.985 140.655 35.365 141.055 ;
        RECT 35.875 140.655 36.205 141.055 ;
        RECT 36.775 140.655 37.105 141.155 ;
        RECT 38.205 140.655 41.715 141.425 ;
        RECT 45.310 141.200 45.650 142.030 ;
        RECT 51.545 141.425 52.295 141.945 ;
        RECT 41.890 140.655 47.235 141.200 ;
        RECT 47.415 140.655 47.745 141.155 ;
        RECT 48.315 140.655 48.645 141.055 ;
        RECT 49.155 140.655 49.535 141.055 ;
        RECT 50.165 140.655 50.455 141.380 ;
        RECT 50.625 140.655 52.295 141.425 ;
        RECT 52.975 140.655 53.225 141.455 ;
        RECT 71.095 141.405 71.615 141.945 ;
        RECT 53.915 140.655 54.140 141.115 ;
        RECT 56.715 140.655 56.985 141.115 ;
        RECT 58.775 140.655 59.100 141.115 ;
        RECT 60.255 140.655 60.560 141.115 ;
        RECT 62.045 140.655 62.235 141.095 ;
        RECT 64.135 140.655 64.465 141.115 ;
        RECT 67.065 140.655 67.395 141.015 ;
        RECT 68.095 140.655 68.425 141.035 ;
        RECT 69.465 140.655 69.795 141.035 ;
        RECT 70.405 140.655 71.615 141.405 ;
        RECT 71.825 140.655 72.055 141.475 ;
        RECT 72.725 140.655 72.935 141.475 ;
        RECT 74.545 141.425 75.755 141.945 ;
        RECT 78.225 141.425 79.435 141.945 ;
        RECT 73.165 140.655 75.755 141.425 ;
        RECT 75.925 140.655 76.215 141.380 ;
        RECT 76.845 140.655 79.435 141.425 ;
        RECT 83.030 141.200 83.370 142.030 ;
        RECT 88.550 141.200 88.890 142.030 ;
        RECT 94.070 141.200 94.410 142.030 ;
        RECT 99.590 141.200 99.930 142.030 ;
        RECT 79.610 140.655 84.955 141.200 ;
        RECT 85.130 140.655 90.475 141.200 ;
        RECT 90.650 140.655 95.995 141.200 ;
        RECT 96.170 140.655 101.515 141.200 ;
        RECT 101.685 140.655 101.975 141.380 ;
        RECT 106.490 141.200 106.830 142.030 ;
        RECT 114.125 141.425 115.775 141.945 ;
        RECT 103.070 140.655 108.415 141.200 ;
        RECT 108.595 140.655 108.925 141.155 ;
        RECT 109.495 140.655 109.825 141.055 ;
        RECT 110.335 140.655 110.715 141.055 ;
        RECT 112.265 140.655 115.775 141.425 ;
        RECT 116.685 140.655 117.195 141.190 ;
        RECT 119.155 140.655 119.485 141.055 ;
        RECT 120.125 140.655 120.355 141.475 ;
        RECT 121.025 140.655 121.235 141.475 ;
        RECT 122.155 141.405 122.675 141.945 ;
        RECT 124.705 141.425 126.355 141.945 ;
        RECT 121.465 140.655 122.675 141.405 ;
        RECT 122.845 140.655 126.355 141.425 ;
        RECT 127.215 141.405 127.735 141.945 ;
        RECT 126.525 140.655 127.735 141.405 ;
        RECT 14.660 140.485 127.820 140.655 ;
        RECT 14.745 139.735 15.955 140.485 ;
        RECT 16.935 140.025 17.220 140.485 ;
        RECT 18.350 140.005 19.010 140.485 ;
        RECT 20.620 140.025 20.940 140.485 ;
        RECT 21.680 140.045 22.090 140.485 ;
        RECT 23.915 140.105 24.245 140.485 ;
        RECT 24.855 140.105 25.185 140.485 ;
        RECT 14.745 139.195 15.265 139.735 ;
        RECT 25.785 139.715 28.375 140.485 ;
        RECT 28.550 139.940 33.895 140.485 ;
        RECT 35.215 140.025 35.465 140.485 ;
        RECT 27.165 139.195 28.375 139.715 ;
        RECT 31.970 139.110 32.310 139.940 ;
        RECT 37.285 139.760 37.575 140.485 ;
        RECT 39.125 140.085 39.505 140.485 ;
        RECT 40.015 140.085 40.345 140.485 ;
        RECT 40.915 139.985 41.245 140.485 ;
        RECT 41.430 139.940 46.775 140.485 ;
        RECT 46.955 139.985 47.285 140.485 ;
        RECT 47.855 140.085 48.185 140.485 ;
        RECT 48.695 140.085 49.075 140.485 ;
        RECT 44.850 139.110 45.190 139.940 ;
        RECT 50.215 139.685 50.465 140.485 ;
        RECT 51.155 140.025 51.380 140.485 ;
        RECT 53.385 139.715 55.055 140.485 ;
        RECT 54.305 139.195 55.055 139.715 ;
        RECT 55.265 139.665 55.495 140.485 ;
        RECT 56.165 139.665 56.375 140.485 ;
        RECT 56.605 139.715 59.195 140.485 ;
        RECT 57.985 139.195 59.195 139.715 ;
        RECT 59.875 139.685 60.125 140.485 ;
        RECT 60.815 140.025 61.040 140.485 ;
        RECT 63.045 139.760 63.335 140.485 ;
        RECT 64.475 139.685 64.725 140.485 ;
        RECT 65.415 140.025 65.640 140.485 ;
        RECT 68.075 140.105 68.405 140.485 ;
        RECT 69.015 140.105 69.345 140.485 ;
        RECT 71.170 140.045 71.580 140.485 ;
        RECT 72.320 140.025 72.640 140.485 ;
        RECT 74.250 140.005 74.910 140.485 ;
        RECT 76.040 140.025 76.325 140.485 ;
        RECT 77.305 139.715 79.895 140.485 ;
        RECT 78.685 139.195 79.895 139.715 ;
        RECT 80.575 139.685 80.825 140.485 ;
        RECT 81.515 140.025 81.740 140.485 ;
        RECT 85.405 139.950 85.915 140.485 ;
        RECT 87.875 140.085 88.205 140.485 ;
        RECT 88.805 139.760 89.095 140.485 ;
        RECT 90.165 140.105 90.495 140.485 ;
        RECT 92.025 139.715 95.535 140.485 ;
        RECT 95.710 139.940 101.055 140.485 ;
        RECT 93.885 139.195 95.535 139.715 ;
        RECT 99.130 139.110 99.470 139.940 ;
        RECT 101.265 139.665 101.495 140.485 ;
        RECT 102.165 139.665 102.375 140.485 ;
        RECT 102.605 139.715 106.115 140.485 ;
        RECT 104.465 139.195 106.115 139.715 ;
        RECT 106.795 139.685 107.045 140.485 ;
        RECT 107.735 140.025 107.960 140.485 ;
        RECT 111.800 140.025 112.025 140.485 ;
        RECT 112.715 139.685 112.965 140.485 ;
        RECT 114.565 139.760 114.855 140.485 ;
        RECT 115.525 139.665 115.755 140.485 ;
        RECT 116.425 139.665 116.635 140.485 ;
        RECT 117.675 140.025 117.960 140.485 ;
        RECT 119.090 140.005 119.750 140.485 ;
        RECT 121.360 140.025 121.680 140.485 ;
        RECT 122.420 140.045 122.830 140.485 ;
        RECT 124.655 140.105 124.985 140.485 ;
        RECT 125.595 140.105 125.925 140.485 ;
        RECT 126.525 139.735 127.735 140.485 ;
        RECT 127.215 139.195 127.735 139.735 ;
        RECT 14.745 135.965 15.265 136.505 ;
        RECT 14.745 135.215 15.955 135.965 ;
        RECT 19.550 135.760 19.890 136.590 ;
        RECT 16.130 135.215 21.475 135.760 ;
        RECT 22.085 135.215 22.415 135.595 ;
        RECT 23.065 135.215 23.295 136.035 ;
        RECT 23.965 135.215 24.175 136.035 ;
        RECT 27.185 135.985 28.835 136.505 ;
        RECT 34.065 135.985 34.815 136.505 ;
        RECT 41.905 135.985 43.555 136.505 ;
        RECT 48.345 135.985 49.995 136.505 ;
        RECT 52.005 135.985 52.755 136.505 ;
        RECT 60.285 135.985 61.035 136.505 ;
        RECT 24.405 135.215 24.695 135.940 ;
        RECT 25.325 135.215 28.835 135.985 ;
        RECT 29.745 135.215 30.255 135.750 ;
        RECT 32.215 135.215 32.545 135.615 ;
        RECT 33.145 135.215 34.815 135.985 ;
        RECT 35.445 135.215 35.825 135.615 ;
        RECT 36.335 135.215 36.665 135.615 ;
        RECT 37.235 135.215 37.565 135.715 ;
        RECT 38.895 135.215 39.145 135.675 ;
        RECT 40.045 135.215 43.555 135.985 ;
        RECT 44.185 135.215 44.565 135.615 ;
        RECT 45.075 135.215 45.405 135.615 ;
        RECT 45.975 135.215 46.305 135.715 ;
        RECT 46.485 135.215 49.995 135.985 ;
        RECT 50.165 135.215 50.455 135.940 ;
        RECT 51.085 135.215 52.755 135.985 ;
        RECT 53.665 135.215 54.175 135.750 ;
        RECT 56.135 135.215 56.465 135.615 ;
        RECT 57.965 135.215 58.295 135.595 ;
        RECT 59.365 135.215 61.035 135.985 ;
        RECT 61.715 135.215 61.965 136.015 ;
        RECT 66.265 135.985 67.015 136.505 ;
        RECT 75.005 135.985 75.755 136.505 ;
        RECT 62.655 135.215 62.880 135.675 ;
        RECT 65.345 135.215 67.015 135.985 ;
        RECT 67.615 135.215 67.945 135.575 ;
        RECT 69.775 135.215 70.230 135.980 ;
        RECT 70.960 135.215 71.285 135.675 ;
        RECT 73.075 135.215 73.345 135.675 ;
        RECT 74.085 135.215 75.755 135.985 ;
        RECT 75.925 135.215 76.215 135.940 ;
        RECT 77.765 135.215 78.145 135.615 ;
        RECT 78.655 135.215 78.985 135.615 ;
        RECT 79.555 135.215 79.885 135.715 ;
        RECT 80.575 135.215 80.825 136.015 ;
        RECT 81.515 135.215 81.740 135.675 ;
        RECT 84.555 135.215 84.840 135.675 ;
        RECT 85.970 135.215 86.630 135.695 ;
        RECT 88.240 135.215 88.560 135.675 ;
        RECT 89.300 135.215 89.710 135.655 ;
        RECT 91.535 135.215 91.865 135.595 ;
        RECT 92.475 135.215 92.805 135.595 ;
        RECT 94.145 135.215 94.655 135.750 ;
        RECT 96.615 135.215 96.945 135.615 ;
        RECT 99.840 135.215 100.065 135.675 ;
        RECT 100.755 135.215 101.005 136.015 ;
        RECT 125.605 135.985 126.355 136.505 ;
        RECT 101.685 135.215 101.975 135.940 ;
        RECT 103.805 135.215 104.315 135.750 ;
        RECT 106.275 135.215 106.605 135.615 ;
        RECT 107.645 135.215 107.975 135.595 ;
        RECT 110.245 135.215 110.755 135.750 ;
        RECT 112.715 135.215 113.045 135.615 ;
        RECT 114.455 135.215 114.740 135.675 ;
        RECT 115.870 135.215 116.530 135.695 ;
        RECT 118.140 135.215 118.460 135.675 ;
        RECT 119.200 135.215 119.610 135.655 ;
        RECT 121.435 135.215 121.765 135.595 ;
        RECT 122.375 135.215 122.705 135.595 ;
        RECT 123.745 135.215 124.075 135.595 ;
        RECT 124.685 135.215 126.355 135.985 ;
        RECT 127.215 135.965 127.735 136.505 ;
        RECT 126.525 135.215 127.735 135.965 ;
        RECT 14.660 135.045 127.820 135.215 ;
        RECT 14.745 134.295 15.955 135.045 ;
        RECT 14.745 133.755 15.265 134.295 ;
        RECT 16.185 134.225 16.395 135.045 ;
        RECT 17.065 134.225 17.295 135.045 ;
        RECT 18.245 134.510 18.755 135.045 ;
        RECT 20.715 134.645 21.045 135.045 ;
        RECT 22.455 134.585 22.740 135.045 ;
        RECT 23.870 134.565 24.530 135.045 ;
        RECT 26.140 134.585 26.460 135.045 ;
        RECT 27.200 134.605 27.610 135.045 ;
        RECT 29.435 134.665 29.765 135.045 ;
        RECT 30.375 134.665 30.705 135.045 ;
        RECT 31.745 134.665 32.075 135.045 ;
        RECT 33.885 134.510 34.395 135.045 ;
        RECT 36.355 134.645 36.685 135.045 ;
        RECT 37.285 134.320 37.575 135.045 ;
        RECT 38.205 134.645 38.585 135.045 ;
        RECT 39.095 134.645 39.425 135.045 ;
        RECT 39.995 134.545 40.325 135.045 ;
        RECT 40.505 134.295 41.715 135.045 ;
        RECT 41.895 134.545 42.225 135.045 ;
        RECT 42.795 134.645 43.125 135.045 ;
        RECT 43.635 134.645 44.015 135.045 ;
        RECT 41.195 133.755 41.715 134.295 ;
        RECT 45.155 134.245 45.405 135.045 ;
        RECT 46.095 134.585 46.320 135.045 ;
        RECT 48.835 134.245 49.085 135.045 ;
        RECT 49.775 134.585 50.000 135.045 ;
        RECT 52.815 134.585 53.100 135.045 ;
        RECT 54.230 134.565 54.890 135.045 ;
        RECT 56.500 134.585 56.820 135.045 ;
        RECT 57.560 134.605 57.970 135.045 ;
        RECT 59.795 134.665 60.125 135.045 ;
        RECT 60.735 134.665 61.065 135.045 ;
        RECT 61.665 134.295 62.875 135.045 ;
        RECT 63.045 134.320 63.335 135.045 ;
        RECT 62.355 133.755 62.875 134.295 ;
        RECT 64.015 134.245 64.265 135.045 ;
        RECT 64.955 134.585 65.180 135.045 ;
        RECT 68.110 134.500 73.455 135.045 ;
        RECT 73.630 134.500 78.975 135.045 ;
        RECT 79.155 134.545 79.485 135.045 ;
        RECT 80.055 134.645 80.385 135.045 ;
        RECT 80.895 134.645 81.275 135.045 ;
        RECT 81.910 134.500 87.255 135.045 ;
        RECT 71.530 133.670 71.870 134.500 ;
        RECT 77.050 133.670 77.390 134.500 ;
        RECT 85.330 133.670 85.670 134.500 ;
        RECT 87.485 134.225 87.695 135.045 ;
        RECT 88.365 134.225 88.595 135.045 ;
        RECT 88.805 134.320 89.095 135.045 ;
        RECT 90.075 134.585 90.360 135.045 ;
        RECT 91.490 134.565 92.150 135.045 ;
        RECT 93.760 134.585 94.080 135.045 ;
        RECT 94.820 134.605 95.230 135.045 ;
        RECT 97.055 134.665 97.385 135.045 ;
        RECT 97.995 134.665 98.325 135.045 ;
        RECT 99.735 134.585 100.020 135.045 ;
        RECT 101.150 134.565 101.810 135.045 ;
        RECT 103.420 134.585 103.740 135.045 ;
        RECT 104.480 134.605 104.890 135.045 ;
        RECT 106.715 134.665 107.045 135.045 ;
        RECT 107.655 134.665 107.985 135.045 ;
        RECT 108.595 134.545 108.925 135.045 ;
        RECT 109.495 134.645 109.825 135.045 ;
        RECT 110.335 134.645 110.715 135.045 ;
        RECT 111.805 134.275 114.395 135.045 ;
        RECT 114.565 134.320 114.855 135.045 ;
        RECT 115.485 134.275 118.995 135.045 ;
        RECT 119.605 134.665 119.935 135.045 ;
        RECT 121.010 134.500 126.355 135.045 ;
        RECT 113.185 133.755 114.395 134.275 ;
        RECT 117.345 133.755 118.995 134.275 ;
        RECT 124.430 133.670 124.770 134.500 ;
        RECT 126.525 134.295 127.735 135.045 ;
        RECT 127.215 133.755 127.735 134.295 ;
        RECT 14.745 130.525 15.265 131.065 ;
        RECT 18.445 130.545 20.095 131.065 ;
        RECT 14.745 129.775 15.955 130.525 ;
        RECT 16.585 129.775 20.095 130.545 ;
        RECT 21.005 129.775 21.515 130.310 ;
        RECT 23.475 129.775 23.805 130.175 ;
        RECT 24.405 129.775 24.695 130.500 ;
        RECT 28.290 130.320 28.630 131.150 ;
        RECT 42.115 130.525 42.635 131.065 ;
        RECT 48.785 130.545 49.995 131.065 ;
        RECT 52.485 130.545 54.135 131.065 ;
        RECT 24.870 129.775 30.215 130.320 ;
        RECT 31.195 129.775 31.480 130.235 ;
        RECT 32.610 129.775 33.270 130.255 ;
        RECT 34.880 129.775 35.200 130.235 ;
        RECT 35.940 129.775 36.350 130.215 ;
        RECT 38.175 129.775 38.505 130.155 ;
        RECT 39.115 129.775 39.445 130.155 ;
        RECT 40.485 129.775 40.815 130.155 ;
        RECT 41.425 129.775 42.635 130.525 ;
        RECT 43.955 129.775 44.205 130.235 ;
        RECT 46.255 129.775 46.505 130.235 ;
        RECT 47.405 129.775 49.995 130.545 ;
        RECT 50.165 129.775 50.455 130.500 ;
        RECT 50.625 129.775 54.135 130.545 ;
        RECT 57.730 130.320 58.070 131.150 ;
        RECT 63.250 130.320 63.590 131.150 ;
        RECT 77.765 130.545 78.515 131.065 ;
        RECT 54.310 129.775 59.655 130.320 ;
        RECT 59.830 129.775 65.175 130.320 ;
        RECT 66.085 129.775 66.595 130.310 ;
        RECT 68.555 129.775 68.885 130.175 ;
        RECT 69.950 129.775 70.285 130.175 ;
        RECT 70.870 129.775 71.145 130.255 ;
        RECT 72.515 129.775 72.765 130.235 ;
        RECT 74.555 129.775 74.830 130.255 ;
        RECT 75.415 129.775 75.750 130.175 ;
        RECT 75.925 129.775 76.215 130.500 ;
        RECT 76.845 129.775 78.515 130.545 ;
        RECT 81.675 130.525 82.195 131.065 ;
        RECT 79.415 129.775 79.665 130.235 ;
        RECT 80.985 129.775 82.195 130.525 ;
        RECT 85.790 130.320 86.130 131.150 ;
        RECT 82.370 129.775 87.715 130.320 ;
        RECT 87.925 129.775 88.155 130.595 ;
        RECT 88.825 129.775 89.035 130.595 ;
        RECT 97.315 130.525 97.835 131.065 ;
        RECT 103.065 130.545 103.815 131.065 ;
        RECT 108.605 130.545 110.255 131.065 ;
        RECT 114.105 130.545 115.315 131.065 ;
        RECT 90.005 129.775 90.515 130.310 ;
        RECT 92.475 129.775 92.805 130.175 ;
        RECT 94.305 129.775 94.635 130.155 ;
        RECT 95.685 129.775 96.015 130.155 ;
        RECT 96.625 129.775 97.835 130.525 ;
        RECT 98.465 129.775 98.845 130.175 ;
        RECT 99.355 129.775 99.685 130.175 ;
        RECT 100.255 129.775 100.585 130.275 ;
        RECT 101.685 129.775 101.975 130.500 ;
        RECT 102.145 129.775 103.815 130.545 ;
        RECT 103.995 129.775 104.325 130.275 ;
        RECT 104.895 129.775 105.225 130.175 ;
        RECT 105.735 129.775 106.115 130.175 ;
        RECT 106.745 129.775 110.255 130.545 ;
        RECT 111.155 129.775 111.405 130.235 ;
        RECT 112.725 129.775 115.315 130.545 ;
        RECT 118.910 130.320 119.250 131.150 ;
        RECT 124.430 130.320 124.770 131.150 ;
        RECT 127.215 130.525 127.735 131.065 ;
        RECT 115.490 129.775 120.835 130.320 ;
        RECT 121.010 129.775 126.355 130.320 ;
        RECT 126.525 129.775 127.735 130.525 ;
        RECT 14.660 129.605 127.820 129.775 ;
        RECT 14.745 128.855 15.955 129.605 ;
        RECT 17.855 129.145 18.140 129.605 ;
        RECT 19.270 129.125 19.930 129.605 ;
        RECT 21.540 129.145 21.860 129.605 ;
        RECT 22.600 129.165 23.010 129.605 ;
        RECT 24.835 129.225 25.165 129.605 ;
        RECT 25.775 129.225 26.105 129.605 ;
        RECT 26.705 128.855 27.915 129.605 ;
        RECT 28.090 129.060 33.435 129.605 ;
        RECT 14.745 128.315 15.265 128.855 ;
        RECT 27.395 128.315 27.915 128.855 ;
        RECT 31.510 128.230 31.850 129.060 ;
        RECT 33.645 128.785 33.875 129.605 ;
        RECT 34.545 128.785 34.755 129.605 ;
        RECT 36.135 129.145 36.385 129.605 ;
        RECT 37.285 128.880 37.575 129.605 ;
        RECT 38.205 128.835 40.795 129.605 ;
        RECT 40.970 129.060 46.315 129.605 ;
        RECT 47.635 129.145 47.885 129.605 ;
        RECT 49.250 129.060 54.595 129.605 ;
        RECT 55.505 129.070 56.015 129.605 ;
        RECT 57.975 129.205 58.305 129.605 ;
        RECT 59.345 129.225 59.675 129.605 ;
        RECT 39.585 128.315 40.795 128.835 ;
        RECT 44.390 128.230 44.730 129.060 ;
        RECT 52.670 128.230 53.010 129.060 ;
        RECT 60.285 128.835 62.875 129.605 ;
        RECT 63.045 128.880 63.335 129.605 ;
        RECT 63.505 128.855 64.715 129.605 ;
        RECT 65.695 129.145 65.980 129.605 ;
        RECT 67.110 129.125 67.770 129.605 ;
        RECT 69.380 129.145 69.700 129.605 ;
        RECT 70.440 129.165 70.850 129.605 ;
        RECT 72.675 129.225 73.005 129.605 ;
        RECT 73.615 129.225 73.945 129.605 ;
        RECT 75.695 129.145 75.945 129.605 ;
        RECT 77.995 129.145 78.245 129.605 ;
        RECT 79.885 129.070 80.395 129.605 ;
        RECT 82.355 129.205 82.685 129.605 ;
        RECT 84.015 129.145 84.265 129.605 ;
        RECT 61.665 128.315 62.875 128.835 ;
        RECT 64.195 128.315 64.715 128.855 ;
        RECT 86.045 128.835 88.635 129.605 ;
        RECT 88.805 128.880 89.095 129.605 ;
        RECT 90.535 129.145 90.820 129.605 ;
        RECT 91.950 129.125 92.610 129.605 ;
        RECT 94.220 129.145 94.540 129.605 ;
        RECT 95.280 129.165 95.690 129.605 ;
        RECT 97.515 129.225 97.845 129.605 ;
        RECT 98.455 129.225 98.785 129.605 ;
        RECT 100.535 129.145 100.785 129.605 ;
        RECT 101.685 128.835 104.275 129.605 ;
        RECT 105.175 129.145 105.425 129.605 ;
        RECT 107.475 129.145 107.725 129.605 ;
        RECT 109.775 129.145 110.025 129.605 ;
        RECT 111.865 129.125 112.145 129.605 ;
        RECT 112.750 129.125 113.005 129.605 ;
        RECT 113.650 129.125 113.925 129.605 ;
        RECT 114.565 128.880 114.855 129.605 ;
        RECT 115.755 129.145 116.005 129.605 ;
        RECT 87.425 128.315 88.635 128.835 ;
        RECT 103.065 128.315 104.275 128.835 ;
        RECT 118.285 128.785 118.515 129.605 ;
        RECT 119.185 128.785 119.395 129.605 ;
        RECT 120.525 129.225 120.855 129.605 ;
        RECT 121.465 128.855 122.675 129.605 ;
        RECT 122.155 128.315 122.675 128.855 ;
        RECT 122.845 128.835 126.355 129.605 ;
        RECT 126.525 128.855 127.735 129.605 ;
        RECT 124.705 128.315 126.355 128.835 ;
        RECT 127.215 128.315 127.735 128.855 ;
        RECT 14.745 125.085 15.265 125.625 ;
        RECT 18.905 125.105 20.555 125.625 ;
        RECT 14.745 124.335 15.955 125.085 ;
        RECT 17.045 124.335 20.555 125.105 ;
        RECT 20.785 124.335 20.995 125.155 ;
        RECT 21.665 124.335 21.895 125.155 ;
        RECT 25.555 125.085 26.075 125.625 ;
        RECT 31.765 125.105 32.975 125.625 ;
        RECT 66.745 125.105 68.395 125.625 ;
        RECT 23.465 124.335 23.795 124.715 ;
        RECT 24.405 124.335 24.695 125.060 ;
        RECT 24.865 124.335 26.075 125.085 ;
        RECT 26.675 124.335 27.005 124.735 ;
        RECT 28.965 124.335 29.475 124.870 ;
        RECT 30.385 124.335 32.975 125.105 ;
        RECT 33.885 124.335 34.395 124.870 ;
        RECT 36.355 124.335 36.685 124.735 ;
        RECT 38.435 124.335 38.685 124.795 ;
        RECT 41.655 124.335 41.905 124.795 ;
        RECT 43.955 124.335 44.205 124.795 ;
        RECT 45.835 124.335 46.085 124.795 ;
        RECT 47.465 124.335 47.745 124.815 ;
        RECT 48.350 124.335 48.605 124.815 ;
        RECT 49.250 124.335 49.525 124.815 ;
        RECT 50.165 124.335 50.455 125.060 ;
        RECT 51.085 124.335 51.390 124.845 ;
        RECT 51.990 124.335 52.250 124.860 ;
        RECT 52.850 124.335 53.110 124.895 ;
        RECT 53.710 124.335 53.970 124.815 ;
        RECT 54.570 124.335 54.830 124.815 ;
        RECT 55.430 124.335 55.675 124.815 ;
        RECT 56.290 124.335 56.535 124.815 ;
        RECT 57.145 124.335 57.395 124.815 ;
        RECT 58.005 124.335 58.255 124.815 ;
        RECT 58.865 124.335 59.125 124.815 ;
        RECT 59.725 124.335 60.025 124.815 ;
        RECT 61.025 124.335 61.535 124.870 ;
        RECT 63.495 124.335 63.825 124.735 ;
        RECT 64.885 124.335 68.395 125.105 ;
        RECT 68.625 124.335 68.835 125.155 ;
        RECT 69.505 124.335 69.735 125.155 ;
        RECT 72.015 125.085 72.535 125.625 ;
        RECT 99.865 125.105 101.515 125.625 ;
        RECT 70.385 124.335 70.715 124.715 ;
        RECT 71.325 124.335 72.535 125.085 ;
        RECT 73.175 124.335 73.450 124.815 ;
        RECT 74.095 124.335 74.350 124.815 ;
        RECT 74.955 124.335 75.235 124.815 ;
        RECT 75.925 124.335 76.215 125.060 ;
        RECT 77.195 124.335 77.480 124.795 ;
        RECT 78.610 124.335 79.270 124.815 ;
        RECT 80.880 124.335 81.200 124.795 ;
        RECT 81.940 124.335 82.350 124.775 ;
        RECT 84.175 124.335 84.505 124.715 ;
        RECT 85.115 124.335 85.445 124.715 ;
        RECT 86.155 124.335 86.325 124.815 ;
        RECT 86.995 124.335 87.165 124.815 ;
        RECT 87.835 124.335 88.005 124.815 ;
        RECT 88.675 124.335 88.845 124.815 ;
        RECT 89.515 124.335 89.685 124.815 ;
        RECT 90.355 124.335 90.525 124.815 ;
        RECT 91.195 124.335 91.365 124.815 ;
        RECT 92.035 124.335 92.205 124.815 ;
        RECT 92.875 124.335 93.045 124.815 ;
        RECT 93.715 124.335 93.885 124.815 ;
        RECT 94.555 124.335 94.725 124.815 ;
        RECT 95.395 124.335 95.565 124.815 ;
        RECT 96.235 124.335 96.405 124.815 ;
        RECT 98.005 124.335 101.515 125.105 ;
        RECT 102.835 125.085 103.355 125.625 ;
        RECT 105.385 125.105 107.035 125.625 ;
        RECT 101.685 124.335 101.975 125.060 ;
        RECT 102.145 124.335 103.355 125.085 ;
        RECT 103.525 124.335 107.035 125.105 ;
        RECT 125.835 125.085 126.355 125.625 ;
        RECT 127.215 125.085 127.735 125.625 ;
        RECT 107.945 124.335 108.455 124.870 ;
        RECT 110.415 124.335 110.745 124.735 ;
        RECT 112.085 124.335 112.595 124.870 ;
        RECT 114.555 124.335 114.885 124.735 ;
        RECT 116.295 124.335 116.580 124.795 ;
        RECT 117.710 124.335 118.370 124.815 ;
        RECT 119.980 124.335 120.300 124.795 ;
        RECT 121.040 124.335 121.450 124.775 ;
        RECT 123.275 124.335 123.605 124.715 ;
        RECT 124.215 124.335 124.545 124.715 ;
        RECT 125.145 124.335 126.355 125.085 ;
        RECT 126.525 124.335 127.735 125.085 ;
        RECT 14.660 124.165 127.820 124.335 ;
        RECT 14.745 123.415 15.955 124.165 ;
        RECT 17.045 123.655 17.350 124.165 ;
        RECT 17.950 123.640 18.210 124.165 ;
        RECT 18.810 123.605 19.070 124.165 ;
        RECT 19.670 123.685 19.930 124.165 ;
        RECT 20.530 123.685 20.790 124.165 ;
        RECT 21.390 123.685 21.635 124.165 ;
        RECT 22.250 123.685 22.495 124.165 ;
        RECT 23.105 123.685 23.355 124.165 ;
        RECT 23.965 123.685 24.215 124.165 ;
        RECT 24.825 123.685 25.085 124.165 ;
        RECT 25.685 123.685 25.985 124.165 ;
        RECT 14.745 122.875 15.265 123.415 ;
        RECT 26.245 123.395 27.915 124.165 ;
        RECT 28.175 123.685 28.475 124.165 ;
        RECT 29.075 123.685 29.335 124.165 ;
        RECT 29.945 123.685 30.195 124.165 ;
        RECT 30.805 123.685 31.055 124.165 ;
        RECT 31.665 123.685 31.910 124.165 ;
        RECT 32.525 123.685 32.770 124.165 ;
        RECT 33.370 123.685 33.630 124.165 ;
        RECT 34.230 123.685 34.490 124.165 ;
        RECT 35.090 123.605 35.350 124.165 ;
        RECT 35.950 123.640 36.210 124.165 ;
        RECT 36.810 123.655 37.115 124.165 ;
        RECT 37.285 123.440 37.575 124.165 ;
        RECT 38.485 123.630 38.995 124.165 ;
        RECT 40.955 123.765 41.285 124.165 ;
        RECT 41.890 123.620 47.235 124.165 ;
        RECT 47.410 123.620 52.755 124.165 ;
        RECT 53.735 123.705 54.020 124.165 ;
        RECT 55.150 123.685 55.810 124.165 ;
        RECT 57.420 123.705 57.740 124.165 ;
        RECT 58.480 123.725 58.890 124.165 ;
        RECT 60.715 123.785 61.045 124.165 ;
        RECT 61.655 123.785 61.985 124.165 ;
        RECT 27.165 122.875 27.915 123.395 ;
        RECT 45.310 122.790 45.650 123.620 ;
        RECT 50.830 122.790 51.170 123.620 ;
        RECT 63.045 123.440 63.335 124.165 ;
        RECT 64.245 123.630 64.755 124.165 ;
        RECT 66.715 123.765 67.045 124.165 ;
        RECT 67.645 123.395 70.235 124.165 ;
        RECT 70.410 123.620 75.755 124.165 ;
        RECT 75.930 123.620 81.275 124.165 ;
        RECT 69.025 122.875 70.235 123.395 ;
        RECT 73.830 122.790 74.170 123.620 ;
        RECT 79.350 122.790 79.690 123.620 ;
        RECT 81.505 123.345 81.715 124.165 ;
        RECT 82.385 123.345 82.615 124.165 ;
        RECT 83.725 123.785 84.055 124.165 ;
        RECT 85.125 123.395 88.635 124.165 ;
        RECT 88.805 123.440 89.095 124.165 ;
        RECT 89.265 123.655 89.570 124.165 ;
        RECT 90.170 123.640 90.430 124.165 ;
        RECT 91.030 123.605 91.290 124.165 ;
        RECT 91.890 123.685 92.150 124.165 ;
        RECT 92.750 123.685 93.010 124.165 ;
        RECT 93.610 123.685 93.855 124.165 ;
        RECT 94.470 123.685 94.715 124.165 ;
        RECT 95.325 123.685 95.575 124.165 ;
        RECT 96.185 123.685 96.435 124.165 ;
        RECT 97.045 123.685 97.305 124.165 ;
        RECT 97.905 123.685 98.205 124.165 ;
        RECT 98.465 123.415 99.675 124.165 ;
        RECT 99.850 123.620 105.195 124.165 ;
        RECT 105.365 123.655 105.670 124.165 ;
        RECT 106.270 123.640 106.530 124.165 ;
        RECT 86.985 122.875 88.635 123.395 ;
        RECT 99.155 122.875 99.675 123.415 ;
        RECT 103.270 122.790 103.610 123.620 ;
        RECT 107.130 123.605 107.390 124.165 ;
        RECT 107.990 123.685 108.250 124.165 ;
        RECT 108.850 123.685 109.110 124.165 ;
        RECT 109.710 123.685 109.955 124.165 ;
        RECT 110.570 123.685 110.815 124.165 ;
        RECT 111.425 123.685 111.675 124.165 ;
        RECT 112.285 123.685 112.535 124.165 ;
        RECT 113.145 123.685 113.405 124.165 ;
        RECT 114.005 123.685 114.305 124.165 ;
        RECT 114.565 123.440 114.855 124.165 ;
        RECT 116.295 123.705 116.580 124.165 ;
        RECT 117.710 123.685 118.370 124.165 ;
        RECT 119.980 123.705 120.300 124.165 ;
        RECT 121.040 123.725 121.450 124.165 ;
        RECT 123.275 123.785 123.605 124.165 ;
        RECT 124.215 123.785 124.545 124.165 ;
        RECT 125.145 123.415 126.355 124.165 ;
        RECT 126.525 123.415 127.735 124.165 ;
        RECT 125.835 122.875 126.355 123.415 ;
        RECT 127.215 122.875 127.735 123.415 ;
        RECT 14.745 119.645 15.265 120.185 ;
        RECT 18.445 119.665 20.095 120.185 ;
        RECT 28.545 119.665 29.295 120.185 ;
        RECT 14.745 118.895 15.955 119.645 ;
        RECT 16.585 118.895 20.095 119.665 ;
        RECT 21.005 118.895 21.515 119.430 ;
        RECT 23.475 118.895 23.805 119.295 ;
        RECT 24.405 118.895 24.695 119.620 ;
        RECT 26.225 118.895 26.555 119.275 ;
        RECT 27.625 118.895 29.295 119.665 ;
        RECT 29.505 118.895 29.735 119.715 ;
        RECT 30.405 118.895 30.615 119.715 ;
        RECT 30.885 118.895 31.115 119.715 ;
        RECT 31.785 118.895 31.995 119.715 ;
        RECT 33.035 118.895 33.320 119.355 ;
        RECT 34.450 118.895 35.110 119.375 ;
        RECT 36.720 118.895 37.040 119.355 ;
        RECT 37.780 118.895 38.190 119.335 ;
        RECT 40.015 118.895 40.345 119.275 ;
        RECT 40.955 118.895 41.285 119.275 ;
        RECT 42.625 118.895 43.135 119.430 ;
        RECT 45.095 118.895 45.425 119.295 ;
        RECT 46.765 118.895 47.275 119.430 ;
        RECT 49.235 118.895 49.565 119.295 ;
        RECT 50.165 118.895 50.455 119.620 ;
        RECT 50.665 118.895 50.895 119.715 ;
        RECT 51.565 118.895 51.775 119.715 ;
        RECT 52.695 119.645 53.215 120.185 ;
        RECT 52.005 118.895 53.215 119.645 ;
        RECT 53.535 118.895 53.865 119.695 ;
        RECT 72.725 119.665 74.375 120.185 ;
        RECT 54.375 118.895 54.705 119.375 ;
        RECT 55.295 118.895 55.535 119.375 ;
        RECT 57.275 118.895 57.605 119.585 ;
        RECT 58.855 118.895 59.185 119.385 ;
        RECT 60.175 118.895 60.460 119.355 ;
        RECT 61.590 118.895 62.250 119.375 ;
        RECT 63.860 118.895 64.180 119.355 ;
        RECT 64.920 118.895 65.330 119.335 ;
        RECT 67.155 118.895 67.485 119.275 ;
        RECT 68.095 118.895 68.425 119.275 ;
        RECT 69.465 118.895 69.795 119.275 ;
        RECT 70.865 118.895 74.375 119.665 ;
        RECT 74.585 118.895 74.815 119.715 ;
        RECT 75.485 118.895 75.695 119.715 ;
        RECT 75.925 118.895 76.215 119.620 ;
        RECT 77.585 118.895 78.095 119.430 ;
        RECT 80.055 118.895 80.385 119.295 ;
        RECT 81.425 118.895 81.755 119.275 ;
        RECT 82.425 118.895 82.635 119.715 ;
        RECT 83.305 118.895 83.535 119.715 ;
        RECT 87.445 119.665 89.095 120.185 ;
        RECT 84.645 118.895 84.975 119.275 ;
        RECT 85.585 118.895 89.095 119.665 ;
        RECT 89.305 118.895 89.535 119.715 ;
        RECT 90.205 118.895 90.415 119.715 ;
        RECT 90.685 118.895 90.915 119.715 ;
        RECT 91.585 118.895 91.795 119.715 ;
        RECT 92.835 118.895 93.120 119.355 ;
        RECT 94.250 118.895 94.910 119.375 ;
        RECT 96.520 118.895 96.840 119.355 ;
        RECT 97.580 118.895 97.990 119.335 ;
        RECT 99.815 118.895 100.145 119.275 ;
        RECT 100.755 118.895 101.085 119.275 ;
        RECT 101.685 118.895 101.975 119.620 ;
        RECT 102.585 118.895 102.915 119.275 ;
        RECT 103.565 118.895 103.795 119.715 ;
        RECT 104.465 118.895 104.675 119.715 ;
        RECT 105.645 118.895 106.155 119.430 ;
        RECT 108.115 118.895 108.445 119.295 ;
        RECT 109.855 118.895 110.140 119.355 ;
        RECT 111.270 118.895 111.930 119.375 ;
        RECT 113.540 118.895 113.860 119.355 ;
        RECT 114.600 118.895 115.010 119.335 ;
        RECT 116.835 118.895 117.165 119.275 ;
        RECT 117.775 118.895 118.105 119.275 ;
        RECT 118.745 118.895 118.975 119.715 ;
        RECT 119.645 118.895 119.855 119.715 ;
        RECT 124.705 119.665 126.355 120.185 ;
        RECT 120.985 118.895 121.315 119.275 ;
        RECT 122.845 118.895 126.355 119.665 ;
        RECT 127.215 119.645 127.735 120.185 ;
        RECT 126.525 118.895 127.735 119.645 ;
        RECT 14.660 118.725 127.820 118.895 ;
        RECT 14.745 117.975 15.955 118.725 ;
        RECT 14.745 117.435 15.265 117.975 ;
        RECT 16.125 117.955 17.795 118.725 ;
        RECT 18.775 118.265 19.060 118.725 ;
        RECT 20.190 118.245 20.850 118.725 ;
        RECT 22.460 118.265 22.780 118.725 ;
        RECT 23.520 118.285 23.930 118.725 ;
        RECT 25.755 118.345 26.085 118.725 ;
        RECT 26.695 118.345 27.025 118.725 ;
        RECT 28.435 118.265 28.720 118.725 ;
        RECT 29.850 118.245 30.510 118.725 ;
        RECT 32.120 118.265 32.440 118.725 ;
        RECT 33.180 118.285 33.590 118.725 ;
        RECT 35.415 118.345 35.745 118.725 ;
        RECT 36.355 118.345 36.685 118.725 ;
        RECT 37.285 118.000 37.575 118.725 ;
        RECT 38.555 118.265 38.840 118.725 ;
        RECT 39.970 118.245 40.630 118.725 ;
        RECT 42.240 118.265 42.560 118.725 ;
        RECT 43.300 118.285 43.710 118.725 ;
        RECT 45.535 118.345 45.865 118.725 ;
        RECT 46.475 118.345 46.805 118.725 ;
        RECT 48.215 118.265 48.500 118.725 ;
        RECT 49.630 118.245 50.290 118.725 ;
        RECT 51.900 118.265 52.220 118.725 ;
        RECT 52.960 118.285 53.370 118.725 ;
        RECT 55.195 118.345 55.525 118.725 ;
        RECT 56.135 118.345 56.465 118.725 ;
        RECT 17.045 117.435 17.795 117.955 ;
        RECT 57.125 117.905 57.335 118.725 ;
        RECT 58.005 117.905 58.235 118.725 ;
        RECT 58.905 117.955 61.495 118.725 ;
        RECT 60.285 117.435 61.495 117.955 ;
        RECT 61.705 117.905 61.935 118.725 ;
        RECT 62.605 117.905 62.815 118.725 ;
        RECT 63.045 118.000 63.335 118.725 ;
        RECT 64.315 118.265 64.600 118.725 ;
        RECT 65.730 118.245 66.390 118.725 ;
        RECT 68.000 118.265 68.320 118.725 ;
        RECT 69.060 118.285 69.470 118.725 ;
        RECT 71.295 118.345 71.625 118.725 ;
        RECT 72.235 118.345 72.565 118.725 ;
        RECT 73.975 118.265 74.260 118.725 ;
        RECT 75.390 118.245 76.050 118.725 ;
        RECT 77.660 118.265 77.980 118.725 ;
        RECT 78.720 118.285 79.130 118.725 ;
        RECT 80.955 118.345 81.285 118.725 ;
        RECT 81.895 118.345 82.225 118.725 ;
        RECT 83.255 118.325 83.585 118.725 ;
        RECT 85.545 118.190 86.055 118.725 ;
        RECT 87.465 117.905 87.695 118.725 ;
        RECT 88.365 117.905 88.575 118.725 ;
        RECT 88.805 118.000 89.095 118.725 ;
        RECT 90.075 118.265 90.360 118.725 ;
        RECT 91.490 118.245 92.150 118.725 ;
        RECT 93.760 118.265 94.080 118.725 ;
        RECT 94.820 118.285 95.230 118.725 ;
        RECT 97.055 118.345 97.385 118.725 ;
        RECT 97.995 118.345 98.325 118.725 ;
        RECT 99.365 118.345 99.695 118.725 ;
        RECT 102.035 118.265 102.320 118.725 ;
        RECT 103.450 118.245 104.110 118.725 ;
        RECT 105.720 118.265 106.040 118.725 ;
        RECT 106.780 118.285 107.190 118.725 ;
        RECT 109.015 118.345 109.345 118.725 ;
        RECT 109.955 118.345 110.285 118.725 ;
        RECT 111.325 118.345 111.655 118.725 ;
        RECT 112.785 117.905 112.995 118.725 ;
        RECT 113.665 117.905 113.895 118.725 ;
        RECT 114.565 118.000 114.855 118.725 ;
        RECT 115.925 118.345 116.255 118.725 ;
        RECT 117.325 118.215 117.630 118.725 ;
        RECT 118.230 118.200 118.490 118.725 ;
        RECT 119.090 118.165 119.350 118.725 ;
        RECT 119.950 118.245 120.210 118.725 ;
        RECT 120.810 118.245 121.070 118.725 ;
        RECT 121.670 118.245 121.915 118.725 ;
        RECT 122.530 118.245 122.775 118.725 ;
        RECT 123.385 118.245 123.635 118.725 ;
        RECT 124.245 118.245 124.495 118.725 ;
        RECT 125.105 118.245 125.365 118.725 ;
        RECT 125.965 118.245 126.265 118.725 ;
        RECT 126.525 117.975 127.735 118.725 ;
        RECT 127.215 117.435 127.735 117.975 ;
        RECT 14.745 114.205 15.265 114.745 ;
        RECT 18.445 114.225 20.095 114.745 ;
        RECT 14.745 113.455 15.955 114.205 ;
        RECT 16.585 113.455 20.095 114.225 ;
        RECT 20.305 113.455 20.535 114.275 ;
        RECT 21.205 113.455 21.415 114.275 ;
        RECT 21.705 113.455 21.915 114.275 ;
        RECT 22.585 113.455 22.815 114.275 ;
        RECT 23.465 113.455 23.795 113.835 ;
        RECT 24.405 113.455 24.695 114.180 ;
        RECT 24.865 113.455 25.170 113.965 ;
        RECT 25.770 113.455 26.030 113.980 ;
        RECT 26.630 113.455 26.890 114.015 ;
        RECT 27.490 113.455 27.750 113.935 ;
        RECT 28.350 113.455 28.610 113.935 ;
        RECT 29.210 113.455 29.455 113.935 ;
        RECT 30.070 113.455 30.315 113.935 ;
        RECT 30.925 113.455 31.175 113.935 ;
        RECT 31.785 113.455 32.035 113.935 ;
        RECT 32.645 113.455 32.905 113.935 ;
        RECT 33.505 113.455 33.805 113.935 ;
        RECT 34.155 113.455 34.455 113.935 ;
        RECT 35.055 113.455 35.315 113.935 ;
        RECT 35.925 113.455 36.175 113.935 ;
        RECT 36.785 113.455 37.035 113.935 ;
        RECT 37.645 113.455 37.890 113.935 ;
        RECT 38.505 113.455 38.750 113.935 ;
        RECT 39.350 113.455 39.610 113.935 ;
        RECT 40.210 113.455 40.470 113.935 ;
        RECT 41.070 113.455 41.330 114.015 ;
        RECT 41.930 113.455 42.190 113.980 ;
        RECT 42.790 113.455 43.095 113.965 ;
        RECT 43.705 113.455 44.035 113.835 ;
        RECT 44.705 113.455 44.915 114.275 ;
        RECT 45.585 113.455 45.815 114.275 ;
        RECT 46.945 114.225 47.695 114.745 ;
        RECT 51.545 114.225 52.295 114.745 ;
        RECT 46.025 113.455 47.695 114.225 ;
        RECT 48.305 113.455 48.635 113.835 ;
        RECT 50.165 113.455 50.455 114.180 ;
        RECT 50.625 113.455 52.295 114.225 ;
        RECT 58.190 114.000 58.530 114.830 ;
        RECT 63.710 114.000 64.050 114.830 ;
        RECT 52.905 113.455 53.235 113.835 ;
        RECT 54.770 113.455 60.115 114.000 ;
        RECT 60.290 113.455 65.635 114.000 ;
        RECT 65.845 113.455 66.075 114.275 ;
        RECT 66.745 113.455 66.955 114.275 ;
        RECT 73.830 114.000 74.170 114.830 ;
        RECT 89.285 114.225 90.935 114.745 ;
        RECT 96.625 114.225 97.375 114.745 ;
        RECT 104.005 114.225 105.655 114.745 ;
        RECT 68.545 113.455 68.875 113.835 ;
        RECT 70.410 113.455 75.755 114.000 ;
        RECT 75.925 113.455 76.215 114.180 ;
        RECT 78.115 113.455 78.400 113.915 ;
        RECT 79.530 113.455 80.190 113.935 ;
        RECT 81.800 113.455 82.120 113.915 ;
        RECT 82.860 113.455 83.270 113.895 ;
        RECT 85.095 113.455 85.425 113.835 ;
        RECT 86.035 113.455 86.365 113.835 ;
        RECT 87.425 113.455 90.935 114.225 ;
        RECT 91.845 113.455 92.355 113.990 ;
        RECT 94.315 113.455 94.645 113.855 ;
        RECT 95.705 113.455 97.375 114.225 ;
        RECT 98.285 113.455 98.795 113.990 ;
        RECT 100.755 113.455 101.085 113.855 ;
        RECT 101.685 113.455 101.975 114.180 ;
        RECT 102.145 113.455 105.655 114.225 ;
        RECT 109.250 114.000 109.590 114.830 ;
        RECT 116.405 114.225 117.155 114.745 ;
        RECT 105.830 113.455 111.175 114.000 ;
        RECT 112.085 113.455 112.595 113.990 ;
        RECT 114.555 113.455 114.885 113.855 ;
        RECT 115.485 113.455 117.155 114.225 ;
        RECT 127.215 114.205 127.735 114.745 ;
        RECT 117.755 113.455 118.085 113.835 ;
        RECT 118.785 113.455 119.115 113.815 ;
        RECT 121.715 113.455 122.045 113.915 ;
        RECT 123.945 113.455 124.135 113.895 ;
        RECT 125.620 113.455 125.925 113.915 ;
        RECT 126.525 113.455 127.735 114.205 ;
        RECT 14.660 113.285 127.820 113.455 ;
        RECT 14.745 112.535 15.955 113.285 ;
        RECT 17.855 112.825 18.140 113.285 ;
        RECT 19.270 112.805 19.930 113.285 ;
        RECT 21.540 112.825 21.860 113.285 ;
        RECT 22.600 112.845 23.010 113.285 ;
        RECT 24.835 112.905 25.165 113.285 ;
        RECT 25.775 112.905 26.105 113.285 ;
        RECT 27.135 112.905 27.465 113.285 ;
        RECT 28.165 112.925 28.495 113.285 ;
        RECT 31.095 112.825 31.425 113.285 ;
        RECT 33.325 112.845 33.515 113.285 ;
        RECT 35.000 112.825 35.305 113.285 ;
        RECT 36.345 112.905 36.675 113.285 ;
        RECT 37.285 112.560 37.575 113.285 ;
        RECT 37.745 112.775 38.050 113.285 ;
        RECT 38.650 112.760 38.910 113.285 ;
        RECT 39.510 112.725 39.770 113.285 ;
        RECT 40.370 112.805 40.630 113.285 ;
        RECT 41.230 112.805 41.490 113.285 ;
        RECT 42.090 112.805 42.335 113.285 ;
        RECT 42.950 112.805 43.195 113.285 ;
        RECT 43.805 112.805 44.055 113.285 ;
        RECT 44.665 112.805 44.915 113.285 ;
        RECT 45.525 112.805 45.785 113.285 ;
        RECT 46.385 112.805 46.685 113.285 ;
        RECT 46.945 112.535 48.155 113.285 ;
        RECT 14.745 111.995 15.265 112.535 ;
        RECT 47.635 111.995 48.155 112.535 ;
        RECT 48.325 112.515 51.835 113.285 ;
        RECT 52.010 112.740 57.355 113.285 ;
        RECT 57.530 112.740 62.875 113.285 ;
        RECT 50.185 111.995 51.835 112.515 ;
        RECT 55.430 111.910 55.770 112.740 ;
        RECT 60.950 111.910 61.290 112.740 ;
        RECT 63.045 112.560 63.335 113.285 ;
        RECT 64.425 112.515 67.935 113.285 ;
        RECT 68.110 112.740 73.455 113.285 ;
        RECT 73.630 112.740 78.975 113.285 ;
        RECT 66.285 111.995 67.935 112.515 ;
        RECT 71.530 111.910 71.870 112.740 ;
        RECT 77.050 111.910 77.390 112.740 ;
        RECT 79.185 112.465 79.415 113.285 ;
        RECT 80.085 112.465 80.295 113.285 ;
        RECT 80.675 112.485 81.005 113.285 ;
        RECT 81.515 112.805 81.845 113.285 ;
        RECT 82.435 112.805 82.675 113.285 ;
        RECT 83.290 112.740 88.635 113.285 ;
        RECT 86.710 111.910 87.050 112.740 ;
        RECT 88.805 112.560 89.095 113.285 ;
        RECT 89.725 112.515 93.235 113.285 ;
        RECT 91.585 111.995 93.235 112.515 ;
        RECT 93.465 112.465 93.675 113.285 ;
        RECT 94.345 112.465 94.575 113.285 ;
        RECT 95.250 112.740 100.595 113.285 ;
        RECT 100.770 112.740 106.115 113.285 ;
        RECT 106.725 112.905 107.055 113.285 ;
        RECT 98.670 111.910 99.010 112.740 ;
        RECT 104.190 111.910 104.530 112.740 ;
        RECT 107.665 112.535 108.875 113.285 ;
        RECT 109.050 112.740 114.395 113.285 ;
        RECT 108.355 111.995 108.875 112.535 ;
        RECT 112.470 111.910 112.810 112.740 ;
        RECT 114.565 112.560 114.855 113.285 ;
        RECT 115.115 112.805 115.415 113.285 ;
        RECT 116.015 112.805 116.275 113.285 ;
        RECT 116.885 112.805 117.135 113.285 ;
        RECT 117.745 112.805 117.995 113.285 ;
        RECT 118.605 112.805 118.850 113.285 ;
        RECT 119.465 112.805 119.710 113.285 ;
        RECT 120.310 112.805 120.570 113.285 ;
        RECT 121.170 112.805 121.430 113.285 ;
        RECT 122.030 112.725 122.290 113.285 ;
        RECT 122.890 112.760 123.150 113.285 ;
        RECT 123.750 112.775 124.055 113.285 ;
        RECT 124.665 112.905 124.995 113.285 ;
        RECT 126.525 112.535 127.735 113.285 ;
        RECT 127.215 111.995 127.735 112.535 ;
        RECT 14.745 108.765 15.265 109.305 ;
        RECT 16.815 108.765 17.335 109.305 ;
        RECT 14.745 108.015 15.955 108.765 ;
        RECT 16.125 108.015 17.335 108.765 ;
        RECT 20.930 108.560 21.270 109.390 ;
        RECT 17.510 108.015 22.855 108.560 ;
        RECT 23.065 108.015 23.295 108.835 ;
        RECT 23.965 108.015 24.175 108.835 ;
        RECT 25.555 108.765 26.075 109.305 ;
        RECT 49.475 108.765 49.995 109.305 ;
        RECT 55.245 108.785 56.895 109.305 ;
        RECT 59.365 108.785 60.115 109.305 ;
        RECT 24.405 108.015 24.695 108.740 ;
        RECT 24.865 108.015 26.075 108.765 ;
        RECT 26.685 108.015 27.015 108.395 ;
        RECT 28.065 108.015 28.395 108.395 ;
        RECT 29.005 108.015 29.310 108.525 ;
        RECT 29.910 108.015 30.170 108.540 ;
        RECT 30.770 108.015 31.030 108.575 ;
        RECT 31.630 108.015 31.890 108.495 ;
        RECT 32.490 108.015 32.750 108.495 ;
        RECT 33.350 108.015 33.595 108.495 ;
        RECT 34.210 108.015 34.455 108.495 ;
        RECT 35.065 108.015 35.315 108.495 ;
        RECT 35.925 108.015 36.175 108.495 ;
        RECT 36.785 108.015 37.045 108.495 ;
        RECT 37.645 108.015 37.945 108.495 ;
        RECT 38.635 108.015 38.965 108.395 ;
        RECT 39.665 108.015 39.995 108.375 ;
        RECT 42.595 108.015 42.925 108.475 ;
        RECT 44.825 108.015 45.015 108.455 ;
        RECT 46.500 108.015 46.805 108.475 ;
        RECT 47.845 108.015 48.175 108.395 ;
        RECT 48.785 108.015 49.995 108.765 ;
        RECT 50.165 108.015 50.455 108.740 ;
        RECT 51.525 108.015 51.855 108.395 ;
        RECT 53.385 108.015 56.895 108.785 ;
        RECT 57.505 108.015 57.835 108.395 ;
        RECT 58.445 108.015 60.115 108.785 ;
        RECT 60.725 108.015 60.965 108.495 ;
        RECT 61.555 108.015 61.885 108.495 ;
        RECT 62.395 108.015 62.725 108.815 ;
        RECT 63.945 108.015 64.275 108.395 ;
        RECT 64.975 108.015 65.275 108.495 ;
        RECT 65.875 108.015 66.135 108.495 ;
        RECT 66.745 108.015 66.995 108.495 ;
        RECT 67.605 108.015 67.855 108.495 ;
        RECT 68.465 108.015 68.710 108.495 ;
        RECT 69.325 108.015 69.570 108.495 ;
        RECT 70.170 108.015 70.430 108.495 ;
        RECT 71.030 108.015 71.290 108.495 ;
        RECT 71.890 108.015 72.150 108.575 ;
        RECT 72.750 108.015 73.010 108.540 ;
        RECT 73.610 108.015 73.915 108.525 ;
        RECT 74.605 108.015 74.815 108.835 ;
        RECT 75.485 108.015 75.715 108.835 ;
        RECT 75.925 108.015 76.215 108.740 ;
        RECT 76.935 108.015 77.235 108.495 ;
        RECT 77.835 108.015 78.095 108.495 ;
        RECT 78.705 108.015 78.955 108.495 ;
        RECT 79.565 108.015 79.815 108.495 ;
        RECT 80.425 108.015 80.670 108.495 ;
        RECT 81.285 108.015 81.530 108.495 ;
        RECT 82.130 108.015 82.390 108.495 ;
        RECT 82.990 108.015 83.250 108.495 ;
        RECT 83.850 108.015 84.110 108.575 ;
        RECT 84.710 108.015 84.970 108.540 ;
        RECT 85.570 108.015 85.875 108.525 ;
        RECT 86.085 108.015 86.315 108.835 ;
        RECT 86.985 108.015 87.195 108.835 ;
        RECT 87.865 108.015 88.195 108.395 ;
        RECT 88.895 108.015 89.195 108.495 ;
        RECT 89.795 108.015 90.055 108.495 ;
        RECT 90.665 108.015 90.915 108.495 ;
        RECT 91.525 108.015 91.775 108.495 ;
        RECT 92.385 108.015 92.630 108.495 ;
        RECT 93.245 108.015 93.490 108.495 ;
        RECT 94.090 108.015 94.350 108.495 ;
        RECT 94.950 108.015 95.210 108.495 ;
        RECT 95.810 108.015 96.070 108.575 ;
        RECT 96.670 108.015 96.930 108.540 ;
        RECT 97.530 108.015 97.835 108.525 ;
        RECT 98.965 108.015 99.195 108.835 ;
        RECT 99.865 108.015 100.075 108.835 ;
        RECT 100.745 108.015 101.075 108.395 ;
        RECT 101.685 108.015 101.975 108.740 ;
        RECT 102.235 108.015 102.535 108.495 ;
        RECT 103.135 108.015 103.395 108.495 ;
        RECT 104.005 108.015 104.255 108.495 ;
        RECT 104.865 108.015 105.115 108.495 ;
        RECT 105.725 108.015 105.970 108.495 ;
        RECT 106.585 108.015 106.830 108.495 ;
        RECT 107.430 108.015 107.690 108.495 ;
        RECT 108.290 108.015 108.550 108.495 ;
        RECT 109.150 108.015 109.410 108.575 ;
        RECT 110.010 108.015 110.270 108.540 ;
        RECT 110.870 108.015 111.175 108.525 ;
        RECT 111.785 108.015 112.115 108.395 ;
        RECT 113.165 108.015 113.495 108.395 ;
        RECT 115.005 108.015 115.335 108.395 ;
        RECT 115.985 108.015 116.215 108.835 ;
        RECT 116.885 108.015 117.095 108.835 ;
        RECT 127.215 108.765 127.735 109.305 ;
        RECT 117.755 108.015 118.060 108.475 ;
        RECT 119.545 108.015 119.735 108.455 ;
        RECT 121.635 108.015 121.965 108.475 ;
        RECT 124.565 108.015 124.895 108.375 ;
        RECT 125.595 108.015 125.925 108.395 ;
        RECT 126.525 108.015 127.735 108.765 ;
        RECT 14.660 107.845 127.820 108.015 ;
        RECT 14.745 107.095 15.955 107.845 ;
        RECT 16.125 107.095 17.335 107.845 ;
        RECT 14.745 106.555 15.265 107.095 ;
        RECT 16.815 106.555 17.335 107.095 ;
        RECT 17.565 107.025 17.775 107.845 ;
        RECT 18.445 107.025 18.675 107.845 ;
        RECT 19.315 107.385 19.620 107.845 ;
        RECT 21.105 107.405 21.295 107.845 ;
        RECT 23.195 107.385 23.525 107.845 ;
        RECT 26.125 107.485 26.455 107.845 ;
        RECT 27.155 107.465 27.485 107.845 ;
        RECT 28.515 107.385 28.820 107.845 ;
        RECT 30.305 107.405 30.495 107.845 ;
        RECT 32.395 107.385 32.725 107.845 ;
        RECT 35.325 107.485 35.655 107.845 ;
        RECT 36.355 107.465 36.685 107.845 ;
        RECT 37.285 107.120 37.575 107.845 ;
        RECT 37.785 107.025 38.015 107.845 ;
        RECT 38.685 107.025 38.895 107.845 ;
        RECT 39.215 107.365 39.515 107.845 ;
        RECT 40.115 107.365 40.375 107.845 ;
        RECT 40.985 107.365 41.235 107.845 ;
        RECT 41.845 107.365 42.095 107.845 ;
        RECT 42.705 107.365 42.950 107.845 ;
        RECT 43.565 107.365 43.810 107.845 ;
        RECT 44.410 107.365 44.670 107.845 ;
        RECT 45.270 107.365 45.530 107.845 ;
        RECT 46.130 107.285 46.390 107.845 ;
        RECT 46.990 107.320 47.250 107.845 ;
        RECT 47.850 107.335 48.155 107.845 ;
        RECT 48.755 107.385 49.060 107.845 ;
        RECT 50.545 107.405 50.735 107.845 ;
        RECT 52.635 107.385 52.965 107.845 ;
        RECT 55.565 107.485 55.895 107.845 ;
        RECT 56.595 107.465 56.925 107.845 ;
        RECT 57.585 107.025 57.795 107.845 ;
        RECT 58.465 107.025 58.695 107.845 ;
        RECT 58.905 107.095 60.115 107.845 ;
        RECT 59.595 106.555 60.115 107.095 ;
        RECT 60.325 107.025 60.555 107.845 ;
        RECT 61.225 107.025 61.435 107.845 ;
        RECT 62.105 107.465 62.435 107.845 ;
        RECT 63.045 107.120 63.335 107.845 ;
        RECT 63.545 107.025 63.775 107.845 ;
        RECT 64.445 107.025 64.655 107.845 ;
        RECT 65.315 107.385 65.620 107.845 ;
        RECT 67.105 107.405 67.295 107.845 ;
        RECT 69.195 107.385 69.525 107.845 ;
        RECT 72.125 107.485 72.455 107.845 ;
        RECT 73.155 107.465 73.485 107.845 ;
        RECT 75.065 107.025 75.275 107.845 ;
        RECT 75.945 107.025 76.175 107.845 ;
        RECT 76.825 107.465 77.155 107.845 ;
        RECT 78.195 107.385 78.500 107.845 ;
        RECT 79.985 107.405 80.175 107.845 ;
        RECT 82.075 107.385 82.405 107.845 ;
        RECT 85.005 107.485 85.335 107.845 ;
        RECT 86.035 107.465 86.365 107.845 ;
        RECT 87.405 107.465 87.735 107.845 ;
        RECT 88.805 107.120 89.095 107.845 ;
        RECT 90.615 107.385 90.920 107.845 ;
        RECT 92.405 107.405 92.595 107.845 ;
        RECT 94.495 107.385 94.825 107.845 ;
        RECT 97.425 107.485 97.755 107.845 ;
        RECT 98.455 107.465 98.785 107.845 ;
        RECT 99.815 107.385 100.120 107.845 ;
        RECT 101.605 107.405 101.795 107.845 ;
        RECT 103.695 107.385 104.025 107.845 ;
        RECT 106.625 107.485 106.955 107.845 ;
        RECT 107.655 107.465 107.985 107.845 ;
        RECT 108.645 107.025 108.855 107.845 ;
        RECT 109.525 107.025 109.755 107.845 ;
        RECT 110.005 107.025 110.235 107.845 ;
        RECT 110.905 107.025 111.115 107.845 ;
        RECT 111.345 107.075 113.015 107.845 ;
        RECT 112.265 106.555 113.015 107.075 ;
        RECT 113.225 107.025 113.455 107.845 ;
        RECT 114.125 107.025 114.335 107.845 ;
        RECT 114.565 107.120 114.855 107.845 ;
        RECT 115.455 107.385 115.760 107.845 ;
        RECT 117.245 107.405 117.435 107.845 ;
        RECT 119.335 107.385 119.665 107.845 ;
        RECT 122.265 107.485 122.595 107.845 ;
        RECT 123.295 107.465 123.625 107.845 ;
        RECT 124.265 107.025 124.495 107.845 ;
        RECT 125.165 107.025 125.375 107.845 ;
        RECT 126.525 107.095 127.735 107.845 ;
        RECT 127.215 106.555 127.735 107.095 ;
        RECT 14.745 103.325 15.265 103.865 ;
        RECT 17.505 103.345 18.715 103.865 ;
        RECT 14.745 102.575 15.955 103.325 ;
        RECT 16.125 102.575 18.715 103.345 ;
        RECT 22.310 103.120 22.650 103.950 ;
        RECT 25.555 103.325 26.075 103.865 ;
        RECT 18.890 102.575 24.235 103.120 ;
        RECT 24.405 102.575 24.695 103.300 ;
        RECT 24.865 102.575 26.075 103.325 ;
        RECT 26.305 102.575 26.515 103.395 ;
        RECT 27.185 102.575 27.415 103.395 ;
        RECT 27.665 102.575 27.895 103.395 ;
        RECT 28.565 102.575 28.775 103.395 ;
        RECT 29.445 102.575 29.775 102.955 ;
        RECT 30.825 102.575 31.155 102.955 ;
        RECT 32.195 102.575 32.500 103.035 ;
        RECT 33.985 102.575 34.175 103.015 ;
        RECT 36.075 102.575 36.405 103.035 ;
        RECT 39.005 102.575 39.335 102.935 ;
        RECT 40.035 102.575 40.365 102.955 ;
        RECT 41.395 102.575 41.700 103.035 ;
        RECT 43.185 102.575 43.375 103.015 ;
        RECT 45.275 102.575 45.605 103.035 ;
        RECT 48.205 102.575 48.535 102.935 ;
        RECT 49.235 102.575 49.565 102.955 ;
        RECT 50.165 102.575 50.455 103.300 ;
        RECT 51.605 102.575 51.815 103.395 ;
        RECT 52.485 102.575 52.715 103.395 ;
        RECT 53.615 103.325 54.135 103.865 ;
        RECT 74.545 103.345 75.755 103.865 ;
        RECT 52.925 102.575 54.135 103.325 ;
        RECT 54.735 102.575 55.040 103.035 ;
        RECT 56.525 102.575 56.715 103.015 ;
        RECT 58.615 102.575 58.945 103.035 ;
        RECT 61.545 102.575 61.875 102.935 ;
        RECT 62.575 102.575 62.905 102.955 ;
        RECT 63.935 102.575 64.240 103.035 ;
        RECT 65.725 102.575 65.915 103.015 ;
        RECT 67.815 102.575 68.145 103.035 ;
        RECT 70.745 102.575 71.075 102.935 ;
        RECT 71.775 102.575 72.105 102.955 ;
        RECT 73.165 102.575 75.755 103.345 ;
        RECT 75.925 102.575 76.215 103.300 ;
        RECT 99.590 103.120 99.930 103.950 ;
        RECT 123.325 103.345 124.975 103.865 ;
        RECT 76.815 102.575 77.120 103.035 ;
        RECT 78.605 102.575 78.795 103.015 ;
        RECT 80.695 102.575 81.025 103.035 ;
        RECT 83.625 102.575 83.955 102.935 ;
        RECT 84.655 102.575 84.985 102.955 ;
        RECT 86.015 102.575 86.320 103.035 ;
        RECT 87.805 102.575 87.995 103.015 ;
        RECT 89.895 102.575 90.225 103.035 ;
        RECT 92.825 102.575 93.155 102.935 ;
        RECT 93.855 102.575 94.185 102.955 ;
        RECT 95.225 102.575 95.555 102.955 ;
        RECT 96.170 102.575 101.515 103.120 ;
        RECT 101.685 102.575 101.975 103.300 ;
        RECT 102.575 102.575 102.905 102.955 ;
        RECT 103.605 102.575 103.935 102.935 ;
        RECT 106.535 102.575 106.865 103.035 ;
        RECT 108.765 102.575 108.955 103.015 ;
        RECT 110.440 102.575 110.745 103.035 ;
        RECT 111.775 102.575 112.080 103.035 ;
        RECT 113.565 102.575 113.755 103.015 ;
        RECT 115.655 102.575 115.985 103.035 ;
        RECT 118.585 102.575 118.915 102.935 ;
        RECT 119.615 102.575 119.945 102.955 ;
        RECT 121.465 102.575 124.975 103.345 ;
        RECT 127.215 103.325 127.735 103.865 ;
        RECT 125.585 102.575 125.915 102.955 ;
        RECT 126.525 102.575 127.735 103.325 ;
        RECT 14.660 102.405 127.820 102.575 ;
        RECT 14.745 101.655 15.955 102.405 ;
        RECT 14.745 101.115 15.265 101.655 ;
        RECT 16.125 101.635 18.715 102.405 ;
        RECT 18.890 101.860 24.235 102.405 ;
        RECT 17.505 101.115 18.715 101.635 ;
        RECT 22.310 101.030 22.650 101.860 ;
        RECT 24.405 101.680 24.695 102.405 ;
        RECT 25.325 101.635 27.915 102.405 ;
        RECT 28.175 101.925 28.475 102.405 ;
        RECT 29.075 101.925 29.335 102.405 ;
        RECT 29.945 101.925 30.195 102.405 ;
        RECT 30.805 101.925 31.055 102.405 ;
        RECT 31.665 101.925 31.910 102.405 ;
        RECT 32.525 101.925 32.770 102.405 ;
        RECT 33.370 101.925 33.630 102.405 ;
        RECT 34.230 101.925 34.490 102.405 ;
        RECT 35.090 101.845 35.350 102.405 ;
        RECT 35.950 101.880 36.210 102.405 ;
        RECT 36.810 101.895 37.115 102.405 ;
        RECT 37.285 101.680 37.575 102.405 ;
        RECT 26.705 101.115 27.915 101.635 ;
        RECT 38.265 101.585 38.475 102.405 ;
        RECT 39.145 101.585 39.375 102.405 ;
        RECT 40.025 102.025 40.355 102.405 ;
        RECT 41.055 101.925 41.355 102.405 ;
        RECT 41.955 101.925 42.215 102.405 ;
        RECT 42.825 101.925 43.075 102.405 ;
        RECT 43.685 101.925 43.935 102.405 ;
        RECT 44.545 101.925 44.790 102.405 ;
        RECT 45.405 101.925 45.650 102.405 ;
        RECT 46.250 101.925 46.510 102.405 ;
        RECT 47.110 101.925 47.370 102.405 ;
        RECT 47.970 101.845 48.230 102.405 ;
        RECT 48.830 101.880 49.090 102.405 ;
        RECT 49.690 101.895 49.995 102.405 ;
        RECT 50.165 101.680 50.455 102.405 ;
        RECT 51.085 101.635 52.755 102.405 ;
        RECT 53.015 101.925 53.315 102.405 ;
        RECT 53.915 101.925 54.175 102.405 ;
        RECT 54.785 101.925 55.035 102.405 ;
        RECT 55.645 101.925 55.895 102.405 ;
        RECT 56.505 101.925 56.750 102.405 ;
        RECT 57.365 101.925 57.610 102.405 ;
        RECT 58.210 101.925 58.470 102.405 ;
        RECT 59.070 101.925 59.330 102.405 ;
        RECT 59.930 101.845 60.190 102.405 ;
        RECT 60.790 101.880 61.050 102.405 ;
        RECT 61.650 101.895 61.955 102.405 ;
        RECT 63.045 101.680 63.335 102.405 ;
        RECT 63.505 101.895 63.810 102.405 ;
        RECT 64.410 101.880 64.670 102.405 ;
        RECT 65.270 101.845 65.530 102.405 ;
        RECT 66.130 101.925 66.390 102.405 ;
        RECT 66.990 101.925 67.250 102.405 ;
        RECT 67.850 101.925 68.095 102.405 ;
        RECT 68.710 101.925 68.955 102.405 ;
        RECT 69.565 101.925 69.815 102.405 ;
        RECT 70.425 101.925 70.675 102.405 ;
        RECT 71.285 101.925 71.545 102.405 ;
        RECT 72.145 101.925 72.445 102.405 ;
        RECT 73.165 101.635 75.755 102.405 ;
        RECT 75.925 101.680 76.215 102.405 ;
        RECT 76.385 101.895 76.690 102.405 ;
        RECT 77.290 101.880 77.550 102.405 ;
        RECT 78.150 101.845 78.410 102.405 ;
        RECT 79.010 101.925 79.270 102.405 ;
        RECT 79.870 101.925 80.130 102.405 ;
        RECT 80.730 101.925 80.975 102.405 ;
        RECT 81.590 101.925 81.835 102.405 ;
        RECT 82.445 101.925 82.695 102.405 ;
        RECT 83.305 101.925 83.555 102.405 ;
        RECT 84.165 101.925 84.425 102.405 ;
        RECT 85.025 101.925 85.325 102.405 ;
        RECT 86.045 101.635 88.635 102.405 ;
        RECT 88.805 101.680 89.095 102.405 ;
        RECT 89.265 101.895 89.570 102.405 ;
        RECT 90.170 101.880 90.430 102.405 ;
        RECT 91.030 101.845 91.290 102.405 ;
        RECT 91.890 101.925 92.150 102.405 ;
        RECT 92.750 101.925 93.010 102.405 ;
        RECT 93.610 101.925 93.855 102.405 ;
        RECT 94.470 101.925 94.715 102.405 ;
        RECT 95.325 101.925 95.575 102.405 ;
        RECT 96.185 101.925 96.435 102.405 ;
        RECT 97.045 101.925 97.305 102.405 ;
        RECT 97.905 101.925 98.205 102.405 ;
        RECT 98.925 101.635 101.515 102.405 ;
        RECT 101.685 101.680 101.975 102.405 ;
        RECT 102.235 101.925 102.535 102.405 ;
        RECT 103.135 101.925 103.395 102.405 ;
        RECT 104.005 101.925 104.255 102.405 ;
        RECT 104.865 101.925 105.115 102.405 ;
        RECT 105.725 101.925 105.970 102.405 ;
        RECT 106.585 101.925 106.830 102.405 ;
        RECT 107.430 101.925 107.690 102.405 ;
        RECT 108.290 101.925 108.550 102.405 ;
        RECT 109.150 101.845 109.410 102.405 ;
        RECT 110.010 101.880 110.270 102.405 ;
        RECT 110.870 101.895 111.175 102.405 ;
        RECT 111.805 101.635 114.395 102.405 ;
        RECT 114.565 101.680 114.855 102.405 ;
        RECT 115.025 101.895 115.330 102.405 ;
        RECT 115.930 101.880 116.190 102.405 ;
        RECT 116.790 101.845 117.050 102.405 ;
        RECT 117.650 101.925 117.910 102.405 ;
        RECT 118.510 101.925 118.770 102.405 ;
        RECT 119.370 101.925 119.615 102.405 ;
        RECT 120.230 101.925 120.475 102.405 ;
        RECT 121.085 101.925 121.335 102.405 ;
        RECT 121.945 101.925 122.195 102.405 ;
        RECT 122.805 101.925 123.065 102.405 ;
        RECT 123.665 101.925 123.965 102.405 ;
        RECT 124.685 101.635 126.355 102.405 ;
        RECT 126.525 101.655 127.735 102.405 ;
        RECT 52.005 101.115 52.755 101.635 ;
        RECT 74.545 101.115 75.755 101.635 ;
        RECT 87.425 101.115 88.635 101.635 ;
        RECT 100.305 101.115 101.515 101.635 ;
        RECT 113.185 101.115 114.395 101.635 ;
        RECT 125.605 101.115 126.355 101.635 ;
        RECT 127.215 101.115 127.735 101.655 ;
        RECT 19.135 48.040 23.045 48.260 ;
        RECT 19.135 45.640 20.855 48.040 ;
        RECT 21.255 46.320 21.425 47.360 ;
        RECT 22.615 45.640 23.045 48.040 ;
        RECT 19.135 45.370 23.045 45.640 ;
        RECT 30.335 48.050 34.245 48.270 ;
        RECT 30.335 45.650 32.055 48.050 ;
        RECT 32.455 46.330 32.625 47.370 ;
        RECT 33.815 45.650 34.245 48.050 ;
        RECT 30.335 45.380 34.245 45.650 ;
        RECT 41.555 48.020 45.465 48.240 ;
        RECT 41.555 45.620 43.275 48.020 ;
        RECT 43.675 46.300 43.845 47.340 ;
        RECT 45.035 45.620 45.465 48.020 ;
        RECT 41.555 45.350 45.465 45.620 ;
        RECT 52.805 48.000 56.715 48.220 ;
        RECT 52.805 45.600 54.525 48.000 ;
        RECT 54.925 46.280 55.095 47.320 ;
        RECT 56.285 45.600 56.715 48.000 ;
        RECT 52.805 45.330 56.715 45.600 ;
        RECT 64.025 47.990 67.935 48.210 ;
        RECT 64.025 45.590 65.745 47.990 ;
        RECT 66.145 46.270 66.315 47.310 ;
        RECT 67.505 45.590 67.935 47.990 ;
        RECT 64.025 45.320 67.935 45.590 ;
        RECT 75.265 47.980 79.175 48.200 ;
        RECT 75.265 45.580 76.985 47.980 ;
        RECT 77.385 46.260 77.555 47.300 ;
        RECT 78.745 45.580 79.175 47.980 ;
        RECT 75.265 45.310 79.175 45.580 ;
        RECT 86.515 47.990 90.425 48.210 ;
        RECT 86.515 45.590 88.235 47.990 ;
        RECT 88.635 46.270 88.805 47.310 ;
        RECT 89.995 45.590 90.425 47.990 ;
        RECT 86.515 45.320 90.425 45.590 ;
        RECT 97.795 47.980 101.705 48.200 ;
        RECT 97.795 45.580 99.515 47.980 ;
        RECT 99.915 46.260 100.085 47.300 ;
        RECT 101.275 45.580 101.705 47.980 ;
        RECT 97.795 45.310 101.705 45.580 ;
        RECT 109.065 47.980 112.975 48.200 ;
        RECT 109.065 45.580 110.785 47.980 ;
        RECT 111.185 46.260 111.355 47.300 ;
        RECT 112.545 45.580 112.975 47.980 ;
        RECT 109.065 45.310 112.975 45.580 ;
        RECT 120.315 47.980 124.225 48.200 ;
        RECT 120.315 45.580 122.035 47.980 ;
        RECT 122.435 46.260 122.605 47.300 ;
        RECT 123.795 45.580 124.225 47.980 ;
        RECT 120.315 45.310 124.225 45.580 ;
        RECT 25.695 39.770 29.605 40.040 ;
        RECT 25.695 37.370 26.125 39.770 ;
        RECT 27.315 38.050 27.485 39.090 ;
        RECT 27.885 37.370 29.605 39.770 ;
        RECT 25.695 37.150 29.605 37.370 ;
        RECT 36.975 39.770 40.885 40.040 ;
        RECT 36.975 37.370 37.405 39.770 ;
        RECT 38.595 38.050 38.765 39.090 ;
        RECT 39.165 37.370 40.885 39.770 ;
        RECT 36.975 37.150 40.885 37.370 ;
        RECT 48.265 39.750 52.175 40.020 ;
        RECT 48.265 37.350 48.695 39.750 ;
        RECT 49.885 38.030 50.055 39.070 ;
        RECT 50.455 37.350 52.175 39.750 ;
        RECT 48.265 37.130 52.175 37.350 ;
        RECT 59.485 39.750 63.395 40.020 ;
        RECT 59.485 37.350 59.915 39.750 ;
        RECT 61.105 38.030 61.275 39.070 ;
        RECT 61.675 37.350 63.395 39.750 ;
        RECT 59.485 37.130 63.395 37.350 ;
        RECT 70.685 39.750 74.595 40.020 ;
        RECT 70.685 37.350 71.115 39.750 ;
        RECT 72.305 38.030 72.475 39.070 ;
        RECT 72.875 37.350 74.595 39.750 ;
        RECT 70.685 37.130 74.595 37.350 ;
        RECT 81.975 39.740 85.885 40.010 ;
        RECT 81.975 37.340 82.405 39.740 ;
        RECT 83.595 38.020 83.765 39.060 ;
        RECT 84.165 37.340 85.885 39.740 ;
        RECT 81.975 37.120 85.885 37.340 ;
        RECT 93.215 39.760 97.125 40.030 ;
        RECT 93.215 37.360 93.645 39.760 ;
        RECT 94.835 38.040 95.005 39.080 ;
        RECT 95.405 37.360 97.125 39.760 ;
        RECT 93.215 37.140 97.125 37.360 ;
        RECT 104.425 39.780 108.335 40.050 ;
        RECT 104.425 37.380 104.855 39.780 ;
        RECT 106.045 38.060 106.215 39.100 ;
        RECT 106.615 37.380 108.335 39.780 ;
        RECT 104.425 37.160 108.335 37.380 ;
        RECT 115.625 39.820 119.535 40.090 ;
        RECT 115.625 37.420 116.055 39.820 ;
        RECT 117.245 38.100 117.415 39.140 ;
        RECT 117.815 37.420 119.535 39.820 ;
        RECT 115.625 37.200 119.535 37.420 ;
        RECT 126.835 39.840 130.745 40.110 ;
        RECT 126.835 37.440 127.265 39.840 ;
        RECT 128.455 38.120 128.625 39.160 ;
        RECT 129.025 37.440 130.745 39.840 ;
        RECT 126.835 37.220 130.745 37.440 ;
      LAYER met1 ;
        RECT 14.660 211.050 127.820 211.530 ;
        RECT 14.660 205.610 127.820 206.090 ;
        RECT 14.660 200.170 127.820 200.650 ;
        RECT 14.660 194.730 127.820 195.210 ;
        RECT 14.660 189.290 127.820 189.770 ;
        RECT 14.660 183.850 127.820 184.330 ;
        RECT 14.660 178.410 127.820 178.890 ;
        RECT 14.660 172.970 127.820 173.450 ;
        RECT 14.660 167.530 127.820 168.010 ;
        RECT 14.660 162.090 127.820 162.570 ;
        RECT 14.660 156.650 127.820 157.130 ;
        RECT 14.660 151.210 127.820 151.690 ;
        RECT 14.660 145.770 127.820 146.250 ;
        RECT 14.660 140.330 127.820 140.810 ;
        RECT 14.660 134.890 127.820 135.370 ;
        RECT 14.660 129.450 127.820 129.930 ;
        RECT 14.660 124.010 127.820 124.490 ;
        RECT 14.660 118.570 127.820 119.050 ;
        RECT 14.660 113.130 127.820 113.610 ;
        RECT 14.660 107.690 127.820 108.170 ;
        RECT 14.660 102.250 127.820 102.730 ;
        RECT 133.330 76.630 136.060 77.830 ;
        RECT 3.910 73.080 6.100 73.190 ;
        RECT 3.910 72.820 12.240 73.080 ;
        RECT 29.635 72.840 43.235 72.850 ;
        RECT 18.435 72.820 43.235 72.840 ;
        RECT 3.910 72.800 54.455 72.820 ;
        RECT 3.910 72.790 65.705 72.800 ;
        RECT 133.960 72.790 135.640 76.630 ;
        RECT 3.910 72.780 76.925 72.790 ;
        RECT 85.815 72.780 99.415 72.790 ;
        RECT 132.085 72.780 140.600 72.790 ;
        RECT 3.910 71.700 140.600 72.780 ;
        RECT 3.910 71.690 32.035 71.700 ;
        RECT 3.910 71.670 19.135 71.690 ;
        RECT 40.855 71.670 140.600 71.700 ;
        RECT 3.910 71.500 12.240 71.670 ;
        RECT 52.105 71.650 140.600 71.670 ;
        RECT 63.325 71.640 140.600 71.650 ;
        RECT 74.565 71.630 88.165 71.640 ;
        RECT 97.095 71.630 133.215 71.640 ;
        RECT 3.910 71.370 6.100 71.500 ;
        RECT 10.800 71.180 11.950 71.500 ;
        RECT 10.800 69.480 11.915 71.180 ;
        RECT 10.800 13.800 11.950 69.480 ;
        RECT 19.295 46.650 20.065 47.720 ;
        RECT 21.225 47.200 21.455 47.340 ;
        RECT 21.085 46.430 21.475 47.200 ;
        RECT 30.495 46.660 31.265 47.730 ;
        RECT 32.425 47.210 32.655 47.350 ;
        RECT 32.285 46.440 32.675 47.210 ;
        RECT 41.715 46.630 42.485 47.700 ;
        RECT 43.645 47.180 43.875 47.320 ;
        RECT 21.225 46.340 21.455 46.430 ;
        RECT 32.425 46.350 32.655 46.440 ;
        RECT 43.505 46.410 43.895 47.180 ;
        RECT 52.965 46.610 53.735 47.680 ;
        RECT 54.895 47.160 55.125 47.300 ;
        RECT 43.645 46.320 43.875 46.410 ;
        RECT 54.755 46.390 55.145 47.160 ;
        RECT 64.185 46.600 64.955 47.670 ;
        RECT 66.115 47.150 66.345 47.290 ;
        RECT 54.895 46.300 55.125 46.390 ;
        RECT 65.975 46.380 66.365 47.150 ;
        RECT 75.425 46.590 76.195 47.660 ;
        RECT 77.355 47.140 77.585 47.280 ;
        RECT 66.115 46.290 66.345 46.380 ;
        RECT 77.215 46.370 77.605 47.140 ;
        RECT 86.675 46.600 87.445 47.670 ;
        RECT 88.605 47.150 88.835 47.290 ;
        RECT 88.465 46.380 88.855 47.150 ;
        RECT 97.955 46.590 98.725 47.660 ;
        RECT 99.885 47.140 100.115 47.280 ;
        RECT 77.355 46.280 77.585 46.370 ;
        RECT 88.605 46.290 88.835 46.380 ;
        RECT 99.745 46.370 100.135 47.140 ;
        RECT 109.225 46.590 109.995 47.660 ;
        RECT 111.155 47.140 111.385 47.280 ;
        RECT 111.015 46.370 111.405 47.140 ;
        RECT 120.475 46.590 121.245 47.660 ;
        RECT 122.405 47.140 122.635 47.280 ;
        RECT 122.265 46.370 122.655 47.140 ;
        RECT 99.885 46.280 100.115 46.370 ;
        RECT 111.155 46.280 111.385 46.370 ;
        RECT 122.405 46.280 122.635 46.370 ;
        RECT 27.285 38.980 27.515 39.070 ;
        RECT 38.565 38.980 38.795 39.070 ;
        RECT 27.265 38.210 27.655 38.980 ;
        RECT 27.285 38.070 27.515 38.210 ;
        RECT 28.675 37.690 29.445 38.760 ;
        RECT 38.545 38.210 38.935 38.980 ;
        RECT 49.855 38.960 50.085 39.050 ;
        RECT 61.075 38.960 61.305 39.050 ;
        RECT 72.275 38.960 72.505 39.050 ;
        RECT 38.565 38.070 38.795 38.210 ;
        RECT 39.955 37.690 40.725 38.760 ;
        RECT 49.835 38.190 50.225 38.960 ;
        RECT 49.855 38.050 50.085 38.190 ;
        RECT 51.245 37.670 52.015 38.740 ;
        RECT 61.055 38.190 61.445 38.960 ;
        RECT 61.075 38.050 61.305 38.190 ;
        RECT 62.465 37.670 63.235 38.740 ;
        RECT 72.255 38.190 72.645 38.960 ;
        RECT 83.565 38.950 83.795 39.040 ;
        RECT 94.805 38.970 95.035 39.060 ;
        RECT 106.015 38.990 106.245 39.080 ;
        RECT 117.215 39.030 117.445 39.120 ;
        RECT 128.425 39.050 128.655 39.140 ;
        RECT 72.275 38.050 72.505 38.190 ;
        RECT 73.665 37.670 74.435 38.740 ;
        RECT 83.545 38.180 83.935 38.950 ;
        RECT 83.565 38.040 83.795 38.180 ;
        RECT 84.955 37.660 85.725 38.730 ;
        RECT 94.785 38.200 95.175 38.970 ;
        RECT 94.805 38.060 95.035 38.200 ;
        RECT 96.195 37.680 96.965 38.750 ;
        RECT 105.995 38.220 106.385 38.990 ;
        RECT 106.015 38.080 106.245 38.220 ;
        RECT 107.405 37.700 108.175 38.770 ;
        RECT 117.195 38.260 117.585 39.030 ;
        RECT 117.215 38.120 117.445 38.260 ;
        RECT 118.605 37.740 119.375 38.810 ;
        RECT 128.405 38.280 128.795 39.050 ;
        RECT 128.425 38.140 128.655 38.280 ;
        RECT 129.815 37.760 130.585 38.830 ;
        RECT 16.965 13.800 17.435 13.810 ;
        RECT 10.800 13.780 17.435 13.800 ;
        RECT 10.800 13.720 17.555 13.780 ;
        RECT 117.845 13.770 131.445 13.790 ;
        RECT 106.635 13.730 131.445 13.770 ;
        RECT 10.800 13.700 41.585 13.720 ;
        RECT 95.435 13.710 131.445 13.730 ;
        RECT 10.800 13.690 75.295 13.700 ;
        RECT 84.225 13.690 131.445 13.710 ;
        RECT 10.800 12.650 131.445 13.690 ;
        RECT 16.705 12.640 131.445 12.650 ;
        RECT 16.705 12.620 120.235 12.640 ;
        RECT 16.705 12.580 109.035 12.620 ;
        RECT 16.705 12.570 97.825 12.580 ;
        RECT 39.275 12.560 97.825 12.570 ;
        RECT 39.275 12.550 86.585 12.560 ;
        RECT 72.985 12.540 86.585 12.550 ;
      LAYER met2 ;
        RECT 28.180 211.105 30.060 211.475 ;
        RECT 58.180 211.105 60.060 211.475 ;
        RECT 88.180 211.105 90.060 211.475 ;
        RECT 118.180 211.105 120.060 211.475 ;
        RECT 28.180 205.665 30.060 206.035 ;
        RECT 58.180 205.665 60.060 206.035 ;
        RECT 88.180 205.665 90.060 206.035 ;
        RECT 118.180 205.665 120.060 206.035 ;
        RECT 28.180 200.225 30.060 200.595 ;
        RECT 58.180 200.225 60.060 200.595 ;
        RECT 88.180 200.225 90.060 200.595 ;
        RECT 118.180 200.225 120.060 200.595 ;
        RECT 28.180 194.785 30.060 195.155 ;
        RECT 58.180 194.785 60.060 195.155 ;
        RECT 88.180 194.785 90.060 195.155 ;
        RECT 118.180 194.785 120.060 195.155 ;
        RECT 28.180 189.345 30.060 189.715 ;
        RECT 58.180 189.345 60.060 189.715 ;
        RECT 88.180 189.345 90.060 189.715 ;
        RECT 118.180 189.345 120.060 189.715 ;
        RECT 28.180 183.905 30.060 184.275 ;
        RECT 58.180 183.905 60.060 184.275 ;
        RECT 88.180 183.905 90.060 184.275 ;
        RECT 118.180 183.905 120.060 184.275 ;
        RECT 28.180 178.465 30.060 178.835 ;
        RECT 58.180 178.465 60.060 178.835 ;
        RECT 88.180 178.465 90.060 178.835 ;
        RECT 118.180 178.465 120.060 178.835 ;
        RECT 28.180 173.025 30.060 173.395 ;
        RECT 58.180 173.025 60.060 173.395 ;
        RECT 88.180 173.025 90.060 173.395 ;
        RECT 118.180 173.025 120.060 173.395 ;
        RECT 28.180 167.585 30.060 167.955 ;
        RECT 58.180 167.585 60.060 167.955 ;
        RECT 88.180 167.585 90.060 167.955 ;
        RECT 118.180 167.585 120.060 167.955 ;
        RECT 28.180 162.145 30.060 162.515 ;
        RECT 58.180 162.145 60.060 162.515 ;
        RECT 88.180 162.145 90.060 162.515 ;
        RECT 118.180 162.145 120.060 162.515 ;
        RECT 28.180 156.705 30.060 157.075 ;
        RECT 58.180 156.705 60.060 157.075 ;
        RECT 88.180 156.705 90.060 157.075 ;
        RECT 118.180 156.705 120.060 157.075 ;
        RECT 28.180 151.265 30.060 151.635 ;
        RECT 58.180 151.265 60.060 151.635 ;
        RECT 88.180 151.265 90.060 151.635 ;
        RECT 118.180 151.265 120.060 151.635 ;
        RECT 28.180 145.825 30.060 146.195 ;
        RECT 58.180 145.825 60.060 146.195 ;
        RECT 88.180 145.825 90.060 146.195 ;
        RECT 118.180 145.825 120.060 146.195 ;
        RECT 28.180 140.385 30.060 140.755 ;
        RECT 58.180 140.385 60.060 140.755 ;
        RECT 88.180 140.385 90.060 140.755 ;
        RECT 118.180 140.385 120.060 140.755 ;
        RECT 28.180 134.945 30.060 135.315 ;
        RECT 58.180 134.945 60.060 135.315 ;
        RECT 88.180 134.945 90.060 135.315 ;
        RECT 118.180 134.945 120.060 135.315 ;
        RECT 28.180 129.505 30.060 129.875 ;
        RECT 58.180 129.505 60.060 129.875 ;
        RECT 88.180 129.505 90.060 129.875 ;
        RECT 118.180 129.505 120.060 129.875 ;
        RECT 28.180 124.065 30.060 124.435 ;
        RECT 58.180 124.065 60.060 124.435 ;
        RECT 88.180 124.065 90.060 124.435 ;
        RECT 118.180 124.065 120.060 124.435 ;
        RECT 28.180 118.625 30.060 118.995 ;
        RECT 58.180 118.625 60.060 118.995 ;
        RECT 88.180 118.625 90.060 118.995 ;
        RECT 118.180 118.625 120.060 118.995 ;
        RECT 28.180 113.185 30.060 113.555 ;
        RECT 58.180 113.185 60.060 113.555 ;
        RECT 88.180 113.185 90.060 113.555 ;
        RECT 118.180 113.185 120.060 113.555 ;
        RECT 28.180 107.745 30.060 108.115 ;
        RECT 58.180 107.745 60.060 108.115 ;
        RECT 88.180 107.745 90.060 108.115 ;
        RECT 118.180 107.745 120.060 108.115 ;
        RECT 28.180 102.305 30.060 102.675 ;
        RECT 58.180 102.305 60.060 102.675 ;
        RECT 88.180 102.305 90.060 102.675 ;
        RECT 118.180 102.305 120.060 102.675 ;
        RECT 133.380 76.580 136.010 77.880 ;
        RECT 3.960 71.320 6.050 73.240 ;
        RECT 19.005 71.800 19.865 72.640 ;
        RECT 30.205 71.810 31.065 72.650 ;
        RECT 19.305 68.570 19.845 71.800 ;
        RECT 30.505 68.580 31.045 71.810 ;
        RECT 41.425 71.780 42.285 72.620 ;
        RECT 19.325 47.770 19.825 68.570 ;
        RECT 30.525 47.780 31.025 68.580 ;
        RECT 41.725 68.550 42.265 71.780 ;
        RECT 52.675 71.760 53.535 72.600 ;
        RECT 19.325 47.060 20.015 47.770 ;
        RECT 21.135 47.060 21.425 47.250 ;
        RECT 19.325 46.620 21.425 47.060 ;
        RECT 19.325 46.600 20.015 46.620 ;
        RECT 21.135 46.380 21.425 46.620 ;
        RECT 30.525 47.070 31.215 47.780 ;
        RECT 41.745 47.750 42.245 68.550 ;
        RECT 52.975 68.530 53.515 71.760 ;
        RECT 63.895 71.750 64.755 72.590 ;
        RECT 32.335 47.070 32.625 47.260 ;
        RECT 30.525 46.630 32.625 47.070 ;
        RECT 30.525 46.610 31.215 46.630 ;
        RECT 32.335 46.390 32.625 46.630 ;
        RECT 41.745 47.040 42.435 47.750 ;
        RECT 52.995 47.730 53.495 68.530 ;
        RECT 64.195 68.520 64.735 71.750 ;
        RECT 75.135 71.740 75.995 72.580 ;
        RECT 86.385 71.750 87.245 72.590 ;
        RECT 43.555 47.040 43.845 47.230 ;
        RECT 41.745 46.600 43.845 47.040 ;
        RECT 41.745 46.580 42.435 46.600 ;
        RECT 43.555 46.360 43.845 46.600 ;
        RECT 52.995 47.020 53.685 47.730 ;
        RECT 64.215 47.720 64.715 68.520 ;
        RECT 75.435 68.510 75.975 71.740 ;
        RECT 86.685 68.520 87.225 71.750 ;
        RECT 97.665 71.740 98.525 72.580 ;
        RECT 108.935 71.740 109.795 72.580 ;
        RECT 120.185 71.740 121.045 72.580 ;
        RECT 54.805 47.020 55.095 47.210 ;
        RECT 52.995 46.580 55.095 47.020 ;
        RECT 52.995 46.560 53.685 46.580 ;
        RECT 54.805 46.340 55.095 46.580 ;
        RECT 64.215 47.010 64.905 47.720 ;
        RECT 75.455 47.710 75.955 68.510 ;
        RECT 86.705 47.720 87.205 68.520 ;
        RECT 97.965 68.510 98.505 71.740 ;
        RECT 109.235 68.510 109.775 71.740 ;
        RECT 120.485 68.510 121.025 71.740 ;
        RECT 66.025 47.010 66.315 47.200 ;
        RECT 64.215 46.570 66.315 47.010 ;
        RECT 64.215 46.550 64.905 46.570 ;
        RECT 66.025 46.330 66.315 46.570 ;
        RECT 75.455 47.000 76.145 47.710 ;
        RECT 77.265 47.000 77.555 47.190 ;
        RECT 75.455 46.560 77.555 47.000 ;
        RECT 75.455 46.540 76.145 46.560 ;
        RECT 77.265 46.320 77.555 46.560 ;
        RECT 86.705 47.010 87.395 47.720 ;
        RECT 97.985 47.710 98.485 68.510 ;
        RECT 109.255 47.710 109.755 68.510 ;
        RECT 120.505 47.710 121.005 68.510 ;
        RECT 88.515 47.010 88.805 47.200 ;
        RECT 86.705 46.570 88.805 47.010 ;
        RECT 86.705 46.550 87.395 46.570 ;
        RECT 88.515 46.330 88.805 46.570 ;
        RECT 97.985 47.000 98.675 47.710 ;
        RECT 99.795 47.000 100.085 47.190 ;
        RECT 97.985 46.560 100.085 47.000 ;
        RECT 97.985 46.540 98.675 46.560 ;
        RECT 99.795 46.320 100.085 46.560 ;
        RECT 109.255 47.000 109.945 47.710 ;
        RECT 111.065 47.000 111.355 47.190 ;
        RECT 109.255 46.560 111.355 47.000 ;
        RECT 109.255 46.540 109.945 46.560 ;
        RECT 111.065 46.320 111.355 46.560 ;
        RECT 120.505 47.000 121.195 47.710 ;
        RECT 122.315 47.000 122.605 47.190 ;
        RECT 120.505 46.560 122.605 47.000 ;
        RECT 120.505 46.540 121.195 46.560 ;
        RECT 122.315 46.320 122.605 46.560 ;
        RECT 27.315 38.790 27.605 39.030 ;
        RECT 28.725 38.790 29.415 38.810 ;
        RECT 27.315 38.350 29.415 38.790 ;
        RECT 27.315 38.160 27.605 38.350 ;
        RECT 28.725 37.640 29.415 38.350 ;
        RECT 38.595 38.790 38.885 39.030 ;
        RECT 40.005 38.790 40.695 38.810 ;
        RECT 38.595 38.350 40.695 38.790 ;
        RECT 38.595 38.160 38.885 38.350 ;
        RECT 40.005 37.640 40.695 38.350 ;
        RECT 49.885 38.770 50.175 39.010 ;
        RECT 51.295 38.770 51.985 38.790 ;
        RECT 49.885 38.330 51.985 38.770 ;
        RECT 49.885 38.140 50.175 38.330 ;
        RECT 28.915 16.840 29.415 37.640 ;
        RECT 40.195 16.840 40.695 37.640 ;
        RECT 51.295 37.620 51.985 38.330 ;
        RECT 61.105 38.770 61.395 39.010 ;
        RECT 62.515 38.770 63.205 38.790 ;
        RECT 61.105 38.330 63.205 38.770 ;
        RECT 61.105 38.140 61.395 38.330 ;
        RECT 62.515 37.620 63.205 38.330 ;
        RECT 72.305 38.770 72.595 39.010 ;
        RECT 73.715 38.770 74.405 38.790 ;
        RECT 72.305 38.330 74.405 38.770 ;
        RECT 72.305 38.140 72.595 38.330 ;
        RECT 73.715 37.620 74.405 38.330 ;
        RECT 83.595 38.760 83.885 39.000 ;
        RECT 94.835 38.780 95.125 39.020 ;
        RECT 106.045 38.800 106.335 39.040 ;
        RECT 117.245 38.840 117.535 39.080 ;
        RECT 128.455 38.860 128.745 39.100 ;
        RECT 129.865 38.860 130.555 38.880 ;
        RECT 118.655 38.840 119.345 38.860 ;
        RECT 107.455 38.800 108.145 38.820 ;
        RECT 96.245 38.780 96.935 38.800 ;
        RECT 85.005 38.760 85.695 38.780 ;
        RECT 83.595 38.320 85.695 38.760 ;
        RECT 83.595 38.130 83.885 38.320 ;
        RECT 28.895 13.610 29.435 16.840 ;
        RECT 40.175 13.610 40.715 16.840 ;
        RECT 51.485 16.820 51.985 37.620 ;
        RECT 62.705 16.820 63.205 37.620 ;
        RECT 73.905 16.820 74.405 37.620 ;
        RECT 85.005 37.610 85.695 38.320 ;
        RECT 94.835 38.340 96.935 38.780 ;
        RECT 94.835 38.150 95.125 38.340 ;
        RECT 96.245 37.630 96.935 38.340 ;
        RECT 106.045 38.360 108.145 38.800 ;
        RECT 106.045 38.170 106.335 38.360 ;
        RECT 107.455 37.650 108.145 38.360 ;
        RECT 117.245 38.400 119.345 38.840 ;
        RECT 117.245 38.210 117.535 38.400 ;
        RECT 118.655 37.690 119.345 38.400 ;
        RECT 128.455 38.420 130.555 38.860 ;
        RECT 128.455 38.230 128.745 38.420 ;
        RECT 129.865 37.710 130.555 38.420 ;
        RECT 28.875 12.770 29.735 13.610 ;
        RECT 40.155 12.770 41.015 13.610 ;
        RECT 51.465 13.590 52.005 16.820 ;
        RECT 62.685 13.590 63.225 16.820 ;
        RECT 73.885 13.590 74.425 16.820 ;
        RECT 85.195 16.810 85.695 37.610 ;
        RECT 96.435 16.830 96.935 37.630 ;
        RECT 107.645 16.850 108.145 37.650 ;
        RECT 118.845 16.890 119.345 37.690 ;
        RECT 130.055 16.910 130.555 37.710 ;
        RECT 51.445 12.750 52.305 13.590 ;
        RECT 62.665 12.750 63.525 13.590 ;
        RECT 73.865 12.750 74.725 13.590 ;
        RECT 85.175 13.580 85.715 16.810 ;
        RECT 96.415 13.600 96.955 16.830 ;
        RECT 107.625 13.620 108.165 16.850 ;
        RECT 118.825 13.660 119.365 16.890 ;
        RECT 130.035 13.680 130.575 16.910 ;
        RECT 85.155 12.740 86.015 13.580 ;
        RECT 96.395 12.760 97.255 13.600 ;
        RECT 107.605 12.780 108.465 13.620 ;
        RECT 118.805 12.820 119.665 13.660 ;
        RECT 130.015 12.840 130.875 13.680 ;
      LAYER met3 ;
        RECT 28.130 211.125 30.110 211.455 ;
        RECT 58.130 211.125 60.110 211.455 ;
        RECT 88.130 211.125 90.110 211.455 ;
        RECT 118.130 211.125 120.110 211.455 ;
        RECT 28.130 205.685 30.110 206.015 ;
        RECT 58.130 205.685 60.110 206.015 ;
        RECT 88.130 205.685 90.110 206.015 ;
        RECT 118.130 205.685 120.110 206.015 ;
        RECT 28.130 200.245 30.110 200.575 ;
        RECT 58.130 200.245 60.110 200.575 ;
        RECT 88.130 200.245 90.110 200.575 ;
        RECT 118.130 200.245 120.110 200.575 ;
        RECT 28.130 194.805 30.110 195.135 ;
        RECT 58.130 194.805 60.110 195.135 ;
        RECT 88.130 194.805 90.110 195.135 ;
        RECT 118.130 194.805 120.110 195.135 ;
        RECT 28.130 189.365 30.110 189.695 ;
        RECT 58.130 189.365 60.110 189.695 ;
        RECT 88.130 189.365 90.110 189.695 ;
        RECT 118.130 189.365 120.110 189.695 ;
        RECT 28.130 183.925 30.110 184.255 ;
        RECT 58.130 183.925 60.110 184.255 ;
        RECT 88.130 183.925 90.110 184.255 ;
        RECT 118.130 183.925 120.110 184.255 ;
        RECT 28.130 178.485 30.110 178.815 ;
        RECT 58.130 178.485 60.110 178.815 ;
        RECT 88.130 178.485 90.110 178.815 ;
        RECT 118.130 178.485 120.110 178.815 ;
        RECT 28.130 173.045 30.110 173.375 ;
        RECT 58.130 173.045 60.110 173.375 ;
        RECT 88.130 173.045 90.110 173.375 ;
        RECT 118.130 173.045 120.110 173.375 ;
        RECT 28.130 167.605 30.110 167.935 ;
        RECT 58.130 167.605 60.110 167.935 ;
        RECT 88.130 167.605 90.110 167.935 ;
        RECT 118.130 167.605 120.110 167.935 ;
        RECT 28.130 162.165 30.110 162.495 ;
        RECT 58.130 162.165 60.110 162.495 ;
        RECT 88.130 162.165 90.110 162.495 ;
        RECT 118.130 162.165 120.110 162.495 ;
        RECT 28.130 156.725 30.110 157.055 ;
        RECT 58.130 156.725 60.110 157.055 ;
        RECT 88.130 156.725 90.110 157.055 ;
        RECT 118.130 156.725 120.110 157.055 ;
        RECT 28.130 151.285 30.110 151.615 ;
        RECT 58.130 151.285 60.110 151.615 ;
        RECT 88.130 151.285 90.110 151.615 ;
        RECT 118.130 151.285 120.110 151.615 ;
        RECT 28.130 145.845 30.110 146.175 ;
        RECT 58.130 145.845 60.110 146.175 ;
        RECT 88.130 145.845 90.110 146.175 ;
        RECT 118.130 145.845 120.110 146.175 ;
        RECT 28.130 140.405 30.110 140.735 ;
        RECT 58.130 140.405 60.110 140.735 ;
        RECT 88.130 140.405 90.110 140.735 ;
        RECT 118.130 140.405 120.110 140.735 ;
        RECT 28.130 134.965 30.110 135.295 ;
        RECT 58.130 134.965 60.110 135.295 ;
        RECT 88.130 134.965 90.110 135.295 ;
        RECT 118.130 134.965 120.110 135.295 ;
        RECT 28.130 129.525 30.110 129.855 ;
        RECT 58.130 129.525 60.110 129.855 ;
        RECT 88.130 129.525 90.110 129.855 ;
        RECT 118.130 129.525 120.110 129.855 ;
        RECT 28.130 124.085 30.110 124.415 ;
        RECT 58.130 124.085 60.110 124.415 ;
        RECT 88.130 124.085 90.110 124.415 ;
        RECT 118.130 124.085 120.110 124.415 ;
        RECT 28.130 118.645 30.110 118.975 ;
        RECT 58.130 118.645 60.110 118.975 ;
        RECT 88.130 118.645 90.110 118.975 ;
        RECT 118.130 118.645 120.110 118.975 ;
        RECT 28.130 113.205 30.110 113.535 ;
        RECT 58.130 113.205 60.110 113.535 ;
        RECT 88.130 113.205 90.110 113.535 ;
        RECT 118.130 113.205 120.110 113.535 ;
        RECT 28.130 107.765 30.110 108.095 ;
        RECT 58.130 107.765 60.110 108.095 ;
        RECT 88.130 107.765 90.110 108.095 ;
        RECT 118.130 107.765 120.110 108.095 ;
        RECT 28.130 102.325 30.110 102.655 ;
        RECT 58.130 102.325 60.110 102.655 ;
        RECT 88.130 102.325 90.110 102.655 ;
        RECT 118.130 102.325 120.110 102.655 ;
        RECT 133.330 76.605 136.060 77.855 ;
        RECT 3.910 71.345 6.100 73.215 ;
      LAYER met4 ;
        RECT 30.670 225.140 30.970 225.760 ;
        RECT 33.430 225.140 33.730 225.760 ;
        RECT 36.190 225.140 36.490 225.760 ;
        RECT 38.950 225.140 39.250 225.760 ;
        RECT 41.710 225.140 42.010 225.760 ;
        RECT 44.470 225.140 44.770 225.760 ;
        RECT 47.230 225.140 47.530 225.760 ;
        RECT 49.990 225.140 50.290 225.760 ;
        RECT 52.750 225.140 53.050 225.760 ;
        RECT 55.510 225.140 55.810 225.760 ;
        RECT 58.270 225.140 58.570 225.760 ;
        RECT 61.030 225.140 61.330 225.760 ;
        RECT 63.790 225.140 64.090 225.760 ;
        RECT 66.550 225.140 66.850 225.760 ;
        RECT 69.310 225.140 69.610 225.760 ;
        RECT 72.070 225.140 72.370 225.760 ;
        RECT 74.830 225.140 75.130 225.760 ;
        RECT 77.590 225.140 77.890 225.760 ;
        RECT 80.350 225.140 80.650 225.760 ;
        RECT 83.110 225.140 83.410 225.760 ;
        RECT 85.870 225.140 86.170 225.760 ;
        RECT 88.630 225.140 88.930 225.760 ;
        RECT 91.390 225.140 91.690 225.760 ;
        RECT 94.150 225.140 94.450 225.760 ;
        RECT 96.910 225.140 97.210 225.760 ;
        RECT 99.670 225.140 99.970 225.760 ;
        RECT 102.430 225.140 102.730 225.760 ;
        RECT 105.190 225.140 105.490 225.760 ;
        RECT 107.950 225.140 108.250 225.760 ;
        RECT 110.710 225.140 111.010 225.760 ;
        RECT 113.470 225.140 113.770 225.760 ;
        RECT 116.230 225.140 116.530 225.760 ;
        RECT 118.990 225.140 119.290 225.760 ;
        RECT 121.750 225.140 122.050 225.760 ;
        RECT 124.510 225.140 124.810 225.760 ;
        RECT 127.270 225.140 127.570 225.760 ;
        RECT 130.030 225.140 130.330 225.760 ;
        RECT 132.790 225.140 133.090 225.760 ;
        RECT 30.420 225.130 133.520 225.140 ;
        RECT 30.300 224.240 133.520 225.130 ;
        RECT 4.000 219.100 6.000 220.760 ;
        RECT 30.300 219.100 31.660 224.240 ;
        RECT 4.000 218.040 31.660 219.100 ;
        RECT 4.000 73.195 6.000 218.040 ;
        RECT 30.300 217.960 31.660 218.040 ;
        RECT 28.120 99.530 30.120 211.530 ;
        RECT 58.120 99.530 60.120 211.530 ;
        RECT 88.120 99.530 90.120 211.530 ;
        RECT 118.120 99.670 120.120 211.530 ;
        RECT 118.110 97.700 120.130 99.670 ;
        RECT 118.130 93.980 120.130 97.700 ;
        RECT 118.130 91.980 135.580 93.980 ;
        RECT 133.580 77.835 135.580 91.980 ;
        RECT 133.375 76.625 136.015 77.835 ;
        RECT 3.955 71.365 6.055 73.195 ;
        RECT 4.000 5.000 6.000 71.365 ;
      LAYER met5 ;
        RECT 14.420 201.590 128.060 203.590 ;
        RECT 14.420 171.590 128.060 173.590 ;
        RECT 14.420 141.590 128.060 143.590 ;
        RECT 14.420 111.590 128.060 113.590 ;
    END
  END vss
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  OBS
      LAYER pwell ;
        RECT 14.805 211.185 14.975 211.375 ;
        RECT 18.485 211.185 18.655 211.375 ;
        RECT 24.005 211.185 24.175 211.375 ;
        RECT 25.845 211.185 26.015 211.375 ;
        RECT 31.365 211.185 31.535 211.375 ;
        RECT 36.885 211.185 37.055 211.375 ;
        RECT 38.725 211.185 38.895 211.375 ;
        RECT 44.245 211.185 44.415 211.375 ;
        RECT 49.765 211.185 49.935 211.375 ;
        RECT 51.605 211.185 51.775 211.375 ;
        RECT 57.125 211.185 57.295 211.375 ;
        RECT 62.645 211.185 62.815 211.375 ;
        RECT 64.485 211.185 64.655 211.375 ;
        RECT 70.005 211.185 70.175 211.375 ;
        RECT 75.525 211.185 75.695 211.375 ;
        RECT 77.365 211.185 77.535 211.375 ;
        RECT 82.885 211.185 83.055 211.375 ;
        RECT 88.405 211.185 88.575 211.375 ;
        RECT 90.245 211.185 90.415 211.375 ;
        RECT 95.765 211.185 95.935 211.375 ;
        RECT 101.285 211.185 101.455 211.375 ;
        RECT 103.125 211.185 103.295 211.375 ;
        RECT 108.645 211.185 108.815 211.375 ;
        RECT 114.165 211.185 114.335 211.375 ;
        RECT 115.140 211.235 115.260 211.345 ;
        RECT 120.605 211.185 120.775 211.375 ;
        RECT 126.125 211.185 126.295 211.375 ;
        RECT 127.505 211.185 127.675 211.375 ;
        RECT 14.665 210.375 16.035 211.185 ;
        RECT 16.045 210.375 18.795 211.185 ;
        RECT 18.805 210.375 24.315 211.185 ;
        RECT 24.785 210.375 26.155 211.185 ;
        RECT 26.165 210.375 31.675 211.185 ;
        RECT 31.685 210.375 37.195 211.185 ;
        RECT 37.665 210.375 39.035 211.185 ;
        RECT 39.045 210.375 44.555 211.185 ;
        RECT 44.565 210.375 50.075 211.185 ;
        RECT 50.545 210.375 51.915 211.185 ;
        RECT 51.925 210.375 57.435 211.185 ;
        RECT 57.445 210.375 62.955 211.185 ;
        RECT 63.425 210.375 64.795 211.185 ;
        RECT 64.805 210.375 70.315 211.185 ;
        RECT 70.325 210.375 75.835 211.185 ;
        RECT 76.305 210.375 77.675 211.185 ;
        RECT 77.685 210.375 83.195 211.185 ;
        RECT 83.205 210.375 88.715 211.185 ;
        RECT 89.185 210.375 90.555 211.185 ;
        RECT 90.565 210.375 96.075 211.185 ;
        RECT 96.085 210.375 101.595 211.185 ;
        RECT 102.065 210.375 103.435 211.185 ;
        RECT 103.445 210.375 108.955 211.185 ;
        RECT 108.965 210.375 114.475 211.185 ;
        RECT 115.405 210.375 120.915 211.185 ;
        RECT 120.925 210.375 126.435 211.185 ;
        RECT 126.445 210.375 127.815 211.185 ;
        RECT 14.665 205.955 16.035 206.765 ;
        RECT 16.045 205.955 18.795 206.765 ;
        RECT 18.805 205.955 24.315 206.765 ;
        RECT 25.245 205.955 27.995 206.765 ;
        RECT 28.005 205.955 33.515 206.765 ;
        RECT 33.525 205.955 39.035 206.765 ;
        RECT 39.045 205.955 44.555 206.765 ;
        RECT 44.565 205.955 50.075 206.765 ;
        RECT 50.545 205.955 52.375 206.765 ;
        RECT 52.385 205.955 57.895 206.765 ;
        RECT 57.905 205.955 63.415 206.765 ;
        RECT 63.425 205.955 68.935 206.765 ;
        RECT 68.945 205.955 74.455 206.765 ;
        RECT 74.475 205.955 75.825 206.865 ;
        RECT 76.305 205.955 77.675 206.765 ;
        RECT 77.685 205.955 80.795 206.865 ;
        RECT 81.365 205.955 85.035 206.765 ;
        RECT 85.045 205.955 90.555 206.765 ;
        RECT 90.565 205.955 96.075 206.765 ;
        RECT 96.085 205.955 101.595 206.765 ;
        RECT 102.525 205.955 104.355 206.765 ;
        RECT 104.365 205.955 109.875 206.765 ;
        RECT 109.885 205.955 115.395 206.765 ;
        RECT 115.405 205.955 120.915 206.765 ;
        RECT 120.925 205.955 126.435 206.765 ;
        RECT 126.445 205.955 127.815 206.765 ;
        RECT 14.805 205.745 14.975 205.955 ;
        RECT 16.645 205.790 16.805 205.900 ;
        RECT 18.485 205.765 18.655 205.955 ;
        RECT 20.325 205.745 20.495 205.935 ;
        RECT 24.005 205.765 24.175 205.955 ;
        RECT 24.980 205.795 25.100 205.905 ;
        RECT 25.845 205.745 26.015 205.935 ;
        RECT 27.685 205.765 27.855 205.955 ;
        RECT 31.365 205.745 31.535 205.935 ;
        RECT 33.205 205.765 33.375 205.955 ;
        RECT 36.885 205.745 37.055 205.935 ;
        RECT 37.860 205.795 37.980 205.905 ;
        RECT 38.725 205.765 38.895 205.955 ;
        RECT 40.565 205.745 40.735 205.935 ;
        RECT 44.245 205.765 44.415 205.955 ;
        RECT 46.085 205.745 46.255 205.935 ;
        RECT 49.765 205.765 49.935 205.955 ;
        RECT 51.605 205.745 51.775 205.935 ;
        RECT 52.065 205.765 52.235 205.955 ;
        RECT 57.125 205.745 57.295 205.935 ;
        RECT 57.585 205.765 57.755 205.955 ;
        RECT 62.645 205.745 62.815 205.935 ;
        RECT 63.105 205.765 63.275 205.955 ;
        RECT 64.945 205.745 65.115 205.935 ;
        RECT 66.325 205.745 66.495 205.935 ;
        RECT 66.840 205.795 66.960 205.905 ;
        RECT 67.245 205.745 67.415 205.935 ;
        RECT 68.625 205.765 68.795 205.955 ;
        RECT 74.145 205.765 74.315 205.955 ;
        RECT 74.605 205.765 74.775 205.955 ;
        RECT 77.365 205.745 77.535 205.955 ;
        RECT 80.585 205.765 80.755 205.955 ;
        RECT 81.100 205.795 81.220 205.905 ;
        RECT 84.725 205.765 84.895 205.955 ;
        RECT 86.565 205.745 86.735 205.935 ;
        RECT 88.405 205.745 88.575 205.935 ;
        RECT 89.380 205.795 89.500 205.905 ;
        RECT 90.245 205.765 90.415 205.955 ;
        RECT 92.085 205.745 92.255 205.935 ;
        RECT 95.765 205.765 95.935 205.955 ;
        RECT 97.605 205.745 97.775 205.935 ;
        RECT 101.285 205.765 101.455 205.955 ;
        RECT 102.260 205.795 102.380 205.905 ;
        RECT 103.125 205.745 103.295 205.935 ;
        RECT 104.045 205.765 104.215 205.955 ;
        RECT 108.645 205.745 108.815 205.935 ;
        RECT 109.565 205.765 109.735 205.955 ;
        RECT 114.165 205.745 114.335 205.935 ;
        RECT 115.085 205.905 115.255 205.955 ;
        RECT 115.085 205.795 115.260 205.905 ;
        RECT 115.085 205.765 115.255 205.795 ;
        RECT 120.605 205.745 120.775 205.955 ;
        RECT 126.125 205.745 126.295 205.955 ;
        RECT 127.505 205.745 127.675 205.955 ;
        RECT 14.665 204.935 16.035 205.745 ;
        RECT 16.965 204.935 20.635 205.745 ;
        RECT 20.645 204.935 26.155 205.745 ;
        RECT 26.165 204.935 31.675 205.745 ;
        RECT 31.685 204.935 37.195 205.745 ;
        RECT 38.125 204.935 40.875 205.745 ;
        RECT 40.885 204.935 46.395 205.745 ;
        RECT 46.405 204.935 51.915 205.745 ;
        RECT 51.925 204.935 57.435 205.745 ;
        RECT 57.445 204.935 62.955 205.745 ;
        RECT 63.425 204.935 65.255 205.745 ;
        RECT 65.275 204.835 66.625 205.745 ;
        RECT 67.115 204.835 68.465 205.745 ;
        RECT 68.485 205.065 77.675 205.745 ;
        RECT 77.685 205.065 86.875 205.745 ;
        RECT 68.485 204.835 69.405 205.065 ;
        RECT 72.235 204.845 73.165 205.065 ;
        RECT 77.685 204.835 78.605 205.065 ;
        RECT 81.435 204.845 82.365 205.065 ;
        RECT 86.885 204.935 88.715 205.745 ;
        RECT 89.645 204.935 92.395 205.745 ;
        RECT 92.405 204.935 97.915 205.745 ;
        RECT 97.925 204.935 103.435 205.745 ;
        RECT 103.445 204.935 108.955 205.745 ;
        RECT 108.965 204.935 114.475 205.745 ;
        RECT 115.405 204.935 120.915 205.745 ;
        RECT 120.925 204.935 126.435 205.745 ;
        RECT 126.445 204.935 127.815 205.745 ;
        RECT 14.665 200.515 16.035 201.325 ;
        RECT 16.045 200.515 18.795 201.325 ;
        RECT 18.805 200.515 24.315 201.325 ;
        RECT 25.245 200.515 27.995 201.325 ;
        RECT 28.005 200.515 33.515 201.325 ;
        RECT 33.525 200.515 39.035 201.325 ;
        RECT 39.045 200.515 44.555 201.325 ;
        RECT 44.565 200.515 50.075 201.325 ;
        RECT 51.005 200.515 54.675 201.325 ;
        RECT 54.685 200.515 60.195 201.325 ;
        RECT 64.715 201.195 65.645 201.415 ;
        RECT 68.365 201.195 70.575 201.425 ;
        RECT 73.110 201.195 74.455 201.425 ;
        RECT 60.205 200.515 70.575 201.195 ;
        RECT 70.785 200.515 72.615 201.195 ;
        RECT 72.625 200.515 74.455 201.195 ;
        RECT 74.465 200.515 75.835 201.325 ;
        RECT 76.305 200.515 78.135 201.195 ;
        RECT 78.145 200.515 79.515 201.295 ;
        RECT 79.525 201.195 80.445 201.425 ;
        RECT 83.275 201.195 84.205 201.415 ;
        RECT 79.525 200.515 88.715 201.195 ;
        RECT 88.725 200.515 90.555 201.325 ;
        RECT 90.565 200.515 96.075 201.325 ;
        RECT 96.085 200.515 101.595 201.325 ;
        RECT 102.525 200.515 104.355 201.325 ;
        RECT 104.365 200.515 109.875 201.325 ;
        RECT 109.885 200.515 115.395 201.325 ;
        RECT 115.405 200.515 120.915 201.325 ;
        RECT 120.925 200.515 126.435 201.325 ;
        RECT 126.445 200.515 127.815 201.325 ;
        RECT 14.805 200.305 14.975 200.515 ;
        RECT 16.645 200.350 16.805 200.460 ;
        RECT 18.485 200.325 18.655 200.515 ;
        RECT 20.325 200.305 20.495 200.495 ;
        RECT 24.005 200.325 24.175 200.515 ;
        RECT 24.980 200.355 25.100 200.465 ;
        RECT 25.845 200.305 26.015 200.495 ;
        RECT 27.685 200.325 27.855 200.515 ;
        RECT 31.365 200.305 31.535 200.495 ;
        RECT 33.205 200.325 33.375 200.515 ;
        RECT 36.885 200.305 37.055 200.495 ;
        RECT 37.860 200.355 37.980 200.465 ;
        RECT 38.725 200.325 38.895 200.515 ;
        RECT 40.565 200.305 40.735 200.495 ;
        RECT 44.245 200.325 44.415 200.515 ;
        RECT 46.085 200.305 46.255 200.495 ;
        RECT 49.765 200.325 49.935 200.515 ;
        RECT 50.740 200.355 50.860 200.465 ;
        RECT 51.605 200.305 51.775 200.495 ;
        RECT 54.365 200.325 54.535 200.515 ;
        RECT 57.125 200.305 57.295 200.495 ;
        RECT 59.885 200.325 60.055 200.515 ;
        RECT 60.345 200.325 60.515 200.515 ;
        RECT 62.645 200.305 62.815 200.495 ;
        RECT 63.620 200.355 63.740 200.465 ;
        RECT 65.405 200.305 65.575 200.495 ;
        RECT 66.785 200.305 66.955 200.495 ;
        RECT 70.465 200.305 70.635 200.495 ;
        RECT 70.925 200.325 71.095 200.515 ;
        RECT 72.765 200.325 72.935 200.515 ;
        RECT 75.065 200.305 75.235 200.495 ;
        RECT 75.525 200.325 75.695 200.515 ;
        RECT 76.445 200.325 76.615 200.515 ;
        RECT 78.285 200.325 78.455 200.515 ;
        RECT 78.745 200.305 78.915 200.495 ;
        RECT 81.045 200.305 81.215 200.495 ;
        RECT 82.430 200.305 82.600 200.495 ;
        RECT 83.805 200.305 83.975 200.495 ;
        RECT 84.265 200.305 84.435 200.495 ;
        RECT 85.700 200.355 85.820 200.465 ;
        RECT 88.405 200.305 88.575 200.515 ;
        RECT 89.380 200.355 89.500 200.465 ;
        RECT 90.245 200.325 90.415 200.515 ;
        RECT 92.085 200.305 92.255 200.495 ;
        RECT 95.765 200.325 95.935 200.515 ;
        RECT 97.605 200.305 97.775 200.495 ;
        RECT 101.285 200.325 101.455 200.515 ;
        RECT 102.260 200.355 102.380 200.465 ;
        RECT 103.125 200.305 103.295 200.495 ;
        RECT 104.045 200.325 104.215 200.515 ;
        RECT 108.645 200.305 108.815 200.495 ;
        RECT 109.565 200.325 109.735 200.515 ;
        RECT 114.165 200.305 114.335 200.495 ;
        RECT 115.085 200.465 115.255 200.515 ;
        RECT 115.085 200.355 115.260 200.465 ;
        RECT 115.085 200.325 115.255 200.355 ;
        RECT 120.605 200.305 120.775 200.515 ;
        RECT 126.125 200.305 126.295 200.515 ;
        RECT 127.505 200.305 127.675 200.515 ;
        RECT 14.665 199.495 16.035 200.305 ;
        RECT 16.965 199.495 20.635 200.305 ;
        RECT 20.645 199.495 26.155 200.305 ;
        RECT 26.165 199.495 31.675 200.305 ;
        RECT 31.685 199.495 37.195 200.305 ;
        RECT 38.125 199.495 40.875 200.305 ;
        RECT 40.885 199.495 46.395 200.305 ;
        RECT 46.405 199.495 51.915 200.305 ;
        RECT 51.925 199.495 57.435 200.305 ;
        RECT 57.445 199.495 62.955 200.305 ;
        RECT 63.885 199.495 65.715 200.305 ;
        RECT 65.725 199.525 67.095 200.305 ;
        RECT 67.105 199.625 70.775 200.305 ;
        RECT 70.795 200.265 71.715 200.305 ;
        RECT 70.785 200.075 71.715 200.265 ;
        RECT 73.805 200.075 75.375 200.305 ;
        RECT 70.785 199.715 75.375 200.075 ;
        RECT 70.795 199.625 75.375 199.715 ;
        RECT 75.480 199.625 78.945 200.305 ;
        RECT 79.065 199.625 81.355 200.305 ;
        RECT 67.105 199.395 68.035 199.625 ;
        RECT 70.795 199.395 73.795 199.625 ;
        RECT 75.480 199.395 76.400 199.625 ;
        RECT 79.065 199.395 79.985 199.625 ;
        RECT 81.365 199.395 82.715 200.305 ;
        RECT 82.755 199.395 84.105 200.305 ;
        RECT 84.135 199.395 85.485 200.305 ;
        RECT 85.965 199.495 88.715 200.305 ;
        RECT 89.645 199.495 92.395 200.305 ;
        RECT 92.405 199.495 97.915 200.305 ;
        RECT 97.925 199.495 103.435 200.305 ;
        RECT 103.445 199.495 108.955 200.305 ;
        RECT 108.965 199.495 114.475 200.305 ;
        RECT 115.405 199.495 120.915 200.305 ;
        RECT 120.925 199.495 126.435 200.305 ;
        RECT 126.445 199.495 127.815 200.305 ;
        RECT 14.665 195.075 16.035 195.885 ;
        RECT 16.045 195.075 18.795 195.885 ;
        RECT 18.805 195.075 24.315 195.885 ;
        RECT 25.245 195.075 27.995 195.885 ;
        RECT 28.005 195.075 33.515 195.885 ;
        RECT 33.525 195.075 39.035 195.885 ;
        RECT 39.045 195.075 44.555 195.885 ;
        RECT 44.565 195.075 50.075 195.885 ;
        RECT 50.545 195.075 52.375 195.885 ;
        RECT 52.395 195.075 53.745 195.985 ;
        RECT 53.765 195.075 55.595 195.885 ;
        RECT 55.615 195.075 56.965 195.985 ;
        RECT 56.985 195.075 58.355 195.885 ;
        RECT 58.365 195.075 63.875 195.885 ;
        RECT 63.885 195.075 69.395 195.885 ;
        RECT 69.405 195.755 70.325 195.985 ;
        RECT 69.405 195.075 71.695 195.755 ;
        RECT 71.705 195.075 74.625 195.985 ;
        RECT 78.275 195.755 79.205 195.985 ;
        RECT 77.370 195.075 79.205 195.755 ;
        RECT 79.525 195.075 85.035 195.885 ;
        RECT 85.045 195.075 90.555 195.885 ;
        RECT 90.565 195.075 96.075 195.885 ;
        RECT 96.085 195.075 101.595 195.885 ;
        RECT 102.065 195.075 107.575 195.885 ;
        RECT 107.595 195.075 108.945 195.985 ;
        RECT 108.965 195.755 109.885 195.985 ;
        RECT 112.715 195.755 113.645 195.975 ;
        RECT 108.965 195.075 118.155 195.755 ;
        RECT 118.165 195.075 120.915 195.885 ;
        RECT 120.925 195.075 126.435 195.885 ;
        RECT 126.445 195.075 127.815 195.885 ;
        RECT 14.805 194.865 14.975 195.075 ;
        RECT 16.645 194.910 16.805 195.020 ;
        RECT 18.485 194.885 18.655 195.075 ;
        RECT 20.325 194.865 20.495 195.055 ;
        RECT 24.005 194.885 24.175 195.075 ;
        RECT 24.980 194.915 25.100 195.025 ;
        RECT 25.845 194.865 26.015 195.055 ;
        RECT 27.685 194.885 27.855 195.075 ;
        RECT 31.365 194.865 31.535 195.055 ;
        RECT 33.205 194.885 33.375 195.075 ;
        RECT 36.885 194.865 37.055 195.055 ;
        RECT 37.860 194.915 37.980 195.025 ;
        RECT 38.725 194.885 38.895 195.075 ;
        RECT 43.325 194.865 43.495 195.055 ;
        RECT 43.785 194.865 43.955 195.055 ;
        RECT 44.245 194.885 44.415 195.075 ;
        RECT 49.765 194.885 49.935 195.075 ;
        RECT 52.065 194.885 52.235 195.075 ;
        RECT 53.445 194.885 53.615 195.075 ;
        RECT 55.285 194.885 55.455 195.075 ;
        RECT 56.665 194.885 56.835 195.075 ;
        RECT 58.045 194.885 58.215 195.075 ;
        RECT 61.725 194.865 61.895 195.055 ;
        RECT 63.565 195.025 63.735 195.075 ;
        RECT 62.645 194.910 62.805 195.020 ;
        RECT 63.565 194.915 63.740 195.025 ;
        RECT 63.565 194.885 63.735 194.915 ;
        RECT 65.405 194.865 65.575 195.055 ;
        RECT 66.785 194.865 66.955 195.055 ;
        RECT 68.165 194.865 68.335 195.055 ;
        RECT 69.085 194.885 69.255 195.075 ;
        RECT 71.385 194.885 71.555 195.075 ;
        RECT 71.850 195.055 72.020 195.075 ;
        RECT 77.370 195.055 77.535 195.075 ;
        RECT 71.845 194.885 72.020 195.055 ;
        RECT 71.845 194.865 72.015 194.885 ;
        RECT 14.665 194.055 16.035 194.865 ;
        RECT 16.965 194.055 20.635 194.865 ;
        RECT 20.645 194.055 26.155 194.865 ;
        RECT 26.165 194.055 31.675 194.865 ;
        RECT 31.685 194.055 37.195 194.865 ;
        RECT 38.125 194.055 43.635 194.865 ;
        RECT 43.645 194.185 52.835 194.865 ;
        RECT 48.155 193.965 49.085 194.185 ;
        RECT 51.915 193.955 52.835 194.185 ;
        RECT 52.845 194.185 62.035 194.865 ;
        RECT 52.845 193.955 53.765 194.185 ;
        RECT 56.595 193.965 57.525 194.185 ;
        RECT 63.885 194.055 65.715 194.865 ;
        RECT 65.735 193.955 67.085 194.865 ;
        RECT 67.105 194.055 68.475 194.865 ;
        RECT 68.485 194.055 72.155 194.865 ;
        RECT 72.305 194.835 72.475 195.055 ;
        RECT 75.525 194.920 75.685 195.030 ;
        RECT 76.905 194.920 77.065 195.030 ;
        RECT 77.365 194.885 77.535 195.055 ;
        RECT 74.430 194.835 75.375 194.865 ;
        RECT 72.305 194.635 75.375 194.835 ;
        RECT 72.165 194.155 75.375 194.635 ;
        RECT 72.165 193.955 73.095 194.155 ;
        RECT 74.430 193.955 75.375 194.155 ;
        RECT 75.385 194.835 76.330 194.865 ;
        RECT 78.285 194.835 78.455 195.055 ;
        RECT 78.800 194.915 78.920 195.025 ;
        RECT 84.265 194.865 84.435 195.055 ;
        RECT 84.725 194.885 84.895 195.075 ;
        RECT 88.130 194.865 88.300 195.055 ;
        RECT 89.380 194.915 89.500 195.025 ;
        RECT 90.245 194.885 90.415 195.075 ;
        RECT 90.705 194.865 90.875 195.055 ;
        RECT 91.220 194.915 91.340 195.025 ;
        RECT 91.625 194.865 91.795 195.055 ;
        RECT 93.060 194.915 93.180 195.025 ;
        RECT 95.765 194.865 95.935 195.075 ;
        RECT 96.225 194.865 96.395 195.055 ;
        RECT 101.285 194.885 101.455 195.075 ;
        RECT 106.345 194.865 106.515 195.055 ;
        RECT 107.265 194.885 107.435 195.075 ;
        RECT 107.725 194.885 107.895 195.075 ;
        RECT 110.025 194.865 110.195 195.055 ;
        RECT 113.890 194.865 114.060 195.055 ;
        RECT 116.005 194.865 116.175 195.055 ;
        RECT 116.925 194.910 117.085 195.020 ;
        RECT 117.845 194.885 118.015 195.075 ;
        RECT 120.605 194.865 120.775 195.075 ;
        RECT 126.125 194.865 126.295 195.075 ;
        RECT 127.505 194.865 127.675 195.075 ;
        RECT 75.385 194.635 78.455 194.835 ;
        RECT 75.385 194.155 78.595 194.635 ;
        RECT 75.385 193.955 76.330 194.155 ;
        RECT 77.665 193.955 78.595 194.155 ;
        RECT 79.065 194.055 84.575 194.865 ;
        RECT 84.815 194.185 88.715 194.865 ;
        RECT 87.785 193.955 88.715 194.185 ;
        RECT 89.655 193.955 91.005 194.865 ;
        RECT 91.485 194.085 92.855 194.865 ;
        RECT 93.325 194.055 96.075 194.865 ;
        RECT 96.095 193.955 97.445 194.865 ;
        RECT 97.465 194.185 106.655 194.865 ;
        RECT 106.760 194.185 110.225 194.865 ;
        RECT 110.575 194.185 114.475 194.865 ;
        RECT 97.465 193.955 98.385 194.185 ;
        RECT 101.215 193.965 102.145 194.185 ;
        RECT 106.760 193.955 107.680 194.185 ;
        RECT 113.545 193.955 114.475 194.185 ;
        RECT 114.955 193.955 116.305 194.865 ;
        RECT 117.245 194.055 120.915 194.865 ;
        RECT 120.925 194.055 126.435 194.865 ;
        RECT 126.445 194.055 127.815 194.865 ;
        RECT 14.665 189.635 16.035 190.445 ;
        RECT 16.045 189.635 18.795 190.445 ;
        RECT 18.805 189.635 24.315 190.445 ;
        RECT 24.785 189.635 26.615 190.445 ;
        RECT 26.625 189.635 32.135 190.445 ;
        RECT 32.145 189.635 37.655 190.445 ;
        RECT 37.665 190.315 38.585 190.545 ;
        RECT 41.415 190.315 42.345 190.535 ;
        RECT 37.665 189.635 46.855 190.315 ;
        RECT 47.325 189.635 50.075 190.445 ;
        RECT 51.465 189.635 52.835 190.415 ;
        RECT 56.045 190.315 56.975 190.545 ;
        RECT 53.075 189.635 56.975 190.315 ;
        RECT 57.905 189.635 59.275 190.415 ;
        RECT 59.285 189.635 62.035 190.445 ;
        RECT 66.555 190.315 67.485 190.535 ;
        RECT 70.315 190.315 71.235 190.545 ;
        RECT 62.045 189.635 71.235 190.315 ;
        RECT 71.245 189.635 74.355 190.545 ;
        RECT 74.465 189.635 75.835 190.445 ;
        RECT 76.305 189.635 78.595 190.545 ;
        RECT 78.605 189.635 80.435 190.445 ;
        RECT 80.445 189.635 85.955 190.445 ;
        RECT 86.335 190.435 87.255 190.545 ;
        RECT 86.335 190.315 88.670 190.435 ;
        RECT 93.335 190.315 94.255 190.535 ;
        RECT 86.335 189.635 95.615 190.315 ;
        RECT 95.625 189.635 97.455 190.445 ;
        RECT 100.665 190.315 101.595 190.545 ;
        RECT 97.695 189.635 101.595 190.315 ;
        RECT 102.525 189.635 103.895 190.415 ;
        RECT 104.365 189.635 106.195 190.445 ;
        RECT 109.405 190.315 110.335 190.545 ;
        RECT 106.435 189.635 110.335 190.315 ;
        RECT 110.345 190.315 111.265 190.545 ;
        RECT 114.095 190.315 115.025 190.535 ;
        RECT 110.345 189.635 119.535 190.315 ;
        RECT 119.545 189.635 120.915 190.445 ;
        RECT 120.925 189.635 126.435 190.445 ;
        RECT 126.445 189.635 127.815 190.445 ;
        RECT 14.805 189.425 14.975 189.635 ;
        RECT 17.565 189.425 17.735 189.615 ;
        RECT 18.485 189.445 18.655 189.635 ;
        RECT 23.085 189.425 23.255 189.615 ;
        RECT 24.005 189.445 24.175 189.635 ;
        RECT 26.305 189.445 26.475 189.635 ;
        RECT 28.605 189.425 28.775 189.615 ;
        RECT 29.985 189.425 30.155 189.615 ;
        RECT 30.500 189.475 30.620 189.585 ;
        RECT 31.825 189.445 31.995 189.635 ;
        RECT 34.125 189.425 34.295 189.615 ;
        RECT 34.585 189.425 34.755 189.615 ;
        RECT 35.965 189.425 36.135 189.615 ;
        RECT 37.345 189.445 37.515 189.635 ;
        RECT 37.805 189.425 37.975 189.615 ;
        RECT 46.545 189.445 46.715 189.635 ;
        RECT 47.060 189.475 47.180 189.585 ;
        RECT 49.765 189.445 49.935 189.635 ;
        RECT 50.870 189.425 51.040 189.615 ;
        RECT 51.145 189.480 51.305 189.590 ;
        RECT 51.605 189.425 51.775 189.615 ;
        RECT 52.525 189.445 52.695 189.635 ;
        RECT 55.340 189.475 55.460 189.585 ;
        RECT 56.390 189.445 56.560 189.635 ;
        RECT 57.125 189.425 57.295 189.615 ;
        RECT 57.585 189.480 57.745 189.590 ;
        RECT 58.045 189.445 58.215 189.635 ;
        RECT 61.725 189.445 61.895 189.635 ;
        RECT 62.185 189.445 62.355 189.635 ;
        RECT 62.645 189.425 62.815 189.615 ;
        RECT 64.485 189.425 64.655 189.615 ;
        RECT 68.165 189.425 68.335 189.615 ;
        RECT 68.625 189.425 68.795 189.615 ;
        RECT 73.225 189.425 73.395 189.615 ;
        RECT 74.145 189.445 74.315 189.635 ;
        RECT 75.525 189.445 75.695 189.635 ;
        RECT 78.280 189.445 78.450 189.635 ;
        RECT 78.745 189.425 78.915 189.615 ;
        RECT 80.125 189.445 80.295 189.635 ;
        RECT 85.645 189.445 85.815 189.635 ;
        RECT 88.405 189.425 88.575 189.615 ;
        RECT 90.245 189.425 90.415 189.615 ;
        RECT 91.625 189.425 91.795 189.615 ;
        RECT 94.385 189.425 94.555 189.615 ;
        RECT 94.845 189.425 95.015 189.615 ;
        RECT 95.305 189.445 95.475 189.635 ;
        RECT 97.145 189.445 97.315 189.635 ;
        RECT 101.010 189.445 101.180 189.635 ;
        RECT 102.260 189.475 102.380 189.585 ;
        RECT 102.665 189.445 102.835 189.635 ;
        RECT 104.100 189.475 104.220 189.585 ;
        RECT 105.885 189.445 106.055 189.635 ;
        RECT 107.265 189.425 107.435 189.615 ;
        RECT 109.750 189.445 109.920 189.635 ;
        RECT 112.785 189.425 112.955 189.615 ;
        RECT 113.245 189.425 113.415 189.615 ;
        RECT 115.545 189.470 115.705 189.580 ;
        RECT 116.005 189.425 116.175 189.615 ;
        RECT 119.225 189.445 119.395 189.635 ;
        RECT 120.605 189.425 120.775 189.635 ;
        RECT 126.125 189.425 126.295 189.635 ;
        RECT 127.505 189.425 127.675 189.635 ;
        RECT 14.665 188.615 16.035 189.425 ;
        RECT 16.045 188.615 17.875 189.425 ;
        RECT 17.885 188.615 23.395 189.425 ;
        RECT 23.405 188.615 28.915 189.425 ;
        RECT 28.935 188.515 30.285 189.425 ;
        RECT 30.765 188.615 34.435 189.425 ;
        RECT 34.455 188.515 35.805 189.425 ;
        RECT 35.825 188.645 37.195 189.425 ;
        RECT 37.665 188.745 46.945 189.425 ;
        RECT 47.555 188.745 51.455 189.425 ;
        RECT 51.575 188.745 55.040 189.425 ;
        RECT 39.025 188.525 39.945 188.745 ;
        RECT 44.610 188.625 46.945 188.745 ;
        RECT 46.025 188.515 46.945 188.625 ;
        RECT 50.525 188.515 51.455 188.745 ;
        RECT 54.120 188.515 55.040 188.745 ;
        RECT 55.605 188.615 57.435 189.425 ;
        RECT 57.445 188.615 62.955 189.425 ;
        RECT 63.425 188.615 64.795 189.425 ;
        RECT 64.805 188.615 68.475 189.425 ;
        RECT 68.595 188.745 72.060 189.425 ;
        RECT 71.140 188.515 72.060 188.745 ;
        RECT 72.165 188.615 73.535 189.425 ;
        RECT 73.545 188.615 79.055 189.425 ;
        RECT 79.435 188.745 88.715 189.425 ;
        RECT 79.435 188.625 81.770 188.745 ;
        RECT 79.435 188.515 80.355 188.625 ;
        RECT 86.435 188.525 87.355 188.745 ;
        RECT 89.195 188.515 90.545 189.425 ;
        RECT 90.565 188.645 91.935 189.425 ;
        RECT 91.945 188.615 94.695 189.425 ;
        RECT 94.815 188.745 98.280 189.425 ;
        RECT 97.360 188.515 98.280 188.745 ;
        RECT 98.385 188.745 107.575 189.425 ;
        RECT 98.385 188.515 99.305 188.745 ;
        RECT 102.135 188.525 103.065 188.745 ;
        RECT 107.585 188.615 113.095 189.425 ;
        RECT 113.105 188.645 114.475 189.425 ;
        RECT 115.865 188.645 117.235 189.425 ;
        RECT 117.245 188.615 120.915 189.425 ;
        RECT 120.925 188.615 126.435 189.425 ;
        RECT 126.445 188.615 127.815 189.425 ;
        RECT 14.665 184.195 16.035 185.005 ;
        RECT 16.045 184.195 18.795 185.005 ;
        RECT 18.805 184.195 24.315 185.005 ;
        RECT 30.215 184.875 31.145 185.095 ;
        RECT 33.975 184.875 34.895 185.105 ;
        RECT 25.705 184.195 34.895 184.875 ;
        RECT 34.905 184.195 37.655 185.005 ;
        RECT 37.675 184.195 39.025 185.105 ;
        RECT 39.045 184.875 39.975 185.105 ;
        RECT 44.105 184.875 45.035 185.105 ;
        RECT 39.045 184.195 42.945 184.875 ;
        RECT 44.105 184.195 48.005 184.875 ;
        RECT 48.715 184.195 50.065 185.105 ;
        RECT 50.545 184.875 51.465 185.105 ;
        RECT 54.295 184.875 55.225 185.095 ;
        RECT 50.545 184.195 59.735 184.875 ;
        RECT 59.745 184.195 61.115 185.005 ;
        RECT 61.125 184.195 64.795 185.005 ;
        RECT 64.805 184.195 70.315 185.005 ;
        RECT 70.325 184.195 75.835 185.005 ;
        RECT 76.765 184.195 79.515 185.005 ;
        RECT 82.180 184.875 83.100 185.105 ;
        RECT 79.635 184.195 83.100 184.875 ;
        RECT 83.205 184.195 85.035 185.005 ;
        RECT 88.245 184.875 89.175 185.105 ;
        RECT 85.275 184.195 89.175 184.875 ;
        RECT 89.195 184.195 90.545 185.105 ;
        RECT 90.565 184.195 92.395 185.005 ;
        RECT 95.060 184.875 95.980 185.105 ;
        RECT 99.285 184.875 100.215 185.105 ;
        RECT 92.515 184.195 95.980 184.875 ;
        RECT 96.315 184.195 100.215 184.875 ;
        RECT 100.225 184.195 101.595 184.975 ;
        RECT 102.075 184.195 103.425 185.105 ;
        RECT 103.905 184.195 107.575 185.005 ;
        RECT 110.240 184.875 111.160 185.105 ;
        RECT 107.695 184.195 111.160 184.875 ;
        RECT 111.725 184.195 115.395 185.005 ;
        RECT 115.405 184.195 120.915 185.005 ;
        RECT 120.925 184.195 126.435 185.005 ;
        RECT 126.445 184.195 127.815 185.005 ;
        RECT 14.805 183.985 14.975 184.195 ;
        RECT 16.240 184.035 16.360 184.145 ;
        RECT 18.485 184.005 18.655 184.195 ;
        RECT 21.705 183.985 21.875 184.175 ;
        RECT 22.165 183.985 22.335 184.175 ;
        RECT 24.005 184.005 24.175 184.195 ;
        RECT 25.385 184.040 25.545 184.150 ;
        RECT 25.845 184.005 26.015 184.195 ;
        RECT 26.765 183.985 26.935 184.175 ;
        RECT 27.225 183.985 27.395 184.175 ;
        RECT 31.180 183.985 31.350 184.175 ;
        RECT 35.100 184.035 35.220 184.145 ;
        RECT 36.885 183.985 37.055 184.175 ;
        RECT 37.345 184.005 37.515 184.195 ;
        RECT 37.805 183.985 37.975 184.195 ;
        RECT 39.460 184.005 39.630 184.195 ;
        RECT 41.540 184.035 41.660 184.145 ;
        RECT 41.945 183.985 42.115 184.175 ;
        RECT 43.325 183.985 43.495 184.175 ;
        RECT 43.785 184.040 43.945 184.150 ;
        RECT 44.520 184.005 44.690 184.195 ;
        RECT 47.005 183.985 47.175 184.175 ;
        RECT 48.440 184.035 48.560 184.145 ;
        RECT 49.765 184.005 49.935 184.195 ;
        RECT 50.960 183.985 51.130 184.175 ;
        RECT 54.880 184.035 55.000 184.145 ;
        RECT 55.285 183.985 55.455 184.175 ;
        RECT 56.665 183.985 56.835 184.175 ;
        RECT 59.425 184.005 59.595 184.195 ;
        RECT 60.345 183.985 60.515 184.175 ;
        RECT 60.805 184.005 60.975 184.195 ;
        RECT 62.645 183.985 62.815 184.175 ;
        RECT 63.620 184.035 63.740 184.145 ;
        RECT 64.485 184.005 64.655 184.195 ;
        RECT 66.325 183.985 66.495 184.175 ;
        RECT 70.005 184.005 70.175 184.195 ;
        RECT 71.845 183.985 72.015 184.175 ;
        RECT 72.305 184.005 72.475 184.175 ;
        RECT 75.525 184.145 75.695 184.195 ;
        RECT 79.205 184.175 79.375 184.195 ;
        RECT 75.525 184.035 75.700 184.145 ;
        RECT 76.500 184.035 76.620 184.145 ;
        RECT 75.525 184.005 75.695 184.035 ;
        RECT 79.200 184.005 79.375 184.175 ;
        RECT 79.665 184.005 79.835 184.195 ;
        RECT 84.725 184.005 84.895 184.195 ;
        RECT 72.405 183.985 72.475 184.005 ;
        RECT 79.200 183.985 79.370 184.005 ;
        RECT 88.405 183.985 88.575 184.175 ;
        RECT 88.590 184.005 88.760 184.195 ;
        RECT 89.785 184.030 89.945 184.140 ;
        RECT 90.245 184.005 90.415 184.195 ;
        RECT 91.165 183.985 91.335 184.175 ;
        RECT 92.085 184.005 92.255 184.195 ;
        RECT 92.545 184.005 92.715 184.195 ;
        RECT 99.630 184.005 99.800 184.195 ;
        RECT 100.365 184.005 100.535 184.195 ;
        RECT 101.285 183.985 101.455 184.175 ;
        RECT 102.205 184.030 102.365 184.140 ;
        RECT 102.940 183.985 103.110 184.175 ;
        RECT 103.125 184.005 103.295 184.195 ;
        RECT 103.640 184.035 103.760 184.145 ;
        RECT 107.265 184.005 107.435 184.195 ;
        RECT 107.725 184.005 107.895 184.195 ;
        RECT 110.025 183.985 110.195 184.175 ;
        RECT 111.460 184.035 111.580 184.145 ;
        RECT 113.890 183.985 114.060 184.175 ;
        RECT 115.085 184.145 115.255 184.195 ;
        RECT 115.085 184.035 115.260 184.145 ;
        RECT 115.085 184.005 115.255 184.035 ;
        RECT 120.605 184.005 120.775 184.195 ;
        RECT 124.285 183.985 124.455 184.175 ;
        RECT 126.125 183.985 126.295 184.195 ;
        RECT 127.505 183.985 127.675 184.195 ;
        RECT 14.665 183.175 16.035 183.985 ;
        RECT 16.505 183.175 22.015 183.985 ;
        RECT 22.025 183.205 23.395 183.985 ;
        RECT 23.500 183.305 26.965 183.985 ;
        RECT 27.195 183.305 30.660 183.985 ;
        RECT 23.500 183.075 24.420 183.305 ;
        RECT 29.740 183.075 30.660 183.305 ;
        RECT 30.765 183.305 34.665 183.985 ;
        RECT 30.765 183.075 31.695 183.305 ;
        RECT 35.365 183.175 37.195 183.985 ;
        RECT 37.775 183.305 41.240 183.985 ;
        RECT 40.320 183.075 41.240 183.305 ;
        RECT 41.805 183.205 43.175 183.985 ;
        RECT 43.295 183.305 46.760 183.985 ;
        RECT 46.975 183.305 50.440 183.985 ;
        RECT 45.840 183.075 46.760 183.305 ;
        RECT 49.520 183.075 50.440 183.305 ;
        RECT 50.545 183.305 54.445 183.985 ;
        RECT 50.545 183.075 51.475 183.305 ;
        RECT 55.155 183.075 56.505 183.985 ;
        RECT 56.635 183.305 60.100 183.985 ;
        RECT 59.180 183.075 60.100 183.305 ;
        RECT 60.205 183.205 61.575 183.985 ;
        RECT 61.585 183.205 62.955 183.985 ;
        RECT 63.885 183.175 66.635 183.985 ;
        RECT 66.645 183.175 72.155 183.985 ;
        RECT 72.405 183.755 74.675 183.985 ;
        RECT 72.405 183.075 75.160 183.755 ;
        RECT 76.040 183.075 79.515 183.985 ;
        RECT 79.525 183.305 88.715 183.985 ;
        RECT 79.525 183.075 80.445 183.305 ;
        RECT 83.275 183.085 84.205 183.305 ;
        RECT 90.105 183.205 91.475 183.985 ;
        RECT 92.405 183.305 101.595 183.985 ;
        RECT 102.525 183.305 106.425 183.985 ;
        RECT 106.760 183.305 110.225 183.985 ;
        RECT 110.575 183.305 114.475 183.985 ;
        RECT 92.405 183.075 93.325 183.305 ;
        RECT 96.155 183.085 97.085 183.305 ;
        RECT 102.525 183.075 103.455 183.305 ;
        RECT 106.760 183.075 107.680 183.305 ;
        RECT 113.545 183.075 114.475 183.305 ;
        RECT 115.405 183.305 124.595 183.985 ;
        RECT 115.405 183.075 116.325 183.305 ;
        RECT 119.155 183.085 120.085 183.305 ;
        RECT 124.605 183.175 126.435 183.985 ;
        RECT 126.445 183.175 127.815 183.985 ;
        RECT 14.665 178.755 16.035 179.565 ;
        RECT 16.045 178.755 18.795 179.565 ;
        RECT 18.805 178.755 24.315 179.565 ;
        RECT 29.295 179.435 30.225 179.655 ;
        RECT 33.055 179.435 33.975 179.665 ;
        RECT 37.100 179.435 38.020 179.665 ;
        RECT 24.785 178.755 33.975 179.435 ;
        RECT 34.555 178.755 38.020 179.435 ;
        RECT 38.585 178.755 39.955 179.535 ;
        RECT 40.885 178.755 46.395 179.565 ;
        RECT 49.060 179.435 49.980 179.665 ;
        RECT 54.120 179.435 55.040 179.665 ;
        RECT 46.515 178.755 49.980 179.435 ;
        RECT 51.575 178.755 55.040 179.435 ;
        RECT 55.145 179.435 56.065 179.665 ;
        RECT 58.895 179.435 59.825 179.655 ;
        RECT 55.145 178.755 64.335 179.435 ;
        RECT 64.815 178.755 66.165 179.665 ;
        RECT 66.185 179.435 67.530 179.665 ;
        RECT 66.185 178.755 68.015 179.435 ;
        RECT 68.265 178.985 71.020 179.665 ;
        RECT 71.255 179.435 74.255 179.665 ;
        RECT 71.255 179.345 75.835 179.435 ;
        RECT 71.245 178.985 75.835 179.345 ;
        RECT 68.265 178.755 70.535 178.985 ;
        RECT 71.245 178.795 72.175 178.985 ;
        RECT 71.255 178.755 72.175 178.795 ;
        RECT 74.265 178.755 75.835 178.985 ;
        RECT 76.545 178.985 79.300 179.665 ;
        RECT 82.725 179.435 83.655 179.665 ;
        RECT 76.545 178.755 78.815 178.985 ;
        RECT 79.755 178.755 83.655 179.435 ;
        RECT 83.665 178.755 92.770 179.435 ;
        RECT 92.865 178.755 94.235 179.565 ;
        RECT 96.900 179.435 97.820 179.665 ;
        RECT 100.580 179.435 101.500 179.665 ;
        RECT 94.355 178.755 97.820 179.435 ;
        RECT 98.035 178.755 101.500 179.435 ;
        RECT 102.065 178.755 103.435 179.535 ;
        RECT 103.905 178.755 107.380 179.665 ;
        RECT 110.785 179.435 111.715 179.665 ;
        RECT 107.815 178.755 111.715 179.435 ;
        RECT 111.725 179.435 112.645 179.665 ;
        RECT 115.475 179.435 116.405 179.655 ;
        RECT 111.725 178.755 120.915 179.435 ;
        RECT 120.925 178.755 122.295 179.535 ;
        RECT 122.305 178.755 123.675 179.535 ;
        RECT 123.685 178.755 126.435 179.565 ;
        RECT 126.445 178.755 127.815 179.565 ;
        RECT 14.805 178.545 14.975 178.755 ;
        RECT 18.485 178.565 18.655 178.755 ;
        RECT 19.405 178.545 19.575 178.735 ;
        RECT 24.005 178.565 24.175 178.755 ;
        RECT 24.925 178.545 25.095 178.755 ;
        RECT 26.305 178.545 26.475 178.735 ;
        RECT 27.685 178.545 27.855 178.735 ;
        RECT 34.180 178.595 34.300 178.705 ;
        RECT 34.585 178.565 34.755 178.755 ;
        RECT 36.885 178.545 37.055 178.735 ;
        RECT 38.080 178.545 38.250 178.735 ;
        RECT 38.320 178.595 38.440 178.705 ;
        RECT 39.645 178.565 39.815 178.755 ;
        RECT 40.565 178.600 40.725 178.710 ;
        RECT 43.325 178.545 43.495 178.735 ;
        RECT 46.085 178.565 46.255 178.755 ;
        RECT 46.545 178.565 46.715 178.755 ;
        RECT 51.605 178.735 51.775 178.755 ;
        RECT 47.000 178.545 47.170 178.735 ;
        RECT 47.520 178.595 47.640 178.705 ;
        RECT 47.930 178.545 48.100 178.735 ;
        RECT 51.145 178.600 51.305 178.710 ;
        RECT 51.605 178.565 51.780 178.735 ;
        RECT 55.340 178.595 55.460 178.705 ;
        RECT 51.610 178.545 51.780 178.565 ;
        RECT 59.150 178.545 59.320 178.735 ;
        RECT 59.940 178.595 60.060 178.705 ;
        RECT 62.645 178.545 62.815 178.735 ;
        RECT 63.620 178.595 63.740 178.705 ;
        RECT 64.025 178.565 64.195 178.755 ;
        RECT 64.540 178.595 64.660 178.705 ;
        RECT 65.405 178.545 65.575 178.735 ;
        RECT 65.865 178.565 66.035 178.755 ;
        RECT 67.245 178.545 67.415 178.735 ;
        RECT 67.705 178.705 67.875 178.755 ;
        RECT 68.265 178.735 68.335 178.755 ;
        RECT 67.705 178.595 67.880 178.705 ;
        RECT 67.705 178.565 67.875 178.595 ;
        RECT 68.165 178.545 68.335 178.735 ;
        RECT 70.925 178.565 71.095 178.735 ;
        RECT 75.525 178.565 75.695 178.755 ;
        RECT 76.545 178.735 76.615 178.755 ;
        RECT 76.445 178.565 76.615 178.735 ;
        RECT 71.025 178.545 71.095 178.565 ;
        RECT 77.360 178.545 77.530 178.735 ;
        RECT 83.070 178.565 83.240 178.755 ;
        RECT 83.805 178.565 83.975 178.755 ;
        RECT 88.400 178.545 88.570 178.735 ;
        RECT 89.785 178.590 89.945 178.700 ;
        RECT 93.925 178.565 94.095 178.755 ;
        RECT 94.385 178.565 94.555 178.755 ;
        RECT 95.305 178.545 95.475 178.735 ;
        RECT 96.685 178.545 96.855 178.735 ;
        RECT 98.065 178.565 98.235 178.755 ;
        RECT 98.525 178.545 98.695 178.735 ;
        RECT 98.990 178.545 99.160 178.735 ;
        RECT 103.125 178.565 103.295 178.755 ;
        RECT 103.640 178.595 103.760 178.705 ;
        RECT 104.050 178.565 104.220 178.755 ;
        RECT 104.965 178.545 105.135 178.735 ;
        RECT 105.430 178.545 105.600 178.735 ;
        RECT 111.130 178.565 111.300 178.755 ;
        RECT 112.325 178.545 112.495 178.735 ;
        RECT 112.840 178.595 112.960 178.705 ;
        RECT 113.245 178.545 113.415 178.735 ;
        RECT 116.465 178.545 116.635 178.735 ;
        RECT 116.925 178.545 117.095 178.735 ;
        RECT 120.605 178.545 120.775 178.755 ;
        RECT 121.985 178.565 122.155 178.755 ;
        RECT 122.445 178.565 122.615 178.755 ;
        RECT 126.125 178.545 126.295 178.755 ;
        RECT 127.505 178.545 127.675 178.755 ;
        RECT 14.665 177.735 16.035 178.545 ;
        RECT 16.045 177.735 19.715 178.545 ;
        RECT 19.725 177.735 25.235 178.545 ;
        RECT 25.255 177.635 26.605 178.545 ;
        RECT 26.625 177.765 27.995 178.545 ;
        RECT 28.005 177.865 37.195 178.545 ;
        RECT 37.665 177.865 41.565 178.545 ;
        RECT 28.005 177.635 28.925 177.865 ;
        RECT 31.755 177.645 32.685 177.865 ;
        RECT 37.665 177.635 38.595 177.865 ;
        RECT 41.805 177.735 43.635 178.545 ;
        RECT 43.840 177.635 47.315 178.545 ;
        RECT 47.785 177.635 51.260 178.545 ;
        RECT 51.465 177.635 54.940 178.545 ;
        RECT 55.835 177.865 59.735 178.545 ;
        RECT 60.215 177.865 62.955 178.545 ;
        RECT 63.885 177.865 65.715 178.545 ;
        RECT 65.725 177.865 67.555 178.545 ;
        RECT 58.805 177.635 59.735 177.865 ;
        RECT 63.885 177.635 65.230 177.865 ;
        RECT 65.725 177.635 67.070 177.865 ;
        RECT 68.025 177.635 70.745 178.545 ;
        RECT 71.025 178.315 73.295 178.545 ;
        RECT 71.025 177.635 73.780 178.315 ;
        RECT 74.200 177.635 77.675 178.545 ;
        RECT 77.705 177.635 88.715 178.545 ;
        RECT 90.105 177.735 95.615 178.545 ;
        RECT 95.635 177.635 96.985 178.545 ;
        RECT 97.005 177.735 98.835 178.545 ;
        RECT 98.845 177.635 102.320 178.545 ;
        RECT 102.525 177.735 105.275 178.545 ;
        RECT 105.285 177.635 108.760 178.545 ;
        RECT 109.060 177.865 112.525 178.545 ;
        RECT 109.060 177.635 109.980 177.865 ;
        RECT 113.115 177.635 114.465 178.545 ;
        RECT 114.945 177.735 116.775 178.545 ;
        RECT 116.795 177.635 118.145 178.545 ;
        RECT 118.165 177.735 120.915 178.545 ;
        RECT 120.925 177.735 126.435 178.545 ;
        RECT 126.445 177.735 127.815 178.545 ;
        RECT 14.665 173.315 16.035 174.125 ;
        RECT 16.045 173.315 18.795 174.125 ;
        RECT 18.805 173.315 24.315 174.125 ;
        RECT 25.715 173.315 27.065 174.225 ;
        RECT 29.740 173.995 30.660 174.225 ;
        RECT 27.195 173.315 30.660 173.995 ;
        RECT 31.225 173.995 32.155 174.225 ;
        RECT 31.225 173.315 35.125 173.995 ;
        RECT 35.560 173.315 39.035 174.225 ;
        RECT 39.045 173.315 42.520 174.225 ;
        RECT 42.920 173.315 46.395 174.225 ;
        RECT 46.405 173.315 49.880 174.225 ;
        RECT 50.545 173.315 51.915 174.125 ;
        RECT 54.580 173.995 55.500 174.225 ;
        RECT 59.725 173.995 60.655 174.225 ;
        RECT 52.035 173.315 55.500 173.995 ;
        RECT 56.755 173.315 60.655 173.995 ;
        RECT 60.665 173.315 62.495 174.125 ;
        RECT 62.505 173.315 63.875 174.095 ;
        RECT 64.345 173.315 68.015 174.125 ;
        RECT 68.025 173.315 70.635 174.225 ;
        RECT 71.245 173.995 72.590 174.225 ;
        RECT 73.570 173.995 74.915 174.225 ;
        RECT 71.245 173.315 73.075 173.995 ;
        RECT 73.085 173.315 74.915 173.995 ;
        RECT 77.420 173.315 80.895 174.225 ;
        RECT 80.905 173.315 84.380 174.225 ;
        RECT 84.680 173.995 85.600 174.225 ;
        RECT 84.680 173.315 88.145 173.995 ;
        RECT 88.265 173.315 91.005 173.995 ;
        RECT 91.025 173.315 92.395 174.125 ;
        RECT 92.405 173.315 96.075 174.125 ;
        RECT 96.085 173.315 101.595 174.125 ;
        RECT 102.065 173.315 111.170 173.995 ;
        RECT 111.265 173.315 114.740 174.225 ;
        RECT 115.140 173.315 118.615 174.225 ;
        RECT 118.635 173.315 119.985 174.225 ;
        RECT 120.925 173.315 126.435 174.125 ;
        RECT 126.445 173.315 127.815 174.125 ;
        RECT 14.805 173.105 14.975 173.315 ;
        RECT 16.645 173.150 16.805 173.260 ;
        RECT 18.485 173.125 18.655 173.315 ;
        RECT 22.165 173.105 22.335 173.295 ;
        RECT 24.005 173.125 24.175 173.315 ;
        RECT 25.385 173.160 25.545 173.270 ;
        RECT 26.765 173.125 26.935 173.315 ;
        RECT 27.225 173.125 27.395 173.315 ;
        RECT 27.685 173.105 27.855 173.295 ;
        RECT 30.960 173.155 31.080 173.265 ;
        RECT 31.640 173.125 31.810 173.315 ;
        RECT 33.205 173.105 33.375 173.295 ;
        RECT 36.880 173.105 37.050 173.295 ;
        RECT 37.860 173.155 37.980 173.265 ;
        RECT 38.270 173.105 38.440 173.295 ;
        RECT 38.720 173.125 38.890 173.315 ;
        RECT 39.190 173.125 39.360 173.315 ;
        RECT 44.245 173.105 44.415 173.295 ;
        RECT 46.080 173.125 46.250 173.315 ;
        RECT 46.550 173.125 46.720 173.315 ;
        RECT 51.605 173.125 51.775 173.315 ;
        RECT 52.065 173.125 52.235 173.315 ;
        RECT 53.445 173.105 53.615 173.295 ;
        RECT 56.205 173.160 56.365 173.270 ;
        RECT 60.070 173.125 60.240 173.315 ;
        RECT 62.185 173.125 62.355 173.315 ;
        RECT 62.645 173.105 62.815 173.295 ;
        RECT 63.565 173.125 63.735 173.315 ;
        RECT 64.080 173.155 64.200 173.265 ;
        RECT 64.485 173.105 64.655 173.295 ;
        RECT 65.405 173.150 65.565 173.260 ;
        RECT 67.705 173.125 67.875 173.315 ;
        RECT 68.170 173.125 68.340 173.315 ;
        RECT 70.925 173.265 71.095 173.295 ;
        RECT 70.925 173.155 71.100 173.265 ;
        RECT 70.925 173.105 71.095 173.155 ;
        RECT 72.765 173.125 72.935 173.315 ;
        RECT 73.225 173.125 73.395 173.315 ;
        RECT 75.525 173.160 75.685 173.270 ;
        RECT 76.445 173.105 76.615 173.295 ;
        RECT 76.905 173.160 77.065 173.270 ;
        RECT 80.580 173.125 80.750 173.315 ;
        RECT 81.050 173.125 81.220 173.315 ;
        RECT 81.965 173.105 82.135 173.295 ;
        RECT 82.430 173.105 82.600 173.295 ;
        RECT 85.185 173.105 85.355 173.295 ;
        RECT 87.945 173.125 88.115 173.315 ;
        RECT 88.405 173.125 88.575 173.315 ;
        RECT 89.380 173.155 89.500 173.265 ;
        RECT 89.785 173.105 89.955 173.295 ;
        RECT 92.085 173.125 92.255 173.315 ;
        RECT 95.765 173.125 95.935 173.315 ;
        RECT 99.905 173.105 100.075 173.295 ;
        RECT 100.825 173.150 100.985 173.260 ;
        RECT 101.285 173.125 101.455 173.315 ;
        RECT 102.205 173.125 102.375 173.315 ;
        RECT 104.505 173.105 104.675 173.295 ;
        RECT 107.725 173.125 107.895 173.295 ;
        RECT 108.190 173.105 108.360 173.295 ;
        RECT 111.410 173.125 111.580 173.315 ;
        RECT 112.785 173.105 112.955 173.295 ;
        RECT 113.245 173.105 113.415 173.295 ;
        RECT 115.545 173.150 115.705 173.260 ;
        RECT 118.300 173.125 118.470 173.315 ;
        RECT 119.685 173.125 119.855 173.315 ;
        RECT 120.605 173.160 120.765 173.270 ;
        RECT 124.745 173.105 124.915 173.295 ;
        RECT 126.125 173.105 126.295 173.315 ;
        RECT 127.505 173.105 127.675 173.315 ;
        RECT 14.665 172.295 16.035 173.105 ;
        RECT 16.965 172.295 22.475 173.105 ;
        RECT 22.485 172.295 27.995 173.105 ;
        RECT 28.005 172.295 33.515 173.105 ;
        RECT 33.720 172.195 37.195 173.105 ;
        RECT 38.125 172.195 41.600 173.105 ;
        RECT 41.805 172.295 44.555 173.105 ;
        RECT 44.650 172.425 53.755 173.105 ;
        RECT 53.765 172.425 62.955 173.105 ;
        RECT 53.765 172.195 54.685 172.425 ;
        RECT 57.515 172.205 58.445 172.425 ;
        RECT 63.435 172.195 64.785 173.105 ;
        RECT 65.725 172.295 71.235 173.105 ;
        RECT 71.245 172.295 76.755 173.105 ;
        RECT 76.765 172.295 82.275 173.105 ;
        RECT 82.285 172.195 84.895 173.105 ;
        RECT 85.155 172.425 88.620 173.105 ;
        RECT 87.700 172.195 88.620 172.425 ;
        RECT 89.655 172.195 91.005 173.105 ;
        RECT 91.025 172.425 100.215 173.105 ;
        RECT 91.025 172.195 91.945 172.425 ;
        RECT 94.775 172.205 95.705 172.425 ;
        RECT 101.145 172.295 104.815 173.105 ;
        RECT 105.205 172.425 107.630 173.105 ;
        RECT 108.045 172.195 111.520 173.105 ;
        RECT 111.725 172.295 113.095 173.105 ;
        RECT 113.115 172.195 114.465 173.105 ;
        RECT 115.865 172.425 125.055 173.105 ;
        RECT 115.865 172.195 116.785 172.425 ;
        RECT 119.615 172.205 120.545 172.425 ;
        RECT 125.065 172.295 126.435 173.105 ;
        RECT 126.445 172.295 127.815 173.105 ;
        RECT 14.665 167.875 16.035 168.685 ;
        RECT 16.045 167.875 18.795 168.685 ;
        RECT 18.805 167.875 24.315 168.685 ;
        RECT 25.245 167.875 27.075 168.685 ;
        RECT 27.095 167.875 28.445 168.785 ;
        RECT 28.465 167.875 30.295 168.685 ;
        RECT 30.315 167.875 31.665 168.785 ;
        RECT 34.340 168.555 35.260 168.785 ;
        RECT 31.795 167.875 35.260 168.555 ;
        RECT 36.025 167.875 38.115 168.685 ;
        RECT 38.125 167.875 39.955 168.685 ;
        RECT 39.965 167.875 45.475 168.685 ;
        RECT 45.485 167.875 48.960 168.785 ;
        RECT 50.545 167.875 52.375 168.685 ;
        RECT 52.765 167.875 55.190 168.555 ;
        RECT 55.605 167.875 57.435 168.685 ;
        RECT 57.445 167.875 62.955 168.685 ;
        RECT 62.965 167.875 68.475 168.685 ;
        RECT 68.970 168.555 70.315 168.785 ;
        RECT 68.485 167.875 70.315 168.555 ;
        RECT 70.325 168.555 71.670 168.785 ;
        RECT 79.505 168.555 80.435 168.785 ;
        RECT 70.325 167.875 72.155 168.555 ;
        RECT 72.625 167.875 75.365 168.555 ;
        RECT 76.535 167.875 80.435 168.555 ;
        RECT 80.815 168.675 81.735 168.785 ;
        RECT 80.815 168.555 83.150 168.675 ;
        RECT 87.815 168.555 88.735 168.775 ;
        RECT 94.225 168.555 95.155 168.785 ;
        RECT 80.815 167.875 90.095 168.555 ;
        RECT 91.255 167.875 95.155 168.555 ;
        RECT 96.085 167.875 97.455 168.655 ;
        RECT 97.925 167.875 101.595 168.685 ;
        RECT 102.525 168.555 103.445 168.785 ;
        RECT 106.275 168.555 107.205 168.775 ;
        RECT 112.645 168.555 113.575 168.785 ;
        RECT 116.880 168.555 117.800 168.785 ;
        RECT 102.525 167.875 111.715 168.555 ;
        RECT 112.645 167.875 116.545 168.555 ;
        RECT 116.880 167.875 120.345 168.555 ;
        RECT 120.475 167.875 121.825 168.785 ;
        RECT 121.845 167.875 123.675 168.555 ;
        RECT 123.685 167.875 125.055 168.655 ;
        RECT 125.065 167.875 126.435 168.685 ;
        RECT 126.445 167.875 127.815 168.685 ;
        RECT 14.805 167.665 14.975 167.875 ;
        RECT 16.240 167.715 16.360 167.825 ;
        RECT 18.025 167.665 18.195 167.855 ;
        RECT 18.485 167.685 18.655 167.875 ;
        RECT 24.005 167.685 24.175 167.875 ;
        RECT 24.980 167.715 25.100 167.825 ;
        RECT 26.765 167.685 26.935 167.875 ;
        RECT 27.225 167.665 27.395 167.855 ;
        RECT 28.145 167.685 28.315 167.875 ;
        RECT 29.985 167.685 30.155 167.875 ;
        RECT 31.365 167.685 31.535 167.875 ;
        RECT 31.825 167.685 31.995 167.875 ;
        RECT 36.425 167.665 36.595 167.855 ;
        RECT 36.940 167.715 37.060 167.825 ;
        RECT 37.805 167.685 37.975 167.875 ;
        RECT 38.725 167.665 38.895 167.855 ;
        RECT 39.645 167.685 39.815 167.875 ;
        RECT 40.105 167.665 40.275 167.855 ;
        RECT 40.620 167.715 40.740 167.825 ;
        RECT 41.025 167.665 41.195 167.855 ;
        RECT 42.405 167.665 42.575 167.855 ;
        RECT 43.785 167.665 43.955 167.855 ;
        RECT 45.165 167.685 45.335 167.875 ;
        RECT 45.630 167.685 45.800 167.875 ;
        RECT 49.765 167.720 49.925 167.830 ;
        RECT 52.065 167.685 52.235 167.875 ;
        RECT 55.285 167.685 55.455 167.855 ;
        RECT 56.205 167.665 56.375 167.855 ;
        RECT 57.125 167.685 57.295 167.875 ;
        RECT 58.505 167.665 58.675 167.855 ;
        RECT 59.425 167.710 59.585 167.820 ;
        RECT 62.180 167.665 62.350 167.855 ;
        RECT 62.645 167.825 62.815 167.875 ;
        RECT 62.645 167.715 62.820 167.825 ;
        RECT 62.645 167.685 62.815 167.715 ;
        RECT 64.025 167.710 64.185 167.820 ;
        RECT 66.780 167.665 66.950 167.855 ;
        RECT 68.165 167.685 68.335 167.875 ;
        RECT 68.625 167.685 68.795 167.875 ;
        RECT 69.545 167.665 69.715 167.855 ;
        RECT 70.925 167.665 71.095 167.855 ;
        RECT 71.385 167.665 71.555 167.855 ;
        RECT 71.845 167.685 72.015 167.875 ;
        RECT 72.360 167.715 72.480 167.825 ;
        RECT 72.765 167.685 72.935 167.875 ;
        RECT 75.065 167.665 75.235 167.855 ;
        RECT 75.580 167.715 75.700 167.825 ;
        RECT 79.850 167.685 80.020 167.875 ;
        RECT 84.725 167.665 84.895 167.855 ;
        RECT 86.105 167.665 86.275 167.855 ;
        RECT 87.485 167.665 87.655 167.855 ;
        RECT 88.405 167.710 88.565 167.820 ;
        RECT 89.380 167.715 89.500 167.825 ;
        RECT 89.785 167.685 89.955 167.875 ;
        RECT 90.705 167.720 90.865 167.830 ;
        RECT 91.165 167.665 91.335 167.855 ;
        RECT 94.570 167.685 94.740 167.875 ;
        RECT 95.765 167.720 95.925 167.830 ;
        RECT 96.225 167.685 96.395 167.875 ;
        RECT 96.685 167.665 96.855 167.855 ;
        RECT 97.660 167.715 97.780 167.825 ;
        RECT 101.285 167.685 101.455 167.875 ;
        RECT 102.260 167.715 102.380 167.825 ;
        RECT 106.345 167.665 106.515 167.855 ;
        RECT 106.860 167.715 106.980 167.825 ;
        RECT 107.265 167.665 107.435 167.855 ;
        RECT 111.405 167.685 111.575 167.875 ;
        RECT 112.325 167.720 112.485 167.830 ;
        RECT 113.060 167.685 113.230 167.875 ;
        RECT 114.165 167.665 114.335 167.855 ;
        RECT 115.545 167.710 115.705 167.820 ;
        RECT 120.145 167.685 120.315 167.875 ;
        RECT 120.605 167.685 120.775 167.875 ;
        RECT 123.365 167.685 123.535 167.875 ;
        RECT 124.745 167.665 124.915 167.875 ;
        RECT 126.125 167.665 126.295 167.875 ;
        RECT 127.505 167.665 127.675 167.875 ;
        RECT 14.665 166.855 16.035 167.665 ;
        RECT 16.505 166.855 18.335 167.665 ;
        RECT 18.345 166.985 27.535 167.665 ;
        RECT 27.630 166.985 36.735 167.665 ;
        RECT 18.345 166.755 19.265 166.985 ;
        RECT 22.095 166.765 23.025 166.985 ;
        RECT 37.665 166.885 39.035 167.665 ;
        RECT 39.055 166.755 40.405 167.665 ;
        RECT 40.885 166.885 42.255 167.665 ;
        RECT 42.275 166.755 43.625 167.665 ;
        RECT 43.755 166.985 47.220 167.665 ;
        RECT 46.300 166.755 47.220 166.985 ;
        RECT 47.325 166.985 56.515 167.665 ;
        RECT 47.325 166.755 48.245 166.985 ;
        RECT 51.075 166.765 52.005 166.985 ;
        RECT 57.455 166.755 58.805 167.665 ;
        RECT 59.885 166.755 62.495 167.665 ;
        RECT 64.485 166.755 67.095 167.665 ;
        RECT 67.115 166.985 69.855 167.665 ;
        RECT 69.865 166.855 71.235 167.665 ;
        RECT 71.245 166.755 73.965 167.665 ;
        RECT 74.005 166.855 75.375 167.665 ;
        RECT 75.755 166.985 85.035 167.665 ;
        RECT 75.755 166.865 78.090 166.985 ;
        RECT 75.755 166.755 76.675 166.865 ;
        RECT 82.755 166.765 83.675 166.985 ;
        RECT 85.055 166.755 86.405 167.665 ;
        RECT 86.435 166.755 87.785 167.665 ;
        RECT 89.645 166.855 91.475 167.665 ;
        RECT 91.485 166.855 96.995 167.665 ;
        RECT 97.375 166.985 106.655 167.665 ;
        RECT 107.235 166.985 110.700 167.665 ;
        RECT 97.375 166.865 99.710 166.985 ;
        RECT 97.375 166.755 98.295 166.865 ;
        RECT 104.375 166.765 105.295 166.985 ;
        RECT 109.780 166.755 110.700 166.985 ;
        RECT 110.900 166.985 114.365 167.665 ;
        RECT 115.865 166.985 125.055 167.665 ;
        RECT 110.900 166.755 111.820 166.985 ;
        RECT 115.865 166.755 116.785 166.985 ;
        RECT 119.615 166.765 120.545 166.985 ;
        RECT 125.065 166.855 126.435 167.665 ;
        RECT 126.445 166.855 127.815 167.665 ;
        RECT 14.665 162.435 16.035 163.245 ;
        RECT 16.045 162.435 18.795 163.245 ;
        RECT 18.805 162.435 24.315 163.245 ;
        RECT 25.705 162.435 27.075 163.215 ;
        RECT 27.085 163.115 28.005 163.345 ;
        RECT 30.835 163.115 31.765 163.335 ;
        RECT 36.285 163.115 37.205 163.345 ;
        RECT 40.035 163.115 40.965 163.335 ;
        RECT 45.485 163.115 46.415 163.345 ;
        RECT 53.745 163.115 54.675 163.345 ;
        RECT 27.085 162.435 36.275 163.115 ;
        RECT 36.285 162.435 45.475 163.115 ;
        RECT 45.485 162.435 49.385 163.115 ;
        RECT 50.775 162.435 54.675 163.115 ;
        RECT 54.685 163.115 55.605 163.345 ;
        RECT 58.435 163.115 59.365 163.335 ;
        RECT 54.685 162.435 63.875 163.115 ;
        RECT 64.345 162.435 67.095 163.245 ;
        RECT 67.115 162.435 69.855 163.115 ;
        RECT 70.325 162.435 75.835 163.245 ;
        RECT 76.305 162.435 78.135 163.245 ;
        RECT 81.345 163.115 82.275 163.345 ;
        RECT 78.375 162.435 82.275 163.115 ;
        RECT 82.285 162.435 83.655 163.215 ;
        RECT 83.665 162.435 85.495 163.245 ;
        RECT 85.505 162.435 86.875 163.215 ;
        RECT 87.805 162.435 93.315 163.245 ;
        RECT 96.525 163.115 97.455 163.345 ;
        RECT 100.665 163.115 101.595 163.345 ;
        RECT 93.555 162.435 97.455 163.115 ;
        RECT 97.695 162.435 101.595 163.115 ;
        RECT 102.160 163.115 103.080 163.345 ;
        RECT 106.665 163.115 107.595 163.345 ;
        RECT 102.160 162.435 105.625 163.115 ;
        RECT 106.665 162.435 110.565 163.115 ;
        RECT 110.815 162.435 112.165 163.345 ;
        RECT 113.105 163.115 114.025 163.345 ;
        RECT 116.855 163.115 117.785 163.335 ;
        RECT 113.105 162.435 122.295 163.115 ;
        RECT 122.305 162.435 123.675 163.215 ;
        RECT 123.685 162.435 126.435 163.245 ;
        RECT 126.445 162.435 127.815 163.245 ;
        RECT 14.805 162.225 14.975 162.435 ;
        RECT 17.565 162.225 17.735 162.415 ;
        RECT 18.485 162.245 18.655 162.435 ;
        RECT 24.005 162.245 24.175 162.435 ;
        RECT 25.385 162.280 25.545 162.390 ;
        RECT 26.765 162.245 26.935 162.435 ;
        RECT 27.225 162.225 27.395 162.415 ;
        RECT 27.960 162.225 28.130 162.415 ;
        RECT 32.745 162.225 32.915 162.415 ;
        RECT 35.965 162.245 36.135 162.435 ;
        RECT 36.610 162.225 36.780 162.415 ;
        RECT 37.860 162.275 37.980 162.385 ;
        RECT 41.485 162.225 41.655 162.415 ;
        RECT 45.165 162.225 45.335 162.435 ;
        RECT 45.900 162.245 46.070 162.435 ;
        RECT 46.545 162.225 46.715 162.415 ;
        RECT 47.005 162.225 47.175 162.415 ;
        RECT 49.820 162.275 49.940 162.385 ;
        RECT 54.090 162.225 54.260 162.435 ;
        RECT 54.825 162.225 54.995 162.415 ;
        RECT 58.560 162.275 58.680 162.385 ;
        RECT 58.965 162.225 59.135 162.415 ;
        RECT 62.645 162.225 62.815 162.415 ;
        RECT 63.565 162.245 63.735 162.435 ;
        RECT 64.080 162.275 64.200 162.385 ;
        RECT 64.485 162.225 64.655 162.415 ;
        RECT 66.325 162.225 66.495 162.415 ;
        RECT 66.785 162.245 66.955 162.435 ;
        RECT 68.165 162.225 68.335 162.415 ;
        RECT 68.625 162.225 68.795 162.415 ;
        RECT 69.545 162.245 69.715 162.435 ;
        RECT 70.060 162.275 70.180 162.385 ;
        RECT 70.465 162.225 70.635 162.415 ;
        RECT 74.605 162.225 74.775 162.415 ;
        RECT 75.525 162.245 75.695 162.435 ;
        RECT 77.825 162.245 77.995 162.435 ;
        RECT 80.125 162.225 80.295 162.415 ;
        RECT 81.505 162.225 81.675 162.415 ;
        RECT 81.690 162.245 81.860 162.435 ;
        RECT 82.425 162.245 82.595 162.435 ;
        RECT 85.185 162.245 85.355 162.435 ;
        RECT 85.370 162.225 85.540 162.415 ;
        RECT 85.645 162.245 85.815 162.435 ;
        RECT 86.160 162.275 86.280 162.385 ;
        RECT 86.565 162.225 86.735 162.415 ;
        RECT 87.485 162.280 87.645 162.390 ;
        RECT 88.405 162.270 88.565 162.380 ;
        RECT 93.005 162.245 93.175 162.435 ;
        RECT 96.870 162.245 97.040 162.435 ;
        RECT 98.525 162.225 98.695 162.415 ;
        RECT 99.445 162.270 99.605 162.380 ;
        RECT 99.905 162.225 100.075 162.415 ;
        RECT 101.010 162.245 101.180 162.435 ;
        RECT 102.205 162.225 102.375 162.415 ;
        RECT 105.425 162.245 105.595 162.435 ;
        RECT 105.885 162.225 106.055 162.415 ;
        RECT 106.345 162.385 106.505 162.390 ;
        RECT 106.345 162.280 106.520 162.385 ;
        RECT 106.400 162.275 106.520 162.280 ;
        RECT 106.805 162.225 106.975 162.415 ;
        RECT 107.080 162.245 107.250 162.435 ;
        RECT 111.865 162.245 112.035 162.435 ;
        RECT 112.785 162.280 112.945 162.390 ;
        RECT 113.890 162.225 114.060 162.415 ;
        RECT 118.490 162.225 118.660 162.415 ;
        RECT 119.225 162.225 119.395 162.415 ;
        RECT 121.985 162.245 122.155 162.435 ;
        RECT 122.905 162.225 123.075 162.415 ;
        RECT 123.365 162.245 123.535 162.435 ;
        RECT 124.340 162.275 124.460 162.385 ;
        RECT 126.125 162.225 126.295 162.435 ;
        RECT 127.505 162.225 127.675 162.435 ;
        RECT 14.665 161.415 16.035 162.225 ;
        RECT 16.045 161.415 17.875 162.225 ;
        RECT 18.255 161.545 27.535 162.225 ;
        RECT 27.545 161.545 31.445 162.225 ;
        RECT 18.255 161.425 20.590 161.545 ;
        RECT 18.255 161.315 19.175 161.425 ;
        RECT 25.255 161.325 26.175 161.545 ;
        RECT 27.545 161.315 28.475 161.545 ;
        RECT 31.685 161.415 33.055 162.225 ;
        RECT 33.295 161.545 37.195 162.225 ;
        RECT 36.265 161.315 37.195 161.545 ;
        RECT 38.125 161.415 41.795 162.225 ;
        RECT 41.900 161.545 45.365 162.225 ;
        RECT 41.900 161.315 42.820 161.545 ;
        RECT 45.485 161.415 46.855 162.225 ;
        RECT 46.975 161.545 50.440 162.225 ;
        RECT 50.775 161.545 54.675 162.225 ;
        RECT 54.795 161.545 58.260 162.225 ;
        RECT 49.520 161.315 50.440 161.545 ;
        RECT 53.745 161.315 54.675 161.545 ;
        RECT 57.340 161.315 58.260 161.545 ;
        RECT 58.825 161.445 60.195 162.225 ;
        RECT 60.205 161.415 62.955 162.225 ;
        RECT 63.425 161.415 64.795 162.225 ;
        RECT 64.805 161.545 66.635 162.225 ;
        RECT 66.645 161.545 68.475 162.225 ;
        RECT 68.485 161.545 70.315 162.225 ;
        RECT 70.325 161.545 72.155 162.225 ;
        RECT 64.805 161.315 66.150 161.545 ;
        RECT 66.645 161.315 67.990 161.545 ;
        RECT 68.970 161.315 70.315 161.545 ;
        RECT 70.810 161.315 72.155 161.545 ;
        RECT 72.165 161.415 74.915 162.225 ;
        RECT 74.925 161.415 80.435 162.225 ;
        RECT 80.455 161.315 81.805 162.225 ;
        RECT 82.055 161.545 85.955 162.225 ;
        RECT 85.025 161.315 85.955 161.545 ;
        RECT 86.425 161.445 87.795 162.225 ;
        RECT 89.555 161.545 98.835 162.225 ;
        RECT 89.555 161.425 91.890 161.545 ;
        RECT 89.555 161.315 90.475 161.425 ;
        RECT 96.555 161.325 97.475 161.545 ;
        RECT 99.765 161.445 101.135 162.225 ;
        RECT 101.155 161.315 102.505 162.225 ;
        RECT 102.620 161.545 106.085 162.225 ;
        RECT 106.775 161.545 110.240 162.225 ;
        RECT 110.575 161.545 114.475 162.225 ;
        RECT 115.175 161.545 119.075 162.225 ;
        RECT 119.195 161.545 122.660 162.225 ;
        RECT 102.620 161.315 103.540 161.545 ;
        RECT 109.320 161.315 110.240 161.545 ;
        RECT 113.545 161.315 114.475 161.545 ;
        RECT 118.145 161.315 119.075 161.545 ;
        RECT 121.740 161.315 122.660 161.545 ;
        RECT 122.765 161.445 124.135 162.225 ;
        RECT 124.605 161.415 126.435 162.225 ;
        RECT 126.445 161.415 127.815 162.225 ;
        RECT 14.665 156.995 16.035 157.805 ;
        RECT 16.045 156.995 17.415 157.805 ;
        RECT 17.435 156.995 18.785 157.905 ;
        RECT 18.815 156.995 20.165 157.905 ;
        RECT 23.385 157.675 24.315 157.905 ;
        RECT 20.415 156.995 24.315 157.675 ;
        RECT 24.785 156.995 26.155 157.775 ;
        RECT 26.625 156.995 32.135 157.805 ;
        RECT 32.240 157.675 33.160 157.905 ;
        RECT 32.240 156.995 35.705 157.675 ;
        RECT 35.825 156.995 37.195 157.805 ;
        RECT 37.205 156.995 42.715 157.805 ;
        RECT 42.920 156.995 46.395 157.905 ;
        RECT 46.405 156.995 49.880 157.905 ;
        RECT 50.545 156.995 54.020 157.905 ;
        RECT 54.685 156.995 56.055 157.775 ;
        RECT 56.065 156.995 61.575 157.805 ;
        RECT 61.725 156.995 64.335 157.905 ;
        RECT 64.805 156.995 68.475 157.805 ;
        RECT 68.970 157.675 70.315 157.905 ;
        RECT 70.810 157.675 72.155 157.905 ;
        RECT 68.485 156.995 70.315 157.675 ;
        RECT 70.325 156.995 72.155 157.675 ;
        RECT 72.360 156.995 75.835 157.905 ;
        RECT 76.765 156.995 80.240 157.905 ;
        RECT 80.815 157.795 81.735 157.905 ;
        RECT 80.815 157.675 83.150 157.795 ;
        RECT 87.815 157.675 88.735 157.895 ;
        RECT 80.815 156.995 90.095 157.675 ;
        RECT 90.105 156.995 92.855 157.805 ;
        RECT 92.875 156.995 94.225 157.905 ;
        RECT 94.245 156.995 96.075 157.805 ;
        RECT 96.085 156.995 97.455 157.775 ;
        RECT 97.925 156.995 101.595 157.805 ;
        RECT 102.525 156.995 105.275 157.805 ;
        RECT 105.285 156.995 106.655 157.775 ;
        RECT 106.665 156.995 108.035 157.805 ;
        RECT 108.045 156.995 113.555 157.805 ;
        RECT 113.565 156.995 119.075 157.805 ;
        RECT 119.225 156.995 121.835 157.905 ;
        RECT 122.765 156.995 126.435 157.805 ;
        RECT 126.445 156.995 127.815 157.805 ;
        RECT 14.805 156.785 14.975 156.995 ;
        RECT 16.240 156.835 16.360 156.945 ;
        RECT 17.105 156.805 17.275 156.995 ;
        RECT 18.485 156.805 18.655 156.995 ;
        RECT 18.945 156.805 19.115 156.995 ;
        RECT 23.730 156.805 23.900 156.995 ;
        RECT 24.925 156.805 25.095 156.995 ;
        RECT 25.845 156.785 26.015 156.975 ;
        RECT 26.360 156.835 26.480 156.945 ;
        RECT 27.225 156.785 27.395 156.975 ;
        RECT 28.145 156.830 28.305 156.940 ;
        RECT 31.825 156.785 31.995 156.995 ;
        RECT 32.285 156.785 32.455 156.975 ;
        RECT 35.505 156.805 35.675 156.995 ;
        RECT 36.885 156.785 37.055 156.995 ;
        RECT 37.860 156.835 37.980 156.945 ;
        RECT 39.645 156.785 39.815 156.975 ;
        RECT 40.110 156.785 40.280 156.975 ;
        RECT 42.405 156.805 42.575 156.995 ;
        RECT 43.790 156.785 43.960 156.975 ;
        RECT 46.080 156.805 46.250 156.995 ;
        RECT 46.550 156.805 46.720 156.995 ;
        RECT 50.690 156.975 50.860 156.995 ;
        RECT 50.680 156.805 50.860 156.975 ;
        RECT 51.200 156.835 51.320 156.945 ;
        RECT 50.680 156.785 50.850 156.805 ;
        RECT 52.985 156.785 53.155 156.975 ;
        RECT 54.420 156.835 54.540 156.945 ;
        RECT 55.745 156.805 55.915 156.995 ;
        RECT 61.265 156.805 61.435 156.995 ;
        RECT 62.645 156.785 62.815 156.975 ;
        RECT 63.565 156.785 63.735 156.975 ;
        RECT 64.020 156.805 64.190 156.995 ;
        RECT 64.540 156.835 64.660 156.945 ;
        RECT 66.325 156.785 66.495 156.975 ;
        RECT 68.165 156.805 68.335 156.995 ;
        RECT 68.625 156.805 68.795 156.995 ;
        RECT 70.465 156.805 70.635 156.995 ;
        RECT 75.520 156.975 75.690 156.995 ;
        RECT 75.520 156.805 75.695 156.975 ;
        RECT 76.500 156.835 76.620 156.945 ;
        RECT 76.910 156.805 77.080 156.995 ;
        RECT 75.525 156.785 75.695 156.805 ;
        RECT 79.200 156.785 79.370 156.975 ;
        RECT 80.125 156.830 80.285 156.940 ;
        RECT 80.590 156.785 80.760 156.975 ;
        RECT 84.725 156.830 84.885 156.940 ;
        RECT 88.405 156.785 88.575 156.975 ;
        RECT 89.785 156.805 89.955 156.995 ;
        RECT 91.625 156.785 91.795 156.975 ;
        RECT 92.545 156.805 92.715 156.995 ;
        RECT 93.925 156.805 94.095 156.995 ;
        RECT 95.765 156.805 95.935 156.995 ;
        RECT 97.145 156.785 97.315 156.995 ;
        RECT 97.610 156.785 97.780 156.975 ;
        RECT 101.285 156.945 101.455 156.995 ;
        RECT 101.285 156.835 101.460 156.945 ;
        RECT 102.260 156.835 102.380 156.945 ;
        RECT 101.285 156.805 101.455 156.835 ;
        RECT 103.125 156.785 103.295 156.975 ;
        RECT 104.965 156.805 105.135 156.995 ;
        RECT 105.425 156.805 105.595 156.995 ;
        RECT 106.800 156.785 106.970 156.975 ;
        RECT 107.725 156.805 107.895 156.995 ;
        RECT 110.480 156.785 110.650 156.975 ;
        RECT 110.950 156.785 111.120 156.975 ;
        RECT 113.245 156.805 113.415 156.995 ;
        RECT 116.005 156.785 116.175 156.975 ;
        RECT 116.470 156.785 116.640 156.975 ;
        RECT 118.765 156.805 118.935 156.995 ;
        RECT 120.605 156.785 120.775 156.975 ;
        RECT 121.520 156.805 121.690 156.995 ;
        RECT 122.445 156.840 122.605 156.950 ;
        RECT 126.125 156.785 126.295 156.995 ;
        RECT 127.505 156.785 127.675 156.995 ;
        RECT 14.665 155.975 16.035 156.785 ;
        RECT 16.875 156.105 26.155 156.785 ;
        RECT 16.875 155.985 19.210 156.105 ;
        RECT 16.875 155.875 17.795 155.985 ;
        RECT 23.875 155.885 24.795 156.105 ;
        RECT 26.165 156.005 27.535 156.785 ;
        RECT 28.465 155.975 32.135 156.785 ;
        RECT 32.255 156.105 35.720 156.785 ;
        RECT 34.800 155.875 35.720 156.105 ;
        RECT 35.825 155.975 37.195 156.785 ;
        RECT 38.125 155.975 39.955 156.785 ;
        RECT 39.965 155.875 43.440 156.785 ;
        RECT 43.645 155.875 47.120 156.785 ;
        RECT 47.520 155.875 50.995 156.785 ;
        RECT 51.465 155.975 53.295 156.785 ;
        RECT 53.675 156.105 62.955 156.785 ;
        RECT 53.675 155.985 56.010 156.105 ;
        RECT 53.675 155.875 54.595 155.985 ;
        RECT 60.675 155.885 61.595 156.105 ;
        RECT 63.435 155.875 64.785 156.785 ;
        RECT 64.805 155.975 66.635 156.785 ;
        RECT 66.730 156.105 75.835 156.785 ;
        RECT 76.040 155.875 79.515 156.785 ;
        RECT 80.445 155.875 83.920 156.785 ;
        RECT 85.045 155.975 88.715 156.785 ;
        RECT 89.185 155.975 91.935 156.785 ;
        RECT 91.945 155.975 97.455 156.785 ;
        RECT 97.465 155.875 100.940 156.785 ;
        RECT 101.605 155.975 103.435 156.785 ;
        RECT 103.640 155.875 107.115 156.785 ;
        RECT 107.320 155.875 110.795 156.785 ;
        RECT 110.805 155.875 114.280 156.785 ;
        RECT 114.945 155.975 116.315 156.785 ;
        RECT 116.325 155.875 118.935 156.785 ;
        RECT 119.085 155.975 120.915 156.785 ;
        RECT 120.925 155.975 126.435 156.785 ;
        RECT 126.445 155.975 127.815 156.785 ;
        RECT 14.665 151.555 16.035 152.365 ;
        RECT 16.505 151.555 20.175 152.365 ;
        RECT 23.385 152.235 24.315 152.465 ;
        RECT 20.415 151.555 24.315 152.235 ;
        RECT 25.245 151.555 30.755 152.365 ;
        RECT 30.775 151.555 32.125 152.465 ;
        RECT 32.145 151.555 33.515 152.335 ;
        RECT 33.525 152.235 34.455 152.465 ;
        RECT 33.525 151.555 37.425 152.235 ;
        RECT 37.665 151.555 41.140 152.465 ;
        RECT 41.805 151.555 44.555 152.365 ;
        RECT 44.565 151.555 50.075 152.365 ;
        RECT 51.465 151.555 56.975 152.365 ;
        RECT 56.995 151.555 58.345 152.465 ;
        RECT 58.735 152.355 59.655 152.465 ;
        RECT 58.735 152.235 61.070 152.355 ;
        RECT 65.735 152.235 66.655 152.455 ;
        RECT 58.735 151.555 68.015 152.235 ;
        RECT 68.485 151.555 71.235 152.365 ;
        RECT 71.730 152.235 73.075 152.465 ;
        RECT 71.245 151.555 73.075 152.235 ;
        RECT 73.085 151.555 75.805 152.465 ;
        RECT 76.765 151.555 79.515 152.365 ;
        RECT 79.525 151.555 85.035 152.365 ;
        RECT 85.045 151.555 90.555 152.365 ;
        RECT 90.575 151.555 91.925 152.465 ;
        RECT 92.405 151.555 96.075 152.365 ;
        RECT 96.085 151.555 101.595 152.365 ;
        RECT 102.525 151.555 105.275 152.365 ;
        RECT 105.285 151.555 108.760 152.465 ;
        RECT 108.965 151.555 112.440 152.465 ;
        RECT 113.105 151.555 118.615 152.365 ;
        RECT 118.635 151.555 119.985 152.465 ;
        RECT 120.465 151.555 121.835 152.335 ;
        RECT 122.765 151.555 126.435 152.365 ;
        RECT 126.445 151.555 127.815 152.365 ;
        RECT 14.805 151.345 14.975 151.555 ;
        RECT 16.240 151.395 16.360 151.505 ;
        RECT 19.865 151.365 20.035 151.555 ;
        RECT 23.730 151.365 23.900 151.555 ;
        RECT 24.980 151.395 25.100 151.505 ;
        RECT 25.385 151.345 25.555 151.535 ;
        RECT 27.225 151.345 27.395 151.535 ;
        RECT 30.445 151.365 30.615 151.555 ;
        RECT 30.905 151.365 31.075 151.555 ;
        RECT 32.285 151.365 32.455 151.555 ;
        RECT 33.940 151.365 34.110 151.555 ;
        RECT 36.885 151.345 37.055 151.535 ;
        RECT 37.810 151.365 37.980 151.555 ;
        RECT 44.245 151.535 44.415 151.555 ;
        RECT 40.565 151.345 40.735 151.535 ;
        RECT 41.540 151.395 41.660 151.505 ;
        RECT 44.240 151.365 44.415 151.535 ;
        RECT 44.240 151.345 44.410 151.365 ;
        RECT 45.625 151.345 45.795 151.535 ;
        RECT 14.665 150.535 16.035 151.345 ;
        RECT 16.415 150.665 25.695 151.345 ;
        RECT 16.415 150.545 18.750 150.665 ;
        RECT 16.415 150.435 17.335 150.545 ;
        RECT 23.415 150.445 24.335 150.665 ;
        RECT 25.705 150.535 27.535 151.345 ;
        RECT 27.915 150.665 37.195 151.345 ;
        RECT 27.915 150.545 30.250 150.665 ;
        RECT 27.915 150.435 28.835 150.545 ;
        RECT 34.915 150.445 35.835 150.665 ;
        RECT 38.125 150.535 40.875 151.345 ;
        RECT 41.080 150.435 44.555 151.345 ;
        RECT 44.565 150.535 45.935 151.345 ;
        RECT 46.090 151.315 46.260 151.535 ;
        RECT 47.750 151.315 48.695 151.345 ;
        RECT 48.850 151.315 49.020 151.535 ;
        RECT 49.765 151.365 49.935 151.555 ;
        RECT 51.145 151.400 51.305 151.510 ;
        RECT 51.610 151.345 51.780 151.535 ;
        RECT 55.340 151.395 55.460 151.505 ;
        RECT 56.665 151.365 56.835 151.555 ;
        RECT 57.125 151.345 57.295 151.555 ;
        RECT 60.990 151.345 61.160 151.535 ;
        RECT 62.645 151.345 62.815 151.535 ;
        RECT 63.620 151.395 63.740 151.505 ;
        RECT 64.025 151.345 64.195 151.535 ;
        RECT 65.460 151.395 65.580 151.505 ;
        RECT 67.245 151.345 67.415 151.535 ;
        RECT 67.705 151.345 67.875 151.555 ;
        RECT 68.220 151.395 68.340 151.505 ;
        RECT 70.925 151.345 71.095 151.555 ;
        RECT 71.385 151.365 71.555 151.555 ;
        RECT 73.225 151.365 73.395 151.555 ;
        RECT 73.685 151.345 73.855 151.535 ;
        RECT 74.605 151.390 74.765 151.500 ;
        RECT 75.065 151.345 75.235 151.535 ;
        RECT 76.500 151.395 76.620 151.505 ;
        RECT 50.510 151.315 51.455 151.345 ;
        RECT 45.945 150.635 48.695 151.315 ;
        RECT 48.705 150.635 51.455 151.315 ;
        RECT 47.750 150.435 48.695 150.635 ;
        RECT 50.510 150.435 51.455 150.635 ;
        RECT 51.465 150.435 54.940 151.345 ;
        RECT 55.605 150.535 57.435 151.345 ;
        RECT 57.675 150.665 61.575 151.345 ;
        RECT 60.645 150.435 61.575 150.665 ;
        RECT 61.585 150.565 62.955 151.345 ;
        RECT 63.885 150.565 65.255 151.345 ;
        RECT 65.725 150.535 67.555 151.345 ;
        RECT 67.565 150.665 69.395 151.345 ;
        RECT 68.050 150.435 69.395 150.665 ;
        RECT 69.405 150.665 71.235 151.345 ;
        RECT 71.255 150.665 73.995 151.345 ;
        RECT 74.925 150.665 77.665 151.345 ;
        RECT 77.830 151.315 78.000 151.535 ;
        RECT 79.205 151.365 79.375 151.555 ;
        RECT 80.640 151.395 80.760 151.505 ;
        RECT 84.265 151.345 84.435 151.535 ;
        RECT 84.725 151.365 84.895 151.555 ;
        RECT 88.130 151.345 88.300 151.535 ;
        RECT 89.325 151.345 89.495 151.535 ;
        RECT 90.245 151.365 90.415 151.555 ;
        RECT 90.705 151.365 90.875 151.555 ;
        RECT 92.140 151.395 92.260 151.505 ;
        RECT 95.765 151.365 95.935 151.555 ;
        RECT 101.285 151.365 101.455 151.555 ;
        RECT 102.260 151.395 102.380 151.505 ;
        RECT 104.045 151.345 104.215 151.535 ;
        RECT 104.965 151.365 105.135 151.555 ;
        RECT 105.430 151.365 105.600 151.555 ;
        RECT 79.490 151.315 80.435 151.345 ;
        RECT 69.405 150.435 70.750 150.665 ;
        RECT 77.685 150.635 80.435 151.315 ;
        RECT 79.490 150.435 80.435 150.635 ;
        RECT 80.905 150.535 84.575 151.345 ;
        RECT 84.815 150.665 88.715 151.345 ;
        RECT 89.185 150.665 98.465 151.345 ;
        RECT 87.785 150.435 88.715 150.665 ;
        RECT 90.545 150.445 91.465 150.665 ;
        RECT 96.130 150.545 98.465 150.665 ;
        RECT 97.545 150.435 98.465 150.545 ;
        RECT 98.845 150.535 104.355 151.345 ;
        RECT 104.365 151.315 105.310 151.345 ;
        RECT 106.800 151.315 106.970 151.535 ;
        RECT 107.270 151.345 107.440 151.535 ;
        RECT 109.110 151.365 109.280 151.555 ;
        RECT 110.945 151.345 111.115 151.535 ;
        RECT 112.840 151.395 112.960 151.505 ;
        RECT 115.545 151.390 115.705 151.500 ;
        RECT 118.305 151.365 118.475 151.555 ;
        RECT 119.685 151.365 119.855 151.555 ;
        RECT 120.200 151.395 120.320 151.505 ;
        RECT 120.605 151.365 120.775 151.555 ;
        RECT 122.445 151.400 122.605 151.510 ;
        RECT 124.745 151.345 124.915 151.535 ;
        RECT 126.125 151.345 126.295 151.555 ;
        RECT 127.505 151.345 127.675 151.555 ;
        RECT 104.365 150.635 107.115 151.315 ;
        RECT 104.365 150.435 105.310 150.635 ;
        RECT 107.125 150.435 110.600 151.345 ;
        RECT 110.915 150.665 114.380 151.345 ;
        RECT 113.460 150.435 114.380 150.665 ;
        RECT 115.865 150.665 125.055 151.345 ;
        RECT 115.865 150.435 116.785 150.665 ;
        RECT 119.615 150.445 120.545 150.665 ;
        RECT 125.065 150.535 126.435 151.345 ;
        RECT 126.445 150.535 127.815 151.345 ;
        RECT 14.665 146.115 16.035 146.925 ;
        RECT 16.505 146.115 20.175 146.925 ;
        RECT 23.385 146.795 24.315 147.025 ;
        RECT 20.415 146.115 24.315 146.795 ;
        RECT 25.255 146.115 26.605 147.025 ;
        RECT 26.625 146.115 27.995 146.895 ;
        RECT 28.005 146.115 29.375 146.895 ;
        RECT 29.385 146.795 30.315 147.025 ;
        RECT 29.385 146.115 33.285 146.795 ;
        RECT 33.985 146.115 35.815 146.925 ;
        RECT 36.020 146.115 39.495 147.025 ;
        RECT 39.505 146.115 42.980 147.025 ;
        RECT 43.185 146.115 44.555 146.925 ;
        RECT 44.565 146.115 50.075 146.925 ;
        RECT 51.465 146.795 52.395 147.025 ;
        RECT 51.465 146.115 55.365 146.795 ;
        RECT 55.605 146.115 59.080 147.025 ;
        RECT 62.945 146.795 63.875 147.025 ;
        RECT 59.975 146.115 63.875 146.795 ;
        RECT 63.885 146.115 65.255 146.925 ;
        RECT 65.265 146.115 70.775 146.925 ;
        RECT 70.785 146.795 72.130 147.025 ;
        RECT 73.110 146.795 74.455 147.025 ;
        RECT 70.785 146.115 72.615 146.795 ;
        RECT 72.625 146.115 74.455 146.795 ;
        RECT 74.465 146.115 75.835 146.925 ;
        RECT 76.500 146.115 79.975 147.025 ;
        RECT 79.985 146.115 83.460 147.025 ;
        RECT 83.675 146.115 85.025 147.025 ;
        RECT 85.415 146.915 86.335 147.025 ;
        RECT 85.415 146.795 87.750 146.915 ;
        RECT 92.415 146.795 93.335 147.015 ;
        RECT 85.415 146.115 94.695 146.795 ;
        RECT 95.635 146.115 96.985 147.025 ;
        RECT 100.205 146.795 101.135 147.025 ;
        RECT 97.235 146.115 101.135 146.795 ;
        RECT 102.065 146.115 103.435 146.895 ;
        RECT 103.905 146.825 104.850 147.025 ;
        RECT 103.905 146.145 106.655 146.825 ;
        RECT 103.905 146.115 104.850 146.145 ;
        RECT 14.805 145.905 14.975 146.115 ;
        RECT 16.240 145.955 16.360 146.065 ;
        RECT 19.865 145.905 20.035 146.115 ;
        RECT 21.245 145.905 21.415 146.095 ;
        RECT 21.760 145.955 21.880 146.065 ;
        RECT 23.730 145.925 23.900 146.115 ;
        RECT 24.980 145.955 25.100 146.065 ;
        RECT 25.385 145.925 25.555 146.115 ;
        RECT 27.685 145.925 27.855 146.115 ;
        RECT 28.145 145.925 28.315 146.115 ;
        RECT 29.800 145.925 29.970 146.115 ;
        RECT 31.365 145.905 31.535 146.095 ;
        RECT 33.720 145.955 33.840 146.065 ;
        RECT 35.505 145.925 35.675 146.115 ;
        RECT 36.885 145.905 37.055 146.095 ;
        RECT 37.860 145.955 37.980 146.065 ;
        RECT 39.180 145.925 39.350 146.115 ;
        RECT 39.650 145.925 39.820 146.115 ;
        RECT 40.565 145.905 40.735 146.095 ;
        RECT 41.025 145.905 41.195 146.095 ;
        RECT 42.405 145.905 42.575 146.095 ;
        RECT 44.245 145.925 44.415 146.115 ;
        RECT 49.765 145.925 49.935 146.115 ;
        RECT 51.145 145.960 51.305 146.070 ;
        RECT 51.880 145.925 52.050 146.115 ;
        RECT 52.985 145.905 53.155 146.095 ;
        RECT 54.365 145.905 54.535 146.095 ;
        RECT 55.750 145.925 55.920 146.115 ;
        RECT 58.045 145.905 58.215 146.095 ;
        RECT 58.505 145.905 58.675 146.095 ;
        RECT 59.480 145.955 59.600 146.065 ;
        RECT 59.940 145.955 60.060 146.065 ;
        RECT 62.645 145.905 62.815 146.095 ;
        RECT 63.290 145.925 63.460 146.115 ;
        RECT 63.620 145.955 63.740 146.065 ;
        RECT 64.945 145.925 65.115 146.115 ;
        RECT 67.430 145.905 67.600 146.095 ;
        RECT 68.220 145.955 68.340 146.065 ;
        RECT 70.465 145.925 70.635 146.115 ;
        RECT 72.305 145.925 72.475 146.115 ;
        RECT 72.765 145.925 72.935 146.115 ;
        RECT 73.685 145.905 73.855 146.095 ;
        RECT 75.525 145.925 75.695 146.115 ;
        RECT 79.660 146.095 79.830 146.115 ;
        RECT 79.205 145.905 79.375 146.095 ;
        RECT 79.660 145.925 79.840 146.095 ;
        RECT 80.130 145.925 80.300 146.115 ;
        RECT 82.480 145.955 82.600 146.065 ;
        RECT 14.665 145.095 16.035 145.905 ;
        RECT 16.505 145.095 20.175 145.905 ;
        RECT 20.195 144.995 21.545 145.905 ;
        RECT 22.395 145.225 31.675 145.905 ;
        RECT 22.395 145.105 24.730 145.225 ;
        RECT 22.395 144.995 23.315 145.105 ;
        RECT 29.395 145.005 30.315 145.225 ;
        RECT 31.685 145.095 37.195 145.905 ;
        RECT 38.125 145.095 40.875 145.905 ;
        RECT 40.895 144.995 42.245 145.905 ;
        RECT 42.265 145.225 51.545 145.905 ;
        RECT 43.625 145.005 44.545 145.225 ;
        RECT 49.210 145.105 51.545 145.225 ;
        RECT 51.925 145.125 53.295 145.905 ;
        RECT 50.625 144.995 51.545 145.105 ;
        RECT 53.305 145.095 54.675 145.905 ;
        RECT 54.685 145.095 58.355 145.905 ;
        RECT 58.375 144.995 59.725 145.905 ;
        RECT 60.205 145.095 62.955 145.905 ;
        RECT 64.115 145.225 68.015 145.905 ;
        RECT 67.085 144.995 68.015 145.225 ;
        RECT 68.485 145.095 73.995 145.905 ;
        RECT 74.005 145.095 79.515 145.905 ;
        RECT 79.670 145.875 79.840 145.925 ;
        RECT 84.265 145.905 84.435 146.095 ;
        RECT 84.725 145.925 84.895 146.115 ;
        RECT 88.130 145.905 88.300 146.095 ;
        RECT 89.785 145.950 89.945 146.060 ;
        RECT 90.245 145.905 90.415 146.095 ;
        RECT 92.545 145.905 92.715 146.095 ;
        RECT 93.005 145.905 93.175 146.095 ;
        RECT 94.385 145.925 94.555 146.115 ;
        RECT 95.305 145.960 95.465 146.070 ;
        RECT 95.765 145.925 95.935 146.115 ;
        RECT 100.550 145.925 100.720 146.115 ;
        RECT 101.340 145.955 101.460 146.065 ;
        RECT 102.205 145.925 102.375 146.115 ;
        RECT 103.640 145.955 103.760 146.065 ;
        RECT 105.425 145.905 105.595 146.095 ;
        RECT 105.940 145.955 106.060 146.065 ;
        RECT 106.340 145.925 106.510 146.145 ;
        RECT 106.665 146.115 110.140 147.025 ;
        RECT 110.345 146.115 112.175 146.925 ;
        RECT 115.385 146.795 116.315 147.025 ;
        RECT 112.415 146.115 116.315 146.795 ;
        RECT 116.695 146.915 117.615 147.025 ;
        RECT 116.695 146.795 119.030 146.915 ;
        RECT 123.695 146.795 124.615 147.015 ;
        RECT 116.695 146.115 125.975 146.795 ;
        RECT 126.445 146.115 127.815 146.925 ;
        RECT 106.810 145.925 106.980 146.115 ;
        RECT 109.565 145.905 109.735 146.095 ;
        RECT 111.865 145.925 112.035 146.115 ;
        RECT 113.240 145.905 113.410 146.095 ;
        RECT 114.165 145.950 114.325 146.060 ;
        RECT 115.140 145.955 115.260 146.065 ;
        RECT 115.730 145.925 115.900 146.115 ;
        RECT 118.950 145.905 119.120 146.095 ;
        RECT 119.685 145.905 119.855 146.095 ;
        RECT 121.120 145.955 121.240 146.065 ;
        RECT 121.525 145.905 121.695 146.095 ;
        RECT 125.665 145.925 125.835 146.115 ;
        RECT 126.125 146.065 126.295 146.095 ;
        RECT 126.125 145.955 126.300 146.065 ;
        RECT 126.125 145.905 126.295 145.955 ;
        RECT 127.505 145.905 127.675 146.115 ;
        RECT 81.330 145.875 82.275 145.905 ;
        RECT 79.525 145.195 82.275 145.875 ;
        RECT 81.330 144.995 82.275 145.195 ;
        RECT 82.745 145.095 84.575 145.905 ;
        RECT 84.815 145.225 88.715 145.905 ;
        RECT 87.785 144.995 88.715 145.225 ;
        RECT 90.105 145.125 91.475 145.905 ;
        RECT 91.485 145.125 92.855 145.905 ;
        RECT 92.975 145.225 96.440 145.905 ;
        RECT 95.520 144.995 96.440 145.225 ;
        RECT 96.545 145.225 105.735 145.905 ;
        RECT 96.545 144.995 97.465 145.225 ;
        RECT 100.295 145.005 101.225 145.225 ;
        RECT 106.205 145.095 109.875 145.905 ;
        RECT 110.080 144.995 113.555 145.905 ;
        RECT 115.635 145.225 119.535 145.905 ;
        RECT 118.605 144.995 119.535 145.225 ;
        RECT 119.555 144.995 120.905 145.905 ;
        RECT 121.385 145.125 122.755 145.905 ;
        RECT 122.765 145.095 126.435 145.905 ;
        RECT 126.445 145.095 127.815 145.905 ;
        RECT 14.665 140.675 16.035 141.485 ;
        RECT 16.045 140.675 18.795 141.485 ;
        RECT 18.805 140.675 24.315 141.485 ;
        RECT 25.245 140.675 28.915 141.485 ;
        RECT 28.925 140.675 34.435 141.485 ;
        RECT 34.445 141.385 35.390 141.585 ;
        RECT 34.445 140.705 37.195 141.385 ;
        RECT 34.445 140.675 35.390 140.705 ;
        RECT 14.805 140.465 14.975 140.675 ;
        RECT 18.485 140.485 18.655 140.675 ;
        RECT 24.005 140.485 24.175 140.675 ;
        RECT 24.980 140.515 25.100 140.625 ;
        RECT 25.385 140.465 25.555 140.655 ;
        RECT 28.145 140.465 28.315 140.655 ;
        RECT 28.605 140.485 28.775 140.675 ;
        RECT 33.665 140.465 33.835 140.655 ;
        RECT 34.125 140.485 34.295 140.675 ;
        RECT 36.880 140.485 37.050 140.705 ;
        RECT 38.125 140.675 41.795 141.485 ;
        RECT 41.805 140.675 47.315 141.485 ;
        RECT 49.130 141.385 50.075 141.585 ;
        RECT 47.325 140.705 50.075 141.385 ;
        RECT 37.805 140.520 37.965 140.630 ;
        RECT 38.265 140.510 38.425 140.620 ;
        RECT 34.145 140.465 34.295 140.485 ;
        RECT 14.665 139.655 16.035 140.465 ;
        RECT 16.415 139.785 25.695 140.465 ;
        RECT 16.415 139.665 18.750 139.785 ;
        RECT 16.415 139.555 17.335 139.665 ;
        RECT 23.415 139.565 24.335 139.785 ;
        RECT 25.705 139.655 28.455 140.465 ;
        RECT 28.465 139.655 33.975 140.465 ;
        RECT 34.145 139.645 36.075 140.465 ;
        RECT 35.125 139.555 36.075 139.645 ;
        RECT 38.585 140.435 39.530 140.465 ;
        RECT 41.020 140.435 41.190 140.655 ;
        RECT 41.485 140.485 41.655 140.675 ;
        RECT 47.005 140.655 47.175 140.675 ;
        RECT 46.545 140.465 46.715 140.655 ;
        RECT 47.005 140.485 47.180 140.655 ;
        RECT 47.470 140.485 47.640 140.705 ;
        RECT 49.130 140.675 50.075 140.705 ;
        RECT 50.545 140.675 52.375 141.485 ;
        RECT 52.385 140.675 55.860 141.585 ;
        RECT 58.720 141.355 59.640 141.585 ;
        RECT 56.175 140.675 59.640 141.355 ;
        RECT 59.745 141.355 60.665 141.585 ;
        RECT 63.495 141.355 64.425 141.575 ;
        RECT 59.745 140.675 68.935 141.355 ;
        RECT 68.945 140.675 70.315 141.455 ;
        RECT 70.325 140.675 71.695 141.485 ;
        RECT 71.715 140.675 73.065 141.585 ;
        RECT 73.085 140.675 75.835 141.485 ;
        RECT 76.765 140.675 79.515 141.485 ;
        RECT 79.525 140.675 85.035 141.485 ;
        RECT 85.045 140.675 90.555 141.485 ;
        RECT 90.565 140.675 96.075 141.485 ;
        RECT 96.085 140.675 101.595 141.485 ;
        RECT 102.985 140.675 108.495 141.485 ;
        RECT 110.310 141.385 111.255 141.585 ;
        RECT 108.505 140.705 111.255 141.385 ;
        RECT 38.585 139.755 41.335 140.435 ;
        RECT 38.585 139.555 39.530 139.755 ;
        RECT 41.345 139.655 46.855 140.465 ;
        RECT 47.010 140.435 47.180 140.485 ;
        RECT 49.770 140.465 49.940 140.655 ;
        RECT 52.065 140.485 52.235 140.675 ;
        RECT 52.530 140.485 52.700 140.675 ;
        RECT 54.825 140.465 54.995 140.655 ;
        RECT 55.285 140.465 55.455 140.655 ;
        RECT 56.205 140.485 56.375 140.675 ;
        RECT 58.965 140.465 59.135 140.655 ;
        RECT 59.430 140.465 59.600 140.655 ;
        RECT 63.620 140.515 63.740 140.625 ;
        RECT 64.030 140.465 64.200 140.655 ;
        RECT 67.705 140.465 67.875 140.655 ;
        RECT 68.625 140.485 68.795 140.675 ;
        RECT 70.005 140.485 70.175 140.675 ;
        RECT 71.385 140.485 71.555 140.675 ;
        RECT 71.845 140.485 72.015 140.675 ;
        RECT 75.525 140.485 75.695 140.675 ;
        RECT 76.500 140.515 76.620 140.625 ;
        RECT 79.205 140.485 79.375 140.675 ;
        RECT 79.665 140.465 79.835 140.655 ;
        RECT 80.130 140.465 80.300 140.655 ;
        RECT 84.265 140.510 84.425 140.620 ;
        RECT 84.725 140.485 84.895 140.675 ;
        RECT 88.130 140.465 88.300 140.655 ;
        RECT 89.380 140.515 89.500 140.625 ;
        RECT 89.785 140.465 89.955 140.655 ;
        RECT 90.245 140.485 90.415 140.675 ;
        RECT 91.625 140.510 91.785 140.620 ;
        RECT 95.305 140.465 95.475 140.655 ;
        RECT 95.765 140.485 95.935 140.675 ;
        RECT 100.825 140.465 100.995 140.655 ;
        RECT 101.285 140.465 101.455 140.675 ;
        RECT 102.665 140.520 102.825 140.630 ;
        RECT 105.885 140.465 106.055 140.655 ;
        RECT 106.350 140.465 106.520 140.655 ;
        RECT 108.185 140.485 108.355 140.675 ;
        RECT 108.650 140.485 108.820 140.705 ;
        RECT 110.310 140.675 111.255 140.705 ;
        RECT 112.185 140.675 115.855 141.485 ;
        RECT 119.065 141.355 119.995 141.585 ;
        RECT 116.095 140.675 119.995 141.355 ;
        RECT 120.015 140.675 121.365 141.585 ;
        RECT 121.385 140.675 122.755 141.485 ;
        RECT 122.765 140.675 126.435 141.485 ;
        RECT 126.445 140.675 127.815 141.485 ;
        RECT 111.865 140.520 112.025 140.630 ;
        RECT 113.240 140.465 113.410 140.655 ;
        RECT 114.165 140.510 114.325 140.620 ;
        RECT 115.140 140.515 115.260 140.625 ;
        RECT 115.545 140.465 115.715 140.675 ;
        RECT 119.410 140.485 119.580 140.675 ;
        RECT 120.145 140.485 120.315 140.675 ;
        RECT 122.445 140.485 122.615 140.675 ;
        RECT 126.125 140.465 126.295 140.675 ;
        RECT 127.505 140.465 127.675 140.675 ;
        RECT 48.670 140.435 49.615 140.465 ;
        RECT 46.865 139.755 49.615 140.435 ;
        RECT 48.670 139.555 49.615 139.755 ;
        RECT 49.625 139.555 53.100 140.465 ;
        RECT 53.305 139.655 55.135 140.465 ;
        RECT 55.155 139.555 56.505 140.465 ;
        RECT 56.525 139.655 59.275 140.465 ;
        RECT 59.285 139.555 62.760 140.465 ;
        RECT 63.885 139.555 67.360 140.465 ;
        RECT 67.565 139.785 76.845 140.465 ;
        RECT 68.925 139.565 69.845 139.785 ;
        RECT 74.510 139.665 76.845 139.785 ;
        RECT 75.925 139.555 76.845 139.665 ;
        RECT 77.225 139.655 79.975 140.465 ;
        RECT 79.985 139.555 83.460 140.465 ;
        RECT 84.815 139.785 88.715 140.465 ;
        RECT 87.785 139.555 88.715 139.785 ;
        RECT 89.645 139.685 91.015 140.465 ;
        RECT 91.945 139.655 95.615 140.465 ;
        RECT 95.625 139.655 101.135 140.465 ;
        RECT 101.155 139.555 102.505 140.465 ;
        RECT 102.525 139.655 106.195 140.465 ;
        RECT 106.205 139.555 109.680 140.465 ;
        RECT 110.080 139.555 113.555 140.465 ;
        RECT 115.415 139.555 116.765 140.465 ;
        RECT 117.155 139.785 126.435 140.465 ;
        RECT 117.155 139.665 119.490 139.785 ;
        RECT 117.155 139.555 118.075 139.665 ;
        RECT 124.155 139.565 125.075 139.785 ;
        RECT 126.445 139.655 127.815 140.465 ;
        RECT 14.665 135.235 16.035 136.045 ;
        RECT 16.045 135.235 21.555 136.045 ;
        RECT 21.565 135.235 22.935 136.015 ;
        RECT 22.955 135.235 24.305 136.145 ;
        RECT 25.245 135.235 28.915 136.045 ;
        RECT 32.125 135.915 33.055 136.145 ;
        RECT 29.155 135.235 33.055 135.915 ;
        RECT 33.065 135.235 34.895 136.045 ;
        RECT 34.905 135.945 35.850 136.145 ;
        RECT 38.805 136.055 39.755 136.145 ;
        RECT 34.905 135.265 37.655 135.945 ;
        RECT 34.905 135.235 35.850 135.265 ;
        RECT 14.805 135.025 14.975 135.235 ;
        RECT 17.105 135.025 17.275 135.215 ;
        RECT 20.970 135.025 21.140 135.215 ;
        RECT 21.245 135.045 21.415 135.235 ;
        RECT 21.705 135.045 21.875 135.235 ;
        RECT 23.085 135.045 23.255 135.235 ;
        RECT 24.980 135.075 25.100 135.185 ;
        RECT 28.605 135.045 28.775 135.235 ;
        RECT 30.905 135.025 31.075 135.215 ;
        RECT 32.285 135.025 32.455 135.215 ;
        RECT 32.470 135.045 32.640 135.235 ;
        RECT 32.800 135.075 32.920 135.185 ;
        RECT 34.585 135.045 34.755 135.235 ;
        RECT 36.610 135.025 36.780 135.215 ;
        RECT 37.340 135.045 37.510 135.265 ;
        RECT 37.825 135.235 39.755 136.055 ;
        RECT 39.965 135.235 43.635 136.045 ;
        RECT 43.645 135.945 44.590 136.145 ;
        RECT 43.645 135.265 46.395 135.945 ;
        RECT 43.645 135.235 44.590 135.265 ;
        RECT 37.825 135.215 37.975 135.235 ;
        RECT 37.805 135.045 37.975 135.215 ;
        RECT 14.665 134.215 16.035 135.025 ;
        RECT 16.055 134.115 17.405 135.025 ;
        RECT 17.655 134.345 21.555 135.025 ;
        RECT 20.625 134.115 21.555 134.345 ;
        RECT 21.935 134.345 31.215 135.025 ;
        RECT 21.935 134.225 24.270 134.345 ;
        RECT 21.935 134.115 22.855 134.225 ;
        RECT 28.935 134.125 29.855 134.345 ;
        RECT 31.225 134.245 32.595 135.025 ;
        RECT 33.295 134.345 37.195 135.025 ;
        RECT 36.265 134.115 37.195 134.345 ;
        RECT 37.665 134.995 38.610 135.025 ;
        RECT 40.100 134.995 40.270 135.215 ;
        RECT 41.485 135.025 41.655 135.215 ;
        RECT 37.665 134.315 40.415 134.995 ;
        RECT 37.665 134.115 38.610 134.315 ;
        RECT 40.425 134.215 41.795 135.025 ;
        RECT 41.950 134.995 42.120 135.215 ;
        RECT 43.325 135.045 43.495 135.235 ;
        RECT 44.710 135.025 44.880 135.215 ;
        RECT 46.080 135.045 46.250 135.265 ;
        RECT 46.405 135.235 50.075 136.045 ;
        RECT 51.005 135.235 52.835 136.045 ;
        RECT 56.045 135.915 56.975 136.145 ;
        RECT 53.075 135.235 56.975 135.915 ;
        RECT 57.445 135.235 58.815 136.015 ;
        RECT 59.285 135.235 61.115 136.045 ;
        RECT 61.125 135.235 64.600 136.145 ;
        RECT 65.265 135.235 67.095 136.045 ;
        RECT 67.105 135.235 70.315 136.145 ;
        RECT 70.420 135.915 71.340 136.145 ;
        RECT 70.420 135.235 73.885 135.915 ;
        RECT 74.005 135.235 75.835 136.045 ;
        RECT 77.225 135.945 78.170 136.145 ;
        RECT 77.225 135.265 79.975 135.945 ;
        RECT 77.225 135.235 78.170 135.265 ;
        RECT 48.390 135.025 48.560 135.215 ;
        RECT 49.765 135.045 49.935 135.235 ;
        RECT 50.740 135.075 50.860 135.185 ;
        RECT 52.525 135.045 52.695 135.235 ;
        RECT 56.390 135.045 56.560 135.235 ;
        RECT 57.180 135.075 57.300 135.185 ;
        RECT 57.585 135.045 57.755 135.235 ;
        RECT 59.020 135.075 59.140 135.185 ;
        RECT 60.805 135.045 60.975 135.235 ;
        RECT 61.270 135.215 61.440 135.235 ;
        RECT 61.265 135.045 61.440 135.215 ;
        RECT 61.265 135.025 61.435 135.045 ;
        RECT 62.645 135.025 62.815 135.215 ;
        RECT 63.570 135.025 63.740 135.215 ;
        RECT 65.000 135.075 65.120 135.185 ;
        RECT 66.785 135.045 66.955 135.235 ;
        RECT 67.705 135.070 67.865 135.180 ;
        RECT 70.005 135.045 70.175 135.235 ;
        RECT 73.225 135.025 73.395 135.215 ;
        RECT 73.685 135.045 73.855 135.235 ;
        RECT 75.525 135.045 75.695 135.235 ;
        RECT 76.905 135.080 77.065 135.190 ;
        RECT 78.745 135.025 78.915 135.215 ;
        RECT 43.610 134.995 44.555 135.025 ;
        RECT 41.805 134.315 44.555 134.995 ;
        RECT 43.610 134.115 44.555 134.315 ;
        RECT 44.565 134.115 48.040 135.025 ;
        RECT 48.245 134.115 51.720 135.025 ;
        RECT 52.295 134.345 61.575 135.025 ;
        RECT 52.295 134.225 54.630 134.345 ;
        RECT 52.295 134.115 53.215 134.225 ;
        RECT 59.295 134.125 60.215 134.345 ;
        RECT 61.585 134.215 62.955 135.025 ;
        RECT 63.425 134.115 66.900 135.025 ;
        RECT 68.025 134.215 73.535 135.025 ;
        RECT 73.545 134.215 79.055 135.025 ;
        RECT 79.210 134.995 79.380 135.215 ;
        RECT 79.660 135.045 79.830 135.265 ;
        RECT 79.985 135.235 83.460 136.145 ;
        RECT 84.035 136.035 84.955 136.145 ;
        RECT 84.035 135.915 86.370 136.035 ;
        RECT 91.035 135.915 91.955 136.135 ;
        RECT 96.525 135.915 97.455 136.145 ;
        RECT 84.035 135.235 93.315 135.915 ;
        RECT 93.555 135.235 97.455 135.915 ;
        RECT 98.120 135.235 101.595 136.145 ;
        RECT 106.185 135.915 107.115 136.145 ;
        RECT 103.215 135.235 107.115 135.915 ;
        RECT 107.125 135.235 108.495 136.015 ;
        RECT 112.625 135.915 113.555 136.145 ;
        RECT 109.655 135.235 113.555 135.915 ;
        RECT 113.935 136.035 114.855 136.145 ;
        RECT 113.935 135.915 116.270 136.035 ;
        RECT 120.935 135.915 121.855 136.135 ;
        RECT 113.935 135.235 123.215 135.915 ;
        RECT 123.225 135.235 124.595 136.015 ;
        RECT 124.605 135.235 126.435 136.045 ;
        RECT 126.445 135.235 127.815 136.045 ;
        RECT 80.130 135.045 80.300 135.235 ;
        RECT 87.025 135.025 87.195 135.215 ;
        RECT 88.405 135.025 88.575 135.215 ;
        RECT 93.005 135.045 93.175 135.235 ;
        RECT 96.870 135.045 97.040 135.235 ;
        RECT 97.660 135.075 97.780 135.185 ;
        RECT 98.525 135.025 98.695 135.215 ;
        RECT 101.280 135.045 101.450 135.235 ;
        RECT 102.665 135.080 102.825 135.190 ;
        RECT 106.530 135.045 106.700 135.235 ;
        RECT 108.185 135.025 108.355 135.235 ;
        RECT 80.870 134.995 81.815 135.025 ;
        RECT 79.065 134.315 81.815 134.995 ;
        RECT 80.870 134.115 81.815 134.315 ;
        RECT 81.825 134.215 87.335 135.025 ;
        RECT 87.355 134.115 88.705 135.025 ;
        RECT 89.555 134.345 98.835 135.025 ;
        RECT 99.215 134.345 108.495 135.025 ;
        RECT 108.650 134.995 108.820 135.215 ;
        RECT 109.105 135.080 109.265 135.190 ;
        RECT 111.460 135.075 111.580 135.185 ;
        RECT 112.970 135.045 113.140 135.235 ;
        RECT 114.165 135.025 114.335 135.215 ;
        RECT 115.140 135.075 115.260 135.185 ;
        RECT 118.765 135.025 118.935 135.215 ;
        RECT 119.225 135.025 119.395 135.215 ;
        RECT 120.660 135.075 120.780 135.185 ;
        RECT 122.905 135.045 123.075 135.235 ;
        RECT 123.365 135.045 123.535 135.235 ;
        RECT 126.125 135.025 126.295 135.235 ;
        RECT 127.505 135.025 127.675 135.235 ;
        RECT 110.310 134.995 111.255 135.025 ;
        RECT 89.555 134.225 91.890 134.345 ;
        RECT 89.555 134.115 90.475 134.225 ;
        RECT 96.555 134.125 97.475 134.345 ;
        RECT 99.215 134.225 101.550 134.345 ;
        RECT 99.215 134.115 100.135 134.225 ;
        RECT 106.215 134.125 107.135 134.345 ;
        RECT 108.505 134.315 111.255 134.995 ;
        RECT 110.310 134.115 111.255 134.315 ;
        RECT 111.725 134.215 114.475 135.025 ;
        RECT 115.405 134.215 119.075 135.025 ;
        RECT 119.085 134.245 120.455 135.025 ;
        RECT 120.925 134.215 126.435 135.025 ;
        RECT 126.445 134.215 127.815 135.025 ;
        RECT 14.665 129.795 16.035 130.605 ;
        RECT 16.505 129.795 20.175 130.605 ;
        RECT 23.385 130.475 24.315 130.705 ;
        RECT 20.415 129.795 24.315 130.475 ;
        RECT 24.785 129.795 30.295 130.605 ;
        RECT 30.675 130.595 31.595 130.705 ;
        RECT 30.675 130.475 33.010 130.595 ;
        RECT 37.675 130.475 38.595 130.695 ;
        RECT 43.865 130.615 44.815 130.705 ;
        RECT 46.165 130.615 47.115 130.705 ;
        RECT 30.675 129.795 39.955 130.475 ;
        RECT 39.965 129.795 41.335 130.575 ;
        RECT 41.345 129.795 42.715 130.605 ;
        RECT 42.885 129.795 44.815 130.615 ;
        RECT 45.185 129.795 47.115 130.615 ;
        RECT 47.325 129.795 50.075 130.605 ;
        RECT 50.545 129.795 54.215 130.605 ;
        RECT 54.225 129.795 59.735 130.605 ;
        RECT 59.745 129.795 65.255 130.605 ;
        RECT 68.465 130.475 69.395 130.705 ;
        RECT 71.905 130.615 72.855 130.705 ;
        RECT 78.805 130.615 79.755 130.705 ;
        RECT 65.495 129.795 69.395 130.475 ;
        RECT 69.865 129.795 71.695 130.475 ;
        RECT 71.905 129.795 73.835 130.615 ;
        RECT 74.005 129.795 75.835 130.475 ;
        RECT 76.765 129.795 78.595 130.605 ;
        RECT 78.805 129.795 80.735 130.615 ;
        RECT 80.905 129.795 82.275 130.605 ;
        RECT 82.285 129.795 87.795 130.605 ;
        RECT 87.815 129.795 89.165 130.705 ;
        RECT 92.385 130.475 93.315 130.705 ;
        RECT 89.415 129.795 93.315 130.475 ;
        RECT 93.785 129.795 95.155 130.575 ;
        RECT 95.165 129.795 96.535 130.575 ;
        RECT 96.545 129.795 97.915 130.605 ;
        RECT 97.925 130.505 98.870 130.705 ;
        RECT 97.925 129.825 100.675 130.505 ;
        RECT 97.925 129.795 98.870 129.825 ;
        RECT 14.805 129.585 14.975 129.795 ;
        RECT 16.240 129.635 16.360 129.745 ;
        RECT 16.645 129.630 16.805 129.740 ;
        RECT 19.865 129.605 20.035 129.795 ;
        RECT 23.730 129.605 23.900 129.795 ;
        RECT 26.305 129.585 26.475 129.775 ;
        RECT 27.685 129.585 27.855 129.775 ;
        RECT 29.985 129.605 30.155 129.795 ;
        RECT 33.205 129.585 33.375 129.775 ;
        RECT 33.665 129.585 33.835 129.775 ;
        RECT 35.045 129.605 35.215 129.775 ;
        RECT 37.860 129.635 37.980 129.745 ;
        RECT 39.645 129.605 39.815 129.795 ;
        RECT 35.065 129.585 35.215 129.605 ;
        RECT 40.565 129.585 40.735 129.775 ;
        RECT 41.025 129.605 41.195 129.795 ;
        RECT 42.405 129.605 42.575 129.795 ;
        RECT 42.885 129.775 43.035 129.795 ;
        RECT 45.185 129.775 45.335 129.795 ;
        RECT 42.865 129.605 43.035 129.775 ;
        RECT 45.165 129.605 45.335 129.775 ;
        RECT 46.085 129.585 46.255 129.775 ;
        RECT 46.545 129.605 46.715 129.775 ;
        RECT 48.900 129.635 49.020 129.745 ;
        RECT 49.765 129.605 49.935 129.795 ;
        RECT 53.905 129.605 54.075 129.795 ;
        RECT 46.565 129.585 46.715 129.605 ;
        RECT 54.365 129.585 54.535 129.775 ;
        RECT 58.230 129.585 58.400 129.775 ;
        RECT 58.965 129.585 59.135 129.775 ;
        RECT 59.425 129.605 59.595 129.795 ;
        RECT 62.645 129.585 62.815 129.775 ;
        RECT 64.485 129.585 64.655 129.775 ;
        RECT 64.945 129.605 65.115 129.795 ;
        RECT 68.810 129.605 68.980 129.795 ;
        RECT 69.600 129.635 69.720 129.745 ;
        RECT 71.385 129.605 71.555 129.795 ;
        RECT 73.685 129.775 73.835 129.795 ;
        RECT 73.685 129.605 73.855 129.775 ;
        RECT 74.145 129.585 74.315 129.795 ;
        RECT 74.605 129.605 74.775 129.775 ;
        RECT 76.500 129.635 76.620 129.745 ;
        RECT 76.905 129.605 77.075 129.775 ;
        RECT 78.285 129.605 78.455 129.795 ;
        RECT 80.585 129.775 80.735 129.795 ;
        RECT 80.585 129.605 80.755 129.775 ;
        RECT 81.965 129.605 82.135 129.795 ;
        RECT 74.625 129.585 74.775 129.605 ;
        RECT 76.925 129.585 77.075 129.605 ;
        RECT 82.610 129.585 82.780 129.775 ;
        RECT 85.185 129.605 85.355 129.775 ;
        RECT 85.700 129.635 85.820 129.745 ;
        RECT 87.485 129.605 87.655 129.795 ;
        RECT 87.945 129.605 88.115 129.795 ;
        RECT 85.185 129.585 85.335 129.605 ;
        RECT 88.405 129.585 88.575 129.775 ;
        RECT 89.380 129.635 89.500 129.745 ;
        RECT 92.730 129.605 92.900 129.795 ;
        RECT 93.520 129.635 93.640 129.745 ;
        RECT 93.925 129.605 94.095 129.795 ;
        RECT 95.305 129.605 95.475 129.795 ;
        RECT 97.605 129.605 97.775 129.795 ;
        RECT 98.985 129.585 99.155 129.775 ;
        RECT 99.445 129.605 99.615 129.775 ;
        RECT 100.360 129.605 100.530 129.825 ;
        RECT 102.065 129.795 103.895 130.605 ;
        RECT 105.710 130.505 106.655 130.705 ;
        RECT 110.545 130.615 111.495 130.705 ;
        RECT 103.905 129.825 106.655 130.505 ;
        RECT 101.285 129.640 101.445 129.750 ;
        RECT 103.585 129.605 103.755 129.795 ;
        RECT 104.050 129.775 104.220 129.825 ;
        RECT 105.710 129.795 106.655 129.825 ;
        RECT 106.665 129.795 110.335 130.605 ;
        RECT 110.545 129.795 112.475 130.615 ;
        RECT 112.645 129.795 115.395 130.605 ;
        RECT 115.405 129.795 120.915 130.605 ;
        RECT 120.925 129.795 126.435 130.605 ;
        RECT 126.445 129.795 127.815 130.605 ;
        RECT 104.045 129.605 104.220 129.775 ;
        RECT 106.345 129.605 106.515 129.775 ;
        RECT 108.645 129.605 108.815 129.775 ;
        RECT 110.025 129.605 110.195 129.795 ;
        RECT 112.325 129.775 112.475 129.795 ;
        RECT 110.945 129.605 111.115 129.775 ;
        RECT 111.460 129.635 111.580 129.745 ;
        RECT 112.325 129.605 112.495 129.775 ;
        RECT 99.465 129.585 99.615 129.605 ;
        RECT 104.045 129.585 104.215 129.605 ;
        RECT 106.345 129.585 106.495 129.605 ;
        RECT 108.645 129.585 108.795 129.605 ;
        RECT 110.945 129.585 111.095 129.605 ;
        RECT 114.165 129.585 114.335 129.775 ;
        RECT 115.085 129.605 115.255 129.795 ;
        RECT 116.925 129.605 117.095 129.775 ;
        RECT 117.845 129.630 118.005 129.740 ;
        RECT 116.925 129.585 117.075 129.605 ;
        RECT 118.305 129.585 118.475 129.775 ;
        RECT 119.740 129.635 119.860 129.745 ;
        RECT 120.145 129.585 120.315 129.775 ;
        RECT 120.605 129.605 120.775 129.795 ;
        RECT 122.445 129.585 122.615 129.775 ;
        RECT 126.125 129.585 126.295 129.795 ;
        RECT 127.505 129.585 127.675 129.795 ;
        RECT 14.665 128.775 16.035 129.585 ;
        RECT 17.335 128.905 26.615 129.585 ;
        RECT 17.335 128.785 19.670 128.905 ;
        RECT 17.335 128.675 18.255 128.785 ;
        RECT 24.335 128.685 25.255 128.905 ;
        RECT 26.625 128.775 27.995 129.585 ;
        RECT 28.005 128.775 33.515 129.585 ;
        RECT 33.535 128.675 34.885 129.585 ;
        RECT 35.065 128.765 36.995 129.585 ;
        RECT 38.125 128.775 40.875 129.585 ;
        RECT 40.885 128.775 46.395 129.585 ;
        RECT 46.565 128.765 48.495 129.585 ;
        RECT 49.165 128.775 54.675 129.585 ;
        RECT 54.915 128.905 58.815 129.585 ;
        RECT 36.045 128.675 36.995 128.765 ;
        RECT 47.545 128.675 48.495 128.765 ;
        RECT 57.885 128.675 58.815 128.905 ;
        RECT 58.825 128.805 60.195 129.585 ;
        RECT 60.205 128.775 62.955 129.585 ;
        RECT 63.425 128.775 64.795 129.585 ;
        RECT 65.175 128.905 74.455 129.585 ;
        RECT 65.175 128.785 67.510 128.905 ;
        RECT 65.175 128.675 66.095 128.785 ;
        RECT 72.175 128.685 73.095 128.905 ;
        RECT 74.625 128.765 76.555 129.585 ;
        RECT 76.925 128.765 78.855 129.585 ;
        RECT 79.295 128.905 83.195 129.585 ;
        RECT 75.605 128.675 76.555 128.765 ;
        RECT 77.905 128.675 78.855 128.765 ;
        RECT 82.265 128.675 83.195 128.905 ;
        RECT 83.405 128.765 85.335 129.585 ;
        RECT 85.965 128.775 88.715 129.585 ;
        RECT 90.015 128.905 99.295 129.585 ;
        RECT 90.015 128.785 92.350 128.905 ;
        RECT 83.405 128.675 84.355 128.765 ;
        RECT 90.015 128.675 90.935 128.785 ;
        RECT 97.015 128.685 97.935 128.905 ;
        RECT 99.465 128.765 101.395 129.585 ;
        RECT 101.605 128.775 104.355 129.585 ;
        RECT 100.445 128.675 101.395 128.765 ;
        RECT 104.565 128.765 106.495 129.585 ;
        RECT 106.865 128.765 108.795 129.585 ;
        RECT 109.165 128.765 111.095 129.585 ;
        RECT 111.735 128.905 114.475 129.585 ;
        RECT 115.145 128.765 117.075 129.585 ;
        RECT 104.565 128.675 105.515 128.765 ;
        RECT 106.865 128.675 107.815 128.765 ;
        RECT 109.165 128.675 110.115 128.765 ;
        RECT 115.145 128.675 116.095 128.765 ;
        RECT 118.175 128.675 119.525 129.585 ;
        RECT 120.005 128.805 121.375 129.585 ;
        RECT 121.385 128.775 122.755 129.585 ;
        RECT 122.765 128.775 126.435 129.585 ;
        RECT 126.445 128.775 127.815 129.585 ;
        RECT 14.665 124.355 16.035 125.165 ;
        RECT 16.965 124.355 20.635 125.165 ;
        RECT 20.655 124.355 22.005 125.265 ;
        RECT 22.945 124.355 24.315 125.135 ;
        RECT 24.785 124.355 26.155 125.165 ;
        RECT 26.165 125.035 27.095 125.265 ;
        RECT 26.165 124.355 30.065 125.035 ;
        RECT 30.305 124.355 33.055 125.165 ;
        RECT 36.265 125.035 37.195 125.265 ;
        RECT 38.345 125.175 39.295 125.265 ;
        RECT 41.565 125.175 42.515 125.265 ;
        RECT 43.865 125.175 44.815 125.265 ;
        RECT 33.295 124.355 37.195 125.035 ;
        RECT 37.365 124.355 39.295 125.175 ;
        RECT 40.585 124.355 42.515 125.175 ;
        RECT 42.885 124.355 44.815 125.175 ;
        RECT 45.225 125.175 46.175 125.265 ;
        RECT 45.225 124.355 47.155 125.175 ;
        RECT 63.405 125.035 64.335 125.265 ;
        RECT 47.335 124.355 50.075 125.035 ;
        RECT 51.005 124.355 60.110 125.035 ;
        RECT 60.435 124.355 64.335 125.035 ;
        RECT 64.805 124.355 68.475 125.165 ;
        RECT 68.495 124.355 69.845 125.265 ;
        RECT 69.865 124.355 71.235 125.135 ;
        RECT 71.245 124.355 72.615 125.165 ;
        RECT 76.675 125.155 77.595 125.265 ;
        RECT 76.675 125.035 79.010 125.155 ;
        RECT 83.675 125.035 84.595 125.255 ;
        RECT 72.625 124.355 75.365 125.035 ;
        RECT 76.675 124.355 85.955 125.035 ;
        RECT 85.985 124.355 96.995 125.265 ;
        RECT 97.925 124.355 101.595 125.165 ;
        RECT 102.065 124.355 103.435 125.165 ;
        RECT 103.445 124.355 107.115 125.165 ;
        RECT 110.325 125.035 111.255 125.265 ;
        RECT 114.465 125.035 115.395 125.265 ;
        RECT 107.355 124.355 111.255 125.035 ;
        RECT 111.495 124.355 115.395 125.035 ;
        RECT 115.775 125.155 116.695 125.265 ;
        RECT 115.775 125.035 118.110 125.155 ;
        RECT 122.775 125.035 123.695 125.255 ;
        RECT 115.775 124.355 125.055 125.035 ;
        RECT 125.065 124.355 126.435 125.165 ;
        RECT 126.445 124.355 127.815 125.165 ;
        RECT 14.805 124.145 14.975 124.355 ;
        RECT 16.645 124.190 16.805 124.310 ;
        RECT 17.105 124.145 17.275 124.335 ;
        RECT 20.325 124.165 20.495 124.355 ;
        RECT 21.705 124.165 21.875 124.355 ;
        RECT 22.625 124.200 22.785 124.310 ;
        RECT 23.085 124.165 23.255 124.355 ;
        RECT 25.845 124.165 26.015 124.355 ;
        RECT 26.580 124.165 26.750 124.355 ;
        RECT 27.685 124.145 27.855 124.335 ;
        RECT 32.745 124.165 32.915 124.355 ;
        RECT 36.610 124.165 36.780 124.355 ;
        RECT 37.365 124.335 37.515 124.355 ;
        RECT 40.585 124.335 40.735 124.355 ;
        RECT 42.885 124.335 43.035 124.355 ;
        RECT 36.885 124.145 37.055 124.335 ;
        RECT 37.345 124.165 37.515 124.335 ;
        RECT 40.105 124.200 40.265 124.310 ;
        RECT 40.565 124.165 40.735 124.335 ;
        RECT 41.210 124.145 41.380 124.335 ;
        RECT 42.865 124.165 43.035 124.335 ;
        RECT 47.005 124.335 47.155 124.355 ;
        RECT 47.005 124.145 47.175 124.335 ;
        RECT 49.765 124.165 49.935 124.355 ;
        RECT 50.740 124.195 50.860 124.305 ;
        RECT 51.145 124.165 51.315 124.355 ;
        RECT 52.525 124.145 52.695 124.335 ;
        RECT 62.185 124.145 62.355 124.335 ;
        RECT 62.700 124.195 62.820 124.305 ;
        RECT 63.750 124.165 63.920 124.355 ;
        RECT 64.540 124.195 64.660 124.305 ;
        RECT 66.970 124.145 67.140 124.335 ;
        RECT 68.165 124.165 68.335 124.355 ;
        RECT 69.545 124.165 69.715 124.355 ;
        RECT 70.005 124.145 70.175 124.355 ;
        RECT 72.305 124.165 72.475 124.355 ;
        RECT 72.765 124.165 72.935 124.355 ;
        RECT 75.525 124.305 75.695 124.335 ;
        RECT 75.525 124.195 75.700 124.305 ;
        RECT 75.525 124.145 75.695 124.195 ;
        RECT 81.045 124.145 81.215 124.335 ;
        RECT 82.425 124.145 82.595 124.335 ;
        RECT 82.940 124.195 83.060 124.305 ;
        RECT 83.345 124.145 83.515 124.335 ;
        RECT 84.780 124.195 84.900 124.305 ;
        RECT 85.645 124.165 85.815 124.355 ;
        RECT 88.405 124.145 88.575 124.335 ;
        RECT 89.325 124.145 89.495 124.335 ;
        RECT 96.680 124.165 96.850 124.355 ;
        RECT 97.605 124.200 97.765 124.310 ;
        RECT 99.445 124.145 99.615 124.335 ;
        RECT 101.285 124.165 101.455 124.355 ;
        RECT 103.125 124.165 103.295 124.355 ;
        RECT 104.965 124.145 105.135 124.335 ;
        RECT 105.425 124.145 105.595 124.335 ;
        RECT 106.805 124.165 106.975 124.355 ;
        RECT 110.670 124.165 110.840 124.355 ;
        RECT 114.810 124.165 114.980 124.355 ;
        RECT 115.140 124.195 115.260 124.305 ;
        RECT 124.745 124.145 124.915 124.355 ;
        RECT 126.125 124.145 126.295 124.355 ;
        RECT 127.505 124.145 127.675 124.355 ;
        RECT 14.665 123.335 16.035 124.145 ;
        RECT 16.965 123.465 26.070 124.145 ;
        RECT 26.165 123.335 27.995 124.145 ;
        RECT 28.090 123.465 37.195 124.145 ;
        RECT 37.895 123.465 41.795 124.145 ;
        RECT 40.865 123.235 41.795 123.465 ;
        RECT 41.805 123.335 47.315 124.145 ;
        RECT 47.325 123.335 52.835 124.145 ;
        RECT 53.215 123.465 62.495 124.145 ;
        RECT 63.655 123.465 67.555 124.145 ;
        RECT 53.215 123.345 55.550 123.465 ;
        RECT 53.215 123.235 54.135 123.345 ;
        RECT 60.215 123.245 61.135 123.465 ;
        RECT 66.625 123.235 67.555 123.465 ;
        RECT 67.565 123.335 70.315 124.145 ;
        RECT 70.325 123.335 75.835 124.145 ;
        RECT 75.845 123.335 81.355 124.145 ;
        RECT 81.375 123.235 82.725 124.145 ;
        RECT 83.205 123.365 84.575 124.145 ;
        RECT 85.045 123.335 88.715 124.145 ;
        RECT 89.185 123.465 98.290 124.145 ;
        RECT 98.385 123.335 99.755 124.145 ;
        RECT 99.765 123.335 105.275 124.145 ;
        RECT 105.285 123.465 114.390 124.145 ;
        RECT 115.775 123.465 125.055 124.145 ;
        RECT 115.775 123.345 118.110 123.465 ;
        RECT 115.775 123.235 116.695 123.345 ;
        RECT 122.775 123.245 123.695 123.465 ;
        RECT 125.065 123.335 126.435 124.145 ;
        RECT 126.445 123.335 127.815 124.145 ;
        RECT 14.665 118.915 16.035 119.725 ;
        RECT 16.505 118.915 20.175 119.725 ;
        RECT 23.385 119.595 24.315 119.825 ;
        RECT 20.415 118.915 24.315 119.595 ;
        RECT 25.705 118.915 27.075 119.695 ;
        RECT 27.545 118.915 29.375 119.725 ;
        RECT 29.395 118.915 30.745 119.825 ;
        RECT 30.775 118.915 32.125 119.825 ;
        RECT 32.515 119.715 33.435 119.825 ;
        RECT 32.515 119.595 34.850 119.715 ;
        RECT 39.515 119.595 40.435 119.815 ;
        RECT 45.005 119.595 45.935 119.825 ;
        RECT 49.145 119.595 50.075 119.825 ;
        RECT 32.515 118.915 41.795 119.595 ;
        RECT 42.035 118.915 45.935 119.595 ;
        RECT 46.175 118.915 50.075 119.595 ;
        RECT 50.555 118.915 51.905 119.825 ;
        RECT 51.925 118.915 53.295 119.725 ;
        RECT 53.445 118.915 56.055 119.825 ;
        RECT 57.185 118.915 59.275 119.725 ;
        RECT 59.655 119.715 60.575 119.825 ;
        RECT 59.655 119.595 61.990 119.715 ;
        RECT 66.655 119.595 67.575 119.815 ;
        RECT 59.655 118.915 68.935 119.595 ;
        RECT 68.945 118.915 70.315 119.695 ;
        RECT 70.785 118.915 74.455 119.725 ;
        RECT 74.475 118.915 75.825 119.825 ;
        RECT 79.965 119.595 80.895 119.825 ;
        RECT 76.995 118.915 80.895 119.595 ;
        RECT 80.905 118.915 82.275 119.695 ;
        RECT 82.295 118.915 83.645 119.825 ;
        RECT 84.125 118.915 85.495 119.695 ;
        RECT 85.505 118.915 89.175 119.725 ;
        RECT 89.195 118.915 90.545 119.825 ;
        RECT 90.575 118.915 91.925 119.825 ;
        RECT 92.315 119.715 93.235 119.825 ;
        RECT 92.315 119.595 94.650 119.715 ;
        RECT 99.315 119.595 100.235 119.815 ;
        RECT 92.315 118.915 101.595 119.595 ;
        RECT 102.065 118.915 103.435 119.695 ;
        RECT 103.455 118.915 104.805 119.825 ;
        RECT 108.025 119.595 108.955 119.825 ;
        RECT 105.055 118.915 108.955 119.595 ;
        RECT 109.335 119.715 110.255 119.825 ;
        RECT 109.335 119.595 111.670 119.715 ;
        RECT 116.335 119.595 117.255 119.815 ;
        RECT 109.335 118.915 118.615 119.595 ;
        RECT 118.635 118.915 119.985 119.825 ;
        RECT 120.465 118.915 121.835 119.695 ;
        RECT 122.765 118.915 126.435 119.725 ;
        RECT 126.445 118.915 127.815 119.725 ;
        RECT 14.805 118.705 14.975 118.915 ;
        RECT 16.240 118.755 16.360 118.865 ;
        RECT 17.565 118.705 17.735 118.895 ;
        RECT 19.865 118.725 20.035 118.915 ;
        RECT 23.730 118.725 23.900 118.915 ;
        RECT 25.385 118.760 25.545 118.870 ;
        RECT 26.765 118.725 26.935 118.915 ;
        RECT 27.225 118.865 27.395 118.895 ;
        RECT 27.225 118.755 27.400 118.865 ;
        RECT 27.225 118.705 27.395 118.755 ;
        RECT 29.065 118.725 29.235 118.915 ;
        RECT 29.525 118.725 29.695 118.915 ;
        RECT 30.905 118.725 31.075 118.915 ;
        RECT 36.885 118.705 37.055 118.895 ;
        RECT 41.485 118.725 41.655 118.915 ;
        RECT 45.350 118.725 45.520 118.915 ;
        RECT 47.005 118.705 47.175 118.895 ;
        RECT 49.490 118.725 49.660 118.915 ;
        RECT 50.685 118.725 50.855 118.915 ;
        RECT 52.985 118.725 53.155 118.915 ;
        RECT 55.740 118.725 55.910 118.915 ;
        RECT 56.260 118.755 56.380 118.865 ;
        RECT 56.665 118.705 56.835 118.895 ;
        RECT 58.045 118.705 58.215 118.895 ;
        RECT 58.560 118.755 58.680 118.865 ;
        RECT 58.965 118.725 59.135 118.915 ;
        RECT 61.265 118.705 61.435 118.895 ;
        RECT 61.725 118.705 61.895 118.895 ;
        RECT 68.625 118.725 68.795 118.915 ;
        RECT 70.005 118.725 70.175 118.915 ;
        RECT 70.520 118.755 70.640 118.865 ;
        RECT 72.765 118.705 72.935 118.895 ;
        RECT 74.145 118.725 74.315 118.915 ;
        RECT 74.605 118.725 74.775 118.915 ;
        RECT 76.500 118.755 76.620 118.865 ;
        RECT 80.310 118.725 80.480 118.915 ;
        RECT 81.965 118.725 82.135 118.915 ;
        RECT 82.425 118.705 82.595 118.895 ;
        RECT 83.160 118.705 83.330 118.895 ;
        RECT 83.345 118.725 83.515 118.915 ;
        RECT 83.860 118.755 83.980 118.865 ;
        RECT 84.265 118.725 84.435 118.915 ;
        RECT 87.080 118.755 87.200 118.865 ;
        RECT 87.485 118.705 87.655 118.895 ;
        RECT 88.865 118.725 89.035 118.915 ;
        RECT 89.325 118.725 89.495 118.915 ;
        RECT 90.705 118.725 90.875 118.915 ;
        RECT 98.525 118.705 98.695 118.895 ;
        RECT 99.905 118.705 100.075 118.895 ;
        RECT 100.825 118.750 100.985 118.860 ;
        RECT 101.285 118.725 101.455 118.915 ;
        RECT 103.125 118.725 103.295 118.915 ;
        RECT 103.585 118.725 103.755 118.915 ;
        RECT 108.370 118.725 108.540 118.915 ;
        RECT 110.485 118.705 110.655 118.895 ;
        RECT 111.865 118.705 112.035 118.895 ;
        RECT 112.380 118.755 112.500 118.865 ;
        RECT 113.705 118.705 113.875 118.895 ;
        RECT 114.220 118.755 114.340 118.865 ;
        RECT 115.140 118.755 115.260 118.865 ;
        RECT 115.545 118.705 115.715 118.895 ;
        RECT 116.980 118.755 117.100 118.865 ;
        RECT 117.385 118.705 117.555 118.895 ;
        RECT 118.305 118.725 118.475 118.915 ;
        RECT 118.765 118.725 118.935 118.915 ;
        RECT 120.200 118.755 120.320 118.865 ;
        RECT 120.605 118.725 120.775 118.915 ;
        RECT 122.445 118.760 122.605 118.870 ;
        RECT 126.125 118.725 126.295 118.915 ;
        RECT 127.505 118.705 127.675 118.915 ;
        RECT 14.665 117.895 16.035 118.705 ;
        RECT 16.045 117.895 17.875 118.705 ;
        RECT 18.255 118.025 27.535 118.705 ;
        RECT 27.915 118.025 37.195 118.705 ;
        RECT 38.035 118.025 47.315 118.705 ;
        RECT 47.695 118.025 56.975 118.705 ;
        RECT 18.255 117.905 20.590 118.025 ;
        RECT 18.255 117.795 19.175 117.905 ;
        RECT 25.255 117.805 26.175 118.025 ;
        RECT 27.915 117.905 30.250 118.025 ;
        RECT 27.915 117.795 28.835 117.905 ;
        RECT 34.915 117.805 35.835 118.025 ;
        RECT 38.035 117.905 40.370 118.025 ;
        RECT 38.035 117.795 38.955 117.905 ;
        RECT 45.035 117.805 45.955 118.025 ;
        RECT 47.695 117.905 50.030 118.025 ;
        RECT 47.695 117.795 48.615 117.905 ;
        RECT 54.695 117.805 55.615 118.025 ;
        RECT 56.995 117.795 58.345 118.705 ;
        RECT 58.825 117.895 61.575 118.705 ;
        RECT 61.595 117.795 62.945 118.705 ;
        RECT 63.795 118.025 73.075 118.705 ;
        RECT 73.455 118.025 82.735 118.705 ;
        RECT 82.745 118.025 86.645 118.705 ;
        RECT 63.795 117.905 66.130 118.025 ;
        RECT 63.795 117.795 64.715 117.905 ;
        RECT 70.795 117.805 71.715 118.025 ;
        RECT 73.455 117.905 75.790 118.025 ;
        RECT 73.455 117.795 74.375 117.905 ;
        RECT 80.455 117.805 81.375 118.025 ;
        RECT 82.745 117.795 83.675 118.025 ;
        RECT 87.355 117.795 88.705 118.705 ;
        RECT 89.555 118.025 98.835 118.705 ;
        RECT 89.555 117.905 91.890 118.025 ;
        RECT 89.555 117.795 90.475 117.905 ;
        RECT 96.555 117.805 97.475 118.025 ;
        RECT 98.845 117.925 100.215 118.705 ;
        RECT 101.515 118.025 110.795 118.705 ;
        RECT 101.515 117.905 103.850 118.025 ;
        RECT 101.515 117.795 102.435 117.905 ;
        RECT 108.515 117.805 109.435 118.025 ;
        RECT 110.805 117.925 112.175 118.705 ;
        RECT 112.655 117.795 114.005 118.705 ;
        RECT 115.405 117.925 116.775 118.705 ;
        RECT 117.245 118.025 126.350 118.705 ;
        RECT 126.445 117.895 127.815 118.705 ;
        RECT 14.665 113.475 16.035 114.285 ;
        RECT 16.505 113.475 20.175 114.285 ;
        RECT 20.195 113.475 21.545 114.385 ;
        RECT 21.575 113.475 22.925 114.385 ;
        RECT 22.945 113.475 24.315 114.255 ;
        RECT 24.785 113.475 33.890 114.155 ;
        RECT 34.070 113.475 43.175 114.155 ;
        RECT 43.185 113.475 44.555 114.255 ;
        RECT 44.575 113.475 45.925 114.385 ;
        RECT 45.945 113.475 47.775 114.285 ;
        RECT 47.785 113.475 49.155 114.255 ;
        RECT 50.545 113.475 52.375 114.285 ;
        RECT 52.385 113.475 53.755 114.255 ;
        RECT 54.685 113.475 60.195 114.285 ;
        RECT 60.205 113.475 65.715 114.285 ;
        RECT 65.735 113.475 67.085 114.385 ;
        RECT 68.025 113.475 69.395 114.255 ;
        RECT 70.325 113.475 75.835 114.285 ;
        RECT 77.595 114.275 78.515 114.385 ;
        RECT 77.595 114.155 79.930 114.275 ;
        RECT 84.595 114.155 85.515 114.375 ;
        RECT 77.595 113.475 86.875 114.155 ;
        RECT 87.345 113.475 91.015 114.285 ;
        RECT 94.225 114.155 95.155 114.385 ;
        RECT 91.255 113.475 95.155 114.155 ;
        RECT 95.625 113.475 97.455 114.285 ;
        RECT 100.665 114.155 101.595 114.385 ;
        RECT 97.695 113.475 101.595 114.155 ;
        RECT 102.065 113.475 105.735 114.285 ;
        RECT 105.745 113.475 111.255 114.285 ;
        RECT 114.465 114.155 115.395 114.385 ;
        RECT 111.495 113.475 115.395 114.155 ;
        RECT 115.405 113.475 117.235 114.285 ;
        RECT 121.755 114.155 122.685 114.375 ;
        RECT 125.515 114.155 126.435 114.385 ;
        RECT 117.245 113.475 126.435 114.155 ;
        RECT 126.445 113.475 127.815 114.285 ;
        RECT 14.805 113.265 14.975 113.475 ;
        RECT 16.240 113.315 16.360 113.425 ;
        RECT 16.645 113.310 16.805 113.420 ;
        RECT 19.865 113.285 20.035 113.475 ;
        RECT 20.325 113.285 20.495 113.475 ;
        RECT 22.625 113.285 22.795 113.475 ;
        RECT 23.085 113.285 23.255 113.475 ;
        RECT 24.925 113.285 25.095 113.475 ;
        RECT 26.305 113.265 26.475 113.455 ;
        RECT 26.765 113.265 26.935 113.455 ;
        RECT 36.885 113.265 37.055 113.455 ;
        RECT 37.805 113.265 37.975 113.455 ;
        RECT 42.865 113.285 43.035 113.475 ;
        RECT 44.245 113.285 44.415 113.475 ;
        RECT 45.625 113.285 45.795 113.475 ;
        RECT 47.465 113.285 47.635 113.475 ;
        RECT 47.925 113.265 48.095 113.455 ;
        RECT 48.845 113.285 49.015 113.475 ;
        RECT 49.765 113.320 49.925 113.430 ;
        RECT 51.605 113.265 51.775 113.455 ;
        RECT 52.065 113.285 52.235 113.475 ;
        RECT 52.525 113.285 52.695 113.475 ;
        RECT 54.365 113.320 54.525 113.430 ;
        RECT 57.125 113.265 57.295 113.455 ;
        RECT 59.885 113.285 60.055 113.475 ;
        RECT 62.645 113.265 62.815 113.455 ;
        RECT 64.025 113.310 64.185 113.420 ;
        RECT 65.405 113.285 65.575 113.475 ;
        RECT 65.865 113.285 66.035 113.475 ;
        RECT 67.705 113.265 67.875 113.455 ;
        RECT 68.165 113.285 68.335 113.475 ;
        RECT 70.005 113.320 70.165 113.430 ;
        RECT 73.225 113.265 73.395 113.455 ;
        RECT 75.525 113.285 75.695 113.475 ;
        RECT 76.905 113.320 77.065 113.430 ;
        RECT 78.745 113.265 78.915 113.455 ;
        RECT 79.205 113.265 79.375 113.455 ;
        RECT 82.880 113.265 83.050 113.455 ;
        RECT 86.565 113.285 86.735 113.475 ;
        RECT 87.080 113.315 87.200 113.425 ;
        RECT 88.405 113.265 88.575 113.455 ;
        RECT 89.380 113.315 89.500 113.425 ;
        RECT 90.705 113.285 90.875 113.475 ;
        RECT 93.005 113.265 93.175 113.455 ;
        RECT 94.385 113.265 94.555 113.455 ;
        RECT 94.570 113.285 94.740 113.475 ;
        RECT 94.900 113.315 95.020 113.425 ;
        RECT 95.360 113.315 95.480 113.425 ;
        RECT 97.145 113.285 97.315 113.475 ;
        RECT 100.365 113.265 100.535 113.455 ;
        RECT 101.010 113.285 101.180 113.475 ;
        RECT 105.425 113.285 105.595 113.475 ;
        RECT 105.885 113.265 106.055 113.455 ;
        RECT 107.265 113.265 107.435 113.455 ;
        RECT 108.645 113.265 108.815 113.455 ;
        RECT 110.945 113.285 111.115 113.475 ;
        RECT 114.165 113.265 114.335 113.455 ;
        RECT 114.810 113.285 114.980 113.475 ;
        RECT 116.925 113.285 117.095 113.475 ;
        RECT 117.385 113.285 117.555 113.475 ;
        RECT 123.825 113.265 123.995 113.455 ;
        RECT 124.285 113.265 124.455 113.455 ;
        RECT 126.125 113.310 126.285 113.420 ;
        RECT 127.505 113.265 127.675 113.475 ;
        RECT 14.665 112.455 16.035 113.265 ;
        RECT 17.335 112.585 26.615 113.265 ;
        RECT 26.625 112.585 35.815 113.265 ;
        RECT 17.335 112.465 19.670 112.585 ;
        RECT 17.335 112.355 18.255 112.465 ;
        RECT 24.335 112.365 25.255 112.585 ;
        RECT 31.135 112.365 32.065 112.585 ;
        RECT 34.895 112.355 35.815 112.585 ;
        RECT 35.825 112.485 37.195 113.265 ;
        RECT 37.665 112.585 46.770 113.265 ;
        RECT 46.865 112.455 48.235 113.265 ;
        RECT 48.245 112.455 51.915 113.265 ;
        RECT 51.925 112.455 57.435 113.265 ;
        RECT 57.445 112.455 62.955 113.265 ;
        RECT 64.345 112.455 68.015 113.265 ;
        RECT 68.025 112.455 73.535 113.265 ;
        RECT 73.545 112.455 79.055 113.265 ;
        RECT 79.075 112.355 80.425 113.265 ;
        RECT 80.585 112.355 83.195 113.265 ;
        RECT 83.205 112.455 88.715 113.265 ;
        RECT 89.645 112.455 93.315 113.265 ;
        RECT 93.335 112.355 94.685 113.265 ;
        RECT 95.165 112.455 100.675 113.265 ;
        RECT 100.685 112.455 106.195 113.265 ;
        RECT 106.205 112.485 107.575 113.265 ;
        RECT 107.585 112.455 108.955 113.265 ;
        RECT 108.965 112.455 114.475 113.265 ;
        RECT 115.030 112.585 124.135 113.265 ;
        RECT 124.145 112.485 125.515 113.265 ;
        RECT 126.445 112.455 127.815 113.265 ;
        RECT 14.665 108.035 16.035 108.845 ;
        RECT 16.045 108.035 17.415 108.845 ;
        RECT 17.425 108.035 22.935 108.845 ;
        RECT 22.955 108.035 24.305 108.945 ;
        RECT 24.785 108.035 26.155 108.845 ;
        RECT 26.165 108.035 27.535 108.815 ;
        RECT 27.545 108.035 28.915 108.815 ;
        RECT 42.635 108.715 43.565 108.935 ;
        RECT 46.395 108.715 47.315 108.945 ;
        RECT 28.925 108.035 38.030 108.715 ;
        RECT 38.125 108.035 47.315 108.715 ;
        RECT 47.325 108.035 48.695 108.815 ;
        RECT 48.705 108.035 50.075 108.845 ;
        RECT 51.005 108.035 52.375 108.815 ;
        RECT 53.305 108.035 56.975 108.845 ;
        RECT 56.985 108.035 58.355 108.815 ;
        RECT 58.365 108.035 60.195 108.845 ;
        RECT 60.205 108.035 62.815 108.945 ;
        RECT 63.425 108.035 64.795 108.815 ;
        RECT 64.890 108.035 73.995 108.715 ;
        RECT 74.475 108.035 75.825 108.945 ;
        RECT 76.850 108.035 85.955 108.715 ;
        RECT 85.975 108.035 87.325 108.945 ;
        RECT 87.345 108.035 88.715 108.815 ;
        RECT 88.810 108.035 97.915 108.715 ;
        RECT 98.855 108.035 100.205 108.945 ;
        RECT 100.225 108.035 101.595 108.815 ;
        RECT 102.150 108.035 111.255 108.715 ;
        RECT 111.265 108.035 112.635 108.815 ;
        RECT 112.645 108.035 114.015 108.815 ;
        RECT 114.485 108.035 115.855 108.815 ;
        RECT 115.875 108.035 117.225 108.945 ;
        RECT 117.245 108.715 118.165 108.945 ;
        RECT 120.995 108.715 121.925 108.935 ;
        RECT 117.245 108.035 126.435 108.715 ;
        RECT 126.445 108.035 127.815 108.845 ;
        RECT 14.805 107.825 14.975 108.035 ;
        RECT 17.105 107.825 17.275 108.035 ;
        RECT 18.485 107.825 18.655 108.015 ;
        RECT 22.625 107.845 22.795 108.035 ;
        RECT 23.085 107.845 23.255 108.035 ;
        RECT 25.845 107.845 26.015 108.035 ;
        RECT 26.305 107.845 26.475 108.035 ;
        RECT 27.685 107.825 27.855 108.035 ;
        RECT 29.065 107.845 29.235 108.035 ;
        RECT 36.885 107.825 37.055 108.015 ;
        RECT 37.805 107.825 37.975 108.015 ;
        RECT 38.265 107.845 38.435 108.035 ;
        RECT 47.465 107.845 47.635 108.035 ;
        RECT 47.925 107.825 48.095 108.015 ;
        RECT 49.765 107.845 49.935 108.035 ;
        RECT 50.740 107.875 50.860 107.985 ;
        RECT 51.145 107.845 51.315 108.035 ;
        RECT 52.985 107.880 53.145 107.990 ;
        RECT 56.665 107.845 56.835 108.035 ;
        RECT 57.125 107.825 57.295 108.035 ;
        RECT 58.505 107.825 58.675 108.015 ;
        RECT 59.885 107.825 60.055 108.035 ;
        RECT 60.350 108.015 60.520 108.035 ;
        RECT 60.345 107.845 60.520 108.015 ;
        RECT 60.345 107.825 60.515 107.845 ;
        RECT 61.725 107.825 61.895 108.015 ;
        RECT 63.160 107.875 63.280 107.985 ;
        RECT 63.565 107.825 63.735 108.035 ;
        RECT 73.685 107.825 73.855 108.035 ;
        RECT 74.200 107.875 74.320 107.985 ;
        RECT 74.605 107.870 74.765 107.980 ;
        RECT 75.525 107.845 75.695 108.035 ;
        RECT 75.985 107.825 76.155 108.015 ;
        RECT 76.445 107.985 76.615 108.015 ;
        RECT 76.445 107.875 76.620 107.985 ;
        RECT 76.445 107.825 76.615 107.875 ;
        RECT 85.645 107.845 85.815 108.035 ;
        RECT 86.105 107.845 86.275 108.035 ;
        RECT 86.565 107.825 86.735 108.015 ;
        RECT 87.485 107.845 87.655 108.035 ;
        RECT 87.945 107.825 88.115 108.015 ;
        RECT 88.460 107.875 88.580 107.985 ;
        RECT 89.785 107.870 89.945 107.980 ;
        RECT 97.605 107.845 97.775 108.035 ;
        RECT 98.525 107.880 98.685 107.990 ;
        RECT 98.985 107.825 99.155 108.035 ;
        RECT 100.365 107.845 100.535 108.035 ;
        RECT 108.185 107.825 108.355 108.015 ;
        RECT 109.565 107.825 109.735 108.015 ;
        RECT 110.025 107.825 110.195 108.015 ;
        RECT 110.945 107.845 111.115 108.035 ;
        RECT 111.405 107.845 111.575 108.035 ;
        RECT 112.785 107.825 112.955 108.035 ;
        RECT 113.245 107.825 113.415 108.015 ;
        RECT 114.220 107.875 114.340 107.985 ;
        RECT 114.625 107.845 114.795 108.035 ;
        RECT 116.005 107.845 116.175 108.035 ;
        RECT 123.825 107.825 123.995 108.015 ;
        RECT 124.285 107.825 124.455 108.015 ;
        RECT 126.125 107.845 126.295 108.035 ;
        RECT 127.505 107.825 127.675 108.035 ;
        RECT 14.665 107.015 16.035 107.825 ;
        RECT 16.045 107.015 17.415 107.825 ;
        RECT 17.435 106.915 18.785 107.825 ;
        RECT 18.805 107.145 27.995 107.825 ;
        RECT 28.005 107.145 37.195 107.825 ;
        RECT 18.805 106.915 19.725 107.145 ;
        RECT 22.555 106.925 23.485 107.145 ;
        RECT 28.005 106.915 28.925 107.145 ;
        RECT 31.755 106.925 32.685 107.145 ;
        RECT 37.675 106.915 39.025 107.825 ;
        RECT 39.130 107.145 48.235 107.825 ;
        RECT 48.245 107.145 57.435 107.825 ;
        RECT 48.245 106.915 49.165 107.145 ;
        RECT 51.995 106.925 52.925 107.145 ;
        RECT 57.455 106.915 58.805 107.825 ;
        RECT 58.825 107.015 60.195 107.825 ;
        RECT 60.215 106.915 61.565 107.825 ;
        RECT 61.585 107.045 62.955 107.825 ;
        RECT 63.435 106.915 64.785 107.825 ;
        RECT 64.805 107.145 73.995 107.825 ;
        RECT 64.805 106.915 65.725 107.145 ;
        RECT 68.555 106.925 69.485 107.145 ;
        RECT 74.935 106.915 76.285 107.825 ;
        RECT 76.305 107.045 77.675 107.825 ;
        RECT 77.685 107.145 86.875 107.825 ;
        RECT 77.685 106.915 78.605 107.145 ;
        RECT 81.435 106.925 82.365 107.145 ;
        RECT 86.885 107.045 88.255 107.825 ;
        RECT 90.105 107.145 99.295 107.825 ;
        RECT 99.305 107.145 108.495 107.825 ;
        RECT 90.105 106.915 91.025 107.145 ;
        RECT 93.855 106.925 94.785 107.145 ;
        RECT 99.305 106.915 100.225 107.145 ;
        RECT 103.055 106.925 103.985 107.145 ;
        RECT 108.515 106.915 109.865 107.825 ;
        RECT 109.895 106.915 111.245 107.825 ;
        RECT 111.265 107.015 113.095 107.825 ;
        RECT 113.115 106.915 114.465 107.825 ;
        RECT 114.945 107.145 124.135 107.825 ;
        RECT 114.945 106.915 115.865 107.145 ;
        RECT 118.695 106.925 119.625 107.145 ;
        RECT 124.155 106.915 125.505 107.825 ;
        RECT 126.445 107.015 127.815 107.825 ;
        RECT 14.665 102.595 16.035 103.405 ;
        RECT 16.045 102.595 18.795 103.405 ;
        RECT 18.805 102.595 24.315 103.405 ;
        RECT 24.785 102.595 26.155 103.405 ;
        RECT 26.175 102.595 27.525 103.505 ;
        RECT 27.555 102.595 28.905 103.505 ;
        RECT 28.925 102.595 30.295 103.375 ;
        RECT 30.305 102.595 31.675 103.375 ;
        RECT 31.685 103.275 32.605 103.505 ;
        RECT 35.435 103.275 36.365 103.495 ;
        RECT 40.885 103.275 41.805 103.505 ;
        RECT 44.635 103.275 45.565 103.495 ;
        RECT 31.685 102.595 40.875 103.275 ;
        RECT 40.885 102.595 50.075 103.275 ;
        RECT 51.475 102.595 52.825 103.505 ;
        RECT 52.845 102.595 54.215 103.405 ;
        RECT 54.225 103.275 55.145 103.505 ;
        RECT 57.975 103.275 58.905 103.495 ;
        RECT 63.425 103.275 64.345 103.505 ;
        RECT 67.175 103.275 68.105 103.495 ;
        RECT 54.225 102.595 63.415 103.275 ;
        RECT 63.425 102.595 72.615 103.275 ;
        RECT 73.085 102.595 75.835 103.405 ;
        RECT 76.305 103.275 77.225 103.505 ;
        RECT 80.055 103.275 80.985 103.495 ;
        RECT 85.505 103.275 86.425 103.505 ;
        RECT 89.255 103.275 90.185 103.495 ;
        RECT 76.305 102.595 85.495 103.275 ;
        RECT 85.505 102.595 94.695 103.275 ;
        RECT 94.705 102.595 96.075 103.375 ;
        RECT 96.085 102.595 101.595 103.405 ;
        RECT 106.575 103.275 107.505 103.495 ;
        RECT 110.335 103.275 111.255 103.505 ;
        RECT 102.065 102.595 111.255 103.275 ;
        RECT 111.265 103.275 112.185 103.505 ;
        RECT 115.015 103.275 115.945 103.495 ;
        RECT 111.265 102.595 120.455 103.275 ;
        RECT 121.385 102.595 125.055 103.405 ;
        RECT 125.065 102.595 126.435 103.375 ;
        RECT 126.445 102.595 127.815 103.405 ;
        RECT 14.805 102.385 14.975 102.595 ;
        RECT 18.485 102.385 18.655 102.595 ;
        RECT 24.005 102.385 24.175 102.595 ;
        RECT 24.980 102.435 25.100 102.545 ;
        RECT 25.845 102.405 26.015 102.595 ;
        RECT 27.225 102.405 27.395 102.595 ;
        RECT 27.685 102.385 27.855 102.595 ;
        RECT 29.985 102.405 30.155 102.595 ;
        RECT 30.445 102.405 30.615 102.595 ;
        RECT 36.885 102.385 37.055 102.575 ;
        RECT 37.860 102.435 37.980 102.545 ;
        RECT 39.185 102.385 39.355 102.575 ;
        RECT 40.565 102.385 40.735 102.595 ;
        RECT 49.765 102.385 49.935 102.595 ;
        RECT 50.740 102.435 50.860 102.545 ;
        RECT 51.145 102.440 51.305 102.550 ;
        RECT 52.525 102.385 52.695 102.595 ;
        RECT 53.905 102.405 54.075 102.595 ;
        RECT 61.725 102.385 61.895 102.575 ;
        RECT 62.645 102.430 62.805 102.540 ;
        RECT 63.105 102.405 63.275 102.595 ;
        RECT 63.565 102.385 63.735 102.575 ;
        RECT 72.305 102.405 72.475 102.595 ;
        RECT 72.820 102.435 72.940 102.545 ;
        RECT 75.525 102.385 75.695 102.595 ;
        RECT 76.445 102.385 76.615 102.575 ;
        RECT 85.185 102.405 85.355 102.595 ;
        RECT 85.700 102.435 85.820 102.545 ;
        RECT 88.405 102.385 88.575 102.575 ;
        RECT 89.325 102.385 89.495 102.575 ;
        RECT 94.385 102.405 94.555 102.595 ;
        RECT 94.845 102.405 95.015 102.595 ;
        RECT 98.580 102.435 98.700 102.545 ;
        RECT 101.285 102.385 101.455 102.595 ;
        RECT 102.205 102.405 102.375 102.595 ;
        RECT 110.945 102.385 111.115 102.575 ;
        RECT 111.460 102.435 111.580 102.545 ;
        RECT 114.165 102.385 114.335 102.575 ;
        RECT 115.085 102.385 115.255 102.575 ;
        RECT 120.145 102.405 120.315 102.595 ;
        RECT 121.065 102.440 121.225 102.550 ;
        RECT 124.340 102.435 124.460 102.545 ;
        RECT 124.745 102.405 124.915 102.595 ;
        RECT 126.115 102.575 126.285 102.595 ;
        RECT 126.115 102.405 126.295 102.575 ;
        RECT 126.125 102.385 126.295 102.405 ;
        RECT 127.505 102.385 127.675 102.595 ;
        RECT 14.665 101.575 16.035 102.385 ;
        RECT 16.045 101.575 18.795 102.385 ;
        RECT 18.805 101.575 24.315 102.385 ;
        RECT 25.245 101.575 27.995 102.385 ;
        RECT 28.090 101.705 37.195 102.385 ;
        RECT 38.135 101.475 39.485 102.385 ;
        RECT 39.505 101.605 40.875 102.385 ;
        RECT 40.970 101.705 50.075 102.385 ;
        RECT 51.005 101.575 52.835 102.385 ;
        RECT 52.930 101.705 62.035 102.385 ;
        RECT 63.425 101.705 72.530 102.385 ;
        RECT 73.085 101.575 75.835 102.385 ;
        RECT 76.305 101.705 85.410 102.385 ;
        RECT 85.965 101.575 88.715 102.385 ;
        RECT 89.185 101.705 98.290 102.385 ;
        RECT 98.845 101.575 101.595 102.385 ;
        RECT 102.150 101.705 111.255 102.385 ;
        RECT 111.725 101.575 114.475 102.385 ;
        RECT 114.945 101.705 124.050 102.385 ;
        RECT 124.605 101.575 126.435 102.385 ;
        RECT 126.445 101.575 127.815 102.385 ;
      LAYER li1 ;
        RECT 74.985 207.335 75.315 208.315 ;
        RECT 78.255 207.975 78.635 208.145 ;
        RECT 78.255 207.805 78.425 207.975 ;
        RECT 80.015 207.805 80.345 208.315 ;
        RECT 74.565 206.925 74.895 207.175 ;
        RECT 75.065 206.735 75.315 207.335 ;
        RECT 74.985 206.105 75.315 206.735 ;
        RECT 77.765 207.605 78.425 207.805 ;
        RECT 78.595 207.635 80.815 207.805 ;
        RECT 77.765 206.675 77.935 207.605 ;
        RECT 78.595 207.435 78.765 207.635 ;
        RECT 78.105 207.265 78.765 207.435 ;
        RECT 78.935 207.295 80.475 207.465 ;
        RECT 78.105 206.845 78.275 207.265 ;
        RECT 78.935 207.095 79.105 207.295 ;
        RECT 78.505 206.925 79.105 207.095 ;
        RECT 79.275 206.925 79.970 207.125 ;
        RECT 80.230 206.845 80.475 207.295 ;
        RECT 78.595 206.675 79.505 206.755 ;
        RECT 80.645 206.675 80.815 207.635 ;
        RECT 77.765 206.195 78.085 206.675 ;
        RECT 78.255 206.585 79.505 206.675 ;
        RECT 78.255 206.505 78.765 206.585 ;
        RECT 78.255 206.105 78.485 206.505 ;
        RECT 79.175 206.105 79.505 206.585 ;
        RECT 80.350 206.130 80.815 206.675 ;
        RECT 65.785 204.965 66.115 205.595 ;
        RECT 67.625 204.965 67.955 205.595 ;
        RECT 65.785 204.365 66.035 204.965 ;
        RECT 66.205 204.525 66.535 204.775 ;
        RECT 67.205 204.525 67.535 204.775 ;
        RECT 67.705 204.365 67.955 204.965 ;
        RECT 65.785 203.385 66.115 204.365 ;
        RECT 67.625 203.385 67.955 204.365 ;
        RECT 68.570 205.055 68.825 205.585 ;
        RECT 69.545 205.385 70.615 205.555 ;
        RECT 68.570 204.405 68.780 205.055 ;
        RECT 69.545 205.030 69.865 205.385 ;
        RECT 69.540 204.855 69.865 205.030 ;
        RECT 68.950 204.555 69.865 204.855 ;
        RECT 70.035 204.815 70.275 205.215 ;
        RECT 70.445 205.155 70.615 205.385 ;
        RECT 71.145 205.315 72.095 205.595 ;
        RECT 72.315 205.405 72.665 205.575 ;
        RECT 70.445 204.985 70.975 205.155 ;
        RECT 68.950 204.525 69.690 204.555 ;
        RECT 68.570 203.525 68.825 204.405 ;
        RECT 69.520 203.935 69.690 204.525 ;
        RECT 70.035 204.445 70.575 204.815 ;
        RECT 70.755 204.705 70.975 204.985 ;
        RECT 71.145 204.535 71.315 205.315 ;
        RECT 70.910 204.365 71.315 204.535 ;
        RECT 71.485 204.525 71.835 205.145 ;
        RECT 70.910 204.275 71.080 204.365 ;
        RECT 72.005 204.355 72.215 205.145 ;
        RECT 69.860 204.105 71.080 204.275 ;
        RECT 71.540 204.195 72.215 204.355 ;
        RECT 69.520 203.765 70.320 203.935 ;
        RECT 70.150 203.475 70.320 203.765 ;
        RECT 70.910 203.725 71.080 204.105 ;
        RECT 71.250 204.185 72.215 204.195 ;
        RECT 72.405 205.015 72.665 205.405 ;
        RECT 74.080 205.375 74.935 205.545 ;
        RECT 75.140 205.375 75.635 205.545 ;
        RECT 72.405 204.325 72.575 205.015 ;
        RECT 72.745 204.665 72.915 204.845 ;
        RECT 73.085 204.835 73.875 205.085 ;
        RECT 74.080 204.665 74.250 205.375 ;
        RECT 74.420 204.865 74.775 205.085 ;
        RECT 72.745 204.495 74.435 204.665 ;
        RECT 71.250 203.895 71.710 204.185 ;
        RECT 72.405 204.155 73.905 204.325 ;
        RECT 72.405 204.015 72.575 204.155 ;
        RECT 72.015 203.845 72.575 204.015 ;
        RECT 70.910 203.385 71.780 203.725 ;
        RECT 72.015 203.385 72.185 203.845 ;
        RECT 73.020 203.815 74.095 203.985 ;
        RECT 73.020 203.475 73.190 203.815 ;
        RECT 73.925 203.475 74.095 203.815 ;
        RECT 74.265 203.715 74.435 204.495 ;
        RECT 74.605 204.275 74.775 204.865 ;
        RECT 74.945 204.465 75.295 205.085 ;
        RECT 74.605 203.885 75.070 204.275 ;
        RECT 75.465 204.015 75.635 205.375 ;
        RECT 75.805 204.185 76.265 205.235 ;
        RECT 75.240 203.845 75.635 204.015 ;
        RECT 75.240 203.715 75.410 203.845 ;
        RECT 74.265 203.385 74.945 203.715 ;
        RECT 75.160 203.385 75.410 203.715 ;
        RECT 76.000 203.400 76.325 204.185 ;
        RECT 76.495 203.385 76.665 205.505 ;
        RECT 77.335 205.215 77.590 205.505 ;
        RECT 76.840 205.045 77.590 205.215 ;
        RECT 77.770 205.055 78.025 205.585 ;
        RECT 78.745 205.385 79.815 205.555 ;
        RECT 76.840 204.055 77.070 205.045 ;
        RECT 77.240 204.225 77.590 204.875 ;
        RECT 77.770 204.405 77.980 205.055 ;
        RECT 78.745 205.030 79.065 205.385 ;
        RECT 78.740 204.855 79.065 205.030 ;
        RECT 78.150 204.555 79.065 204.855 ;
        RECT 79.235 204.815 79.475 205.215 ;
        RECT 79.645 205.155 79.815 205.385 ;
        RECT 80.345 205.315 81.295 205.595 ;
        RECT 81.515 205.405 81.865 205.575 ;
        RECT 79.645 204.985 80.175 205.155 ;
        RECT 78.150 204.525 78.890 204.555 ;
        RECT 76.840 203.885 77.590 204.055 ;
        RECT 77.335 203.385 77.590 203.885 ;
        RECT 77.770 203.525 78.025 204.405 ;
        RECT 78.720 203.935 78.890 204.525 ;
        RECT 79.235 204.445 79.775 204.815 ;
        RECT 79.955 204.705 80.175 204.985 ;
        RECT 80.345 204.535 80.515 205.315 ;
        RECT 80.110 204.365 80.515 204.535 ;
        RECT 80.685 204.525 81.035 205.145 ;
        RECT 80.110 204.275 80.280 204.365 ;
        RECT 81.205 204.355 81.415 205.145 ;
        RECT 79.060 204.105 80.280 204.275 ;
        RECT 80.740 204.195 81.415 204.355 ;
        RECT 78.720 203.765 79.520 203.935 ;
        RECT 79.350 203.475 79.520 203.765 ;
        RECT 80.110 203.725 80.280 204.105 ;
        RECT 80.450 204.185 81.415 204.195 ;
        RECT 81.605 205.015 81.865 205.405 ;
        RECT 83.280 205.375 84.135 205.545 ;
        RECT 84.340 205.375 84.835 205.545 ;
        RECT 81.605 204.325 81.775 205.015 ;
        RECT 81.945 204.665 82.115 204.845 ;
        RECT 82.285 204.835 83.075 205.085 ;
        RECT 83.280 204.665 83.450 205.375 ;
        RECT 83.620 204.865 83.975 205.085 ;
        RECT 81.945 204.495 83.635 204.665 ;
        RECT 80.450 203.895 80.910 204.185 ;
        RECT 81.605 204.155 83.105 204.325 ;
        RECT 81.605 204.015 81.775 204.155 ;
        RECT 81.215 203.845 81.775 204.015 ;
        RECT 80.110 203.385 80.980 203.725 ;
        RECT 81.215 203.385 81.385 203.845 ;
        RECT 82.220 203.815 83.295 203.985 ;
        RECT 82.220 203.475 82.390 203.815 ;
        RECT 83.125 203.475 83.295 203.815 ;
        RECT 83.465 203.715 83.635 204.495 ;
        RECT 83.805 204.275 83.975 204.865 ;
        RECT 84.145 204.465 84.495 205.085 ;
        RECT 83.805 203.885 84.270 204.275 ;
        RECT 84.665 204.015 84.835 205.375 ;
        RECT 85.005 204.185 85.465 205.235 ;
        RECT 84.440 203.845 84.835 204.015 ;
        RECT 84.440 203.715 84.610 203.845 ;
        RECT 83.465 203.385 84.145 203.715 ;
        RECT 84.360 203.385 84.610 203.715 ;
        RECT 85.200 203.400 85.525 204.185 ;
        RECT 85.695 203.385 85.865 205.505 ;
        RECT 86.535 205.215 86.790 205.505 ;
        RECT 86.040 205.045 86.790 205.215 ;
        RECT 86.040 204.055 86.270 205.045 ;
        RECT 86.440 204.225 86.790 204.875 ;
        RECT 86.040 203.885 86.790 204.055 ;
        RECT 86.535 203.385 86.790 203.885 ;
        RECT 60.290 202.375 60.545 202.875 ;
        RECT 60.290 202.205 61.040 202.375 ;
        RECT 60.290 201.385 60.640 202.035 ;
        RECT 60.810 201.215 61.040 202.205 ;
        RECT 60.290 201.045 61.040 201.215 ;
        RECT 60.290 200.755 60.545 201.045 ;
        RECT 61.215 200.755 61.385 202.875 ;
        RECT 61.555 202.075 61.880 202.860 ;
        RECT 62.470 202.545 62.720 202.875 ;
        RECT 62.935 202.545 63.615 202.875 ;
        RECT 62.470 202.415 62.640 202.545 ;
        RECT 62.245 202.245 62.640 202.415 ;
        RECT 61.615 201.025 62.075 202.075 ;
        RECT 62.245 200.885 62.415 202.245 ;
        RECT 62.810 201.985 63.275 202.375 ;
        RECT 62.585 201.175 62.935 201.795 ;
        RECT 63.105 201.395 63.275 201.985 ;
        RECT 63.445 201.765 63.615 202.545 ;
        RECT 63.785 202.445 63.955 202.785 ;
        RECT 64.690 202.445 64.860 202.785 ;
        RECT 63.785 202.275 64.860 202.445 ;
        RECT 65.695 202.415 65.865 202.875 ;
        RECT 66.100 202.535 66.970 202.875 ;
        RECT 65.305 202.245 65.865 202.415 ;
        RECT 65.305 202.105 65.475 202.245 ;
        RECT 63.975 201.935 65.475 202.105 ;
        RECT 66.170 202.075 66.630 202.365 ;
        RECT 63.445 201.595 65.135 201.765 ;
        RECT 63.105 201.175 63.460 201.395 ;
        RECT 63.630 200.885 63.800 201.595 ;
        RECT 64.005 201.175 64.795 201.425 ;
        RECT 64.965 201.415 65.135 201.595 ;
        RECT 65.305 201.245 65.475 201.935 ;
        RECT 62.245 200.715 62.740 200.885 ;
        RECT 62.945 200.715 63.800 200.885 ;
        RECT 65.215 200.855 65.475 201.245 ;
        RECT 65.665 202.065 66.630 202.075 ;
        RECT 66.800 202.155 66.970 202.535 ;
        RECT 67.560 202.495 67.730 202.785 ;
        RECT 67.560 202.325 68.360 202.495 ;
        RECT 65.665 201.905 66.340 202.065 ;
        RECT 66.800 201.985 68.020 202.155 ;
        RECT 65.665 201.115 65.875 201.905 ;
        RECT 66.800 201.895 66.970 201.985 ;
        RECT 66.045 201.115 66.395 201.735 ;
        RECT 66.565 201.725 66.970 201.895 ;
        RECT 66.565 200.945 66.735 201.725 ;
        RECT 66.905 201.275 67.125 201.555 ;
        RECT 67.305 201.445 67.845 201.815 ;
        RECT 68.190 201.705 68.360 202.325 ;
        RECT 68.915 202.035 69.205 202.875 ;
        RECT 69.755 202.035 70.005 202.875 ;
        RECT 70.865 202.075 71.135 202.845 ;
        RECT 71.840 202.440 72.025 202.845 ;
        RECT 71.840 202.265 72.505 202.440 ;
        RECT 68.915 201.865 70.640 202.035 ;
        RECT 66.905 201.105 67.435 201.275 ;
        RECT 65.215 200.685 65.565 200.855 ;
        RECT 65.785 200.665 66.735 200.945 ;
        RECT 67.265 200.875 67.435 201.105 ;
        RECT 67.605 201.045 67.845 201.445 ;
        RECT 68.015 201.695 68.360 201.705 ;
        RECT 68.015 201.485 70.045 201.695 ;
        RECT 68.015 201.230 68.340 201.485 ;
        RECT 70.230 201.315 70.640 201.865 ;
        RECT 68.015 200.875 68.335 201.230 ;
        RECT 67.265 200.705 68.335 200.875 ;
        RECT 68.875 201.145 70.640 201.315 ;
        RECT 70.865 201.905 71.995 202.075 ;
        RECT 68.875 200.665 69.205 201.145 ;
        RECT 69.715 200.665 70.045 201.145 ;
        RECT 70.865 200.995 71.035 201.905 ;
        RECT 71.205 201.155 71.565 201.735 ;
        RECT 71.745 201.405 71.995 201.905 ;
        RECT 72.165 201.235 72.505 202.265 ;
        RECT 72.795 202.115 72.965 202.875 ;
        RECT 72.795 201.945 73.510 202.115 ;
        RECT 73.680 201.970 73.935 202.875 ;
        RECT 72.705 201.395 73.060 201.765 ;
        RECT 73.340 201.735 73.510 201.945 ;
        RECT 73.340 201.405 73.595 201.735 ;
        RECT 71.820 201.065 72.505 201.235 ;
        RECT 73.340 201.215 73.510 201.405 ;
        RECT 73.765 201.240 73.935 201.970 ;
        RECT 70.865 200.665 71.125 200.995 ;
        RECT 71.820 200.665 72.025 201.065 ;
        RECT 72.795 201.045 73.510 201.215 ;
        RECT 72.795 200.665 72.965 201.045 ;
        RECT 73.680 200.665 73.935 201.240 ;
        RECT 76.385 202.075 76.655 202.845 ;
        RECT 77.360 202.440 77.545 202.845 ;
        RECT 77.360 202.265 78.025 202.440 ;
        RECT 76.385 201.905 77.515 202.075 ;
        RECT 76.385 200.995 76.555 201.905 ;
        RECT 76.725 201.155 77.085 201.735 ;
        RECT 77.265 201.405 77.515 201.905 ;
        RECT 77.685 201.235 78.025 202.265 ;
        RECT 78.315 202.115 78.485 202.875 ;
        RECT 78.315 201.945 78.980 202.115 ;
        RECT 79.165 201.970 79.435 202.875 ;
        RECT 78.810 201.800 78.980 201.945 ;
        RECT 78.245 201.395 78.575 201.765 ;
        RECT 78.810 201.470 79.095 201.800 ;
        RECT 77.340 201.065 78.025 201.235 ;
        RECT 78.810 201.215 78.980 201.470 ;
        RECT 76.385 200.665 76.645 200.995 ;
        RECT 77.340 200.665 77.545 201.065 ;
        RECT 78.315 201.045 78.980 201.215 ;
        RECT 79.265 201.170 79.435 201.970 ;
        RECT 78.315 200.665 78.485 201.045 ;
        RECT 79.175 200.665 79.435 201.170 ;
        RECT 79.610 201.855 79.865 202.735 ;
        RECT 81.190 202.495 81.360 202.785 ;
        RECT 80.560 202.325 81.360 202.495 ;
        RECT 81.950 202.535 82.820 202.875 ;
        RECT 79.610 201.205 79.820 201.855 ;
        RECT 80.560 201.735 80.730 202.325 ;
        RECT 81.950 202.155 82.120 202.535 ;
        RECT 83.055 202.415 83.225 202.875 ;
        RECT 84.060 202.445 84.230 202.785 ;
        RECT 84.965 202.445 85.135 202.785 ;
        RECT 80.900 201.985 82.120 202.155 ;
        RECT 82.290 202.075 82.750 202.365 ;
        RECT 83.055 202.245 83.615 202.415 ;
        RECT 84.060 202.275 85.135 202.445 ;
        RECT 85.305 202.545 85.985 202.875 ;
        RECT 86.200 202.545 86.450 202.875 ;
        RECT 83.445 202.105 83.615 202.245 ;
        RECT 82.290 202.065 83.255 202.075 ;
        RECT 81.950 201.895 82.120 201.985 ;
        RECT 82.580 201.905 83.255 202.065 ;
        RECT 79.990 201.705 80.730 201.735 ;
        RECT 79.990 201.405 80.905 201.705 ;
        RECT 80.580 201.230 80.905 201.405 ;
        RECT 79.610 200.675 79.865 201.205 ;
        RECT 80.585 200.875 80.905 201.230 ;
        RECT 81.075 201.445 81.615 201.815 ;
        RECT 81.950 201.725 82.355 201.895 ;
        RECT 81.075 201.045 81.315 201.445 ;
        RECT 81.795 201.275 82.015 201.555 ;
        RECT 81.485 201.105 82.015 201.275 ;
        RECT 81.485 200.875 81.655 201.105 ;
        RECT 80.585 200.705 81.655 200.875 ;
        RECT 82.185 200.945 82.355 201.725 ;
        RECT 82.525 201.115 82.875 201.735 ;
        RECT 83.045 201.115 83.255 201.905 ;
        RECT 83.445 201.935 84.945 202.105 ;
        RECT 83.445 201.245 83.615 201.935 ;
        RECT 85.305 201.765 85.475 202.545 ;
        RECT 86.280 202.415 86.450 202.545 ;
        RECT 83.785 201.595 85.475 201.765 ;
        RECT 85.645 201.985 86.110 202.375 ;
        RECT 86.280 202.245 86.675 202.415 ;
        RECT 83.785 201.415 83.955 201.595 ;
        RECT 82.185 200.665 83.135 200.945 ;
        RECT 83.445 200.855 83.705 201.245 ;
        RECT 84.125 201.175 84.915 201.425 ;
        RECT 83.355 200.685 83.705 200.855 ;
        RECT 85.120 200.885 85.290 201.595 ;
        RECT 85.645 201.395 85.815 201.985 ;
        RECT 85.460 201.175 85.815 201.395 ;
        RECT 85.985 201.175 86.335 201.795 ;
        RECT 86.505 200.885 86.675 202.245 ;
        RECT 87.040 202.075 87.365 202.860 ;
        RECT 86.845 201.025 87.305 202.075 ;
        RECT 85.120 200.715 85.975 200.885 ;
        RECT 86.180 200.715 86.675 200.885 ;
        RECT 87.535 200.755 87.705 202.875 ;
        RECT 88.375 202.375 88.630 202.875 ;
        RECT 87.880 202.205 88.630 202.375 ;
        RECT 87.880 201.215 88.110 202.205 ;
        RECT 88.280 201.385 88.630 202.035 ;
        RECT 87.880 201.045 88.630 201.215 ;
        RECT 88.375 200.755 88.630 201.045 ;
        RECT 65.805 199.650 66.065 200.155 ;
        RECT 66.755 199.775 66.925 200.155 ;
        RECT 67.190 200.070 67.525 200.115 ;
        RECT 65.805 198.850 65.975 199.650 ;
        RECT 66.260 199.605 66.925 199.775 ;
        RECT 67.185 199.605 67.525 200.070 ;
        RECT 66.260 199.350 66.430 199.605 ;
        RECT 66.145 199.020 66.430 199.350 ;
        RECT 66.665 199.055 66.995 199.425 ;
        RECT 66.260 198.875 66.430 199.020 ;
        RECT 67.185 198.915 67.355 199.605 ;
        RECT 67.525 199.085 67.785 199.415 ;
        RECT 65.805 197.945 66.075 198.850 ;
        RECT 66.260 198.705 66.925 198.875 ;
        RECT 66.755 197.945 66.925 198.705 ;
        RECT 67.185 197.945 67.445 198.915 ;
        RECT 67.615 198.535 67.785 199.085 ;
        RECT 67.955 198.715 68.295 199.745 ;
        RECT 68.485 199.645 68.755 199.990 ;
        RECT 68.485 199.475 68.795 199.645 ;
        RECT 68.485 198.715 68.755 199.475 ;
        RECT 68.980 198.715 69.260 199.990 ;
        RECT 69.460 199.825 69.690 200.155 ;
        RECT 69.460 198.535 69.630 199.825 ;
        RECT 70.435 199.755 70.610 200.155 ;
        RECT 69.980 199.585 70.610 199.755 ;
        RECT 69.980 199.415 70.150 199.585 ;
        RECT 69.800 199.085 70.150 199.415 ;
        RECT 67.615 198.365 69.630 198.535 ;
        RECT 69.980 198.565 70.150 199.085 ;
        RECT 70.330 198.735 70.695 199.415 ;
        RECT 69.980 198.395 70.610 198.565 ;
        RECT 68.170 197.945 68.340 198.365 ;
        RECT 69.460 197.945 69.630 198.365 ;
        RECT 70.435 197.945 70.610 198.395 ;
        RECT 70.865 197.945 71.125 200.155 ;
        RECT 71.835 199.415 72.030 199.990 ;
        RECT 72.300 199.415 72.485 199.995 ;
        RECT 71.295 198.495 71.465 199.415 ;
        RECT 71.775 199.085 72.030 199.415 ;
        RECT 72.255 199.085 72.485 199.415 ;
        RECT 72.735 199.985 74.215 200.155 ;
        RECT 72.735 199.085 72.905 199.985 ;
        RECT 73.075 199.485 73.625 199.815 ;
        RECT 73.815 199.655 74.215 199.985 ;
        RECT 75.035 199.825 75.295 200.155 ;
        RECT 71.835 198.775 72.030 199.085 ;
        RECT 72.300 198.775 72.485 199.085 ;
        RECT 73.075 198.495 73.245 199.485 ;
        RECT 73.815 199.175 73.985 199.655 ;
        RECT 74.565 199.465 74.775 199.645 ;
        RECT 74.155 199.295 74.775 199.465 ;
        RECT 71.295 198.325 73.245 198.495 ;
        RECT 73.415 199.005 73.985 199.175 ;
        RECT 75.125 199.125 75.295 199.825 ;
        RECT 73.415 198.495 73.585 199.005 ;
        RECT 74.165 198.955 75.295 199.125 ;
        RECT 74.165 198.835 74.335 198.955 ;
        RECT 73.755 198.665 74.335 198.835 ;
        RECT 73.415 198.325 74.155 198.495 ;
        RECT 74.605 198.455 74.955 198.785 ;
        RECT 72.050 197.945 72.220 198.325 ;
        RECT 73.005 197.945 73.175 198.325 ;
        RECT 73.965 197.945 74.155 198.325 ;
        RECT 75.125 198.275 75.295 198.955 ;
        RECT 75.035 197.945 75.295 198.275 ;
        RECT 75.465 199.585 75.850 200.155 ;
        RECT 76.865 199.695 77.145 200.155 ;
        RECT 75.465 198.915 75.745 199.585 ;
        RECT 76.020 199.525 77.145 199.695 ;
        RECT 76.020 199.415 76.470 199.525 ;
        RECT 75.915 199.085 76.470 199.415 ;
        RECT 77.335 199.355 77.735 200.155 ;
        RECT 78.575 199.695 78.860 200.155 ;
        RECT 75.465 197.945 75.850 198.915 ;
        RECT 76.020 198.625 76.470 199.085 ;
        RECT 76.640 198.795 77.735 199.355 ;
        RECT 76.020 198.405 77.145 198.625 ;
        RECT 76.865 197.945 77.145 198.405 ;
        RECT 77.335 197.945 77.735 198.795 ;
        RECT 77.905 199.525 78.860 199.695 ;
        RECT 79.145 199.675 79.405 200.155 ;
        RECT 77.905 198.625 78.115 199.525 ;
        RECT 78.285 198.795 78.975 199.355 ;
        RECT 79.145 198.645 79.315 199.675 ;
        RECT 79.995 199.645 80.215 200.105 ;
        RECT 79.965 199.620 80.215 199.645 ;
        RECT 79.485 199.025 79.715 199.420 ;
        RECT 79.885 199.195 80.215 199.620 ;
        RECT 80.385 199.945 81.275 200.115 ;
        RECT 80.385 199.220 80.555 199.945 ;
        RECT 80.725 199.390 81.275 199.775 ;
        RECT 81.445 199.525 82.140 200.155 ;
        RECT 81.965 199.475 82.140 199.525 ;
        RECT 80.385 199.150 81.275 199.220 ;
        RECT 80.380 199.125 81.275 199.150 ;
        RECT 80.370 199.110 81.275 199.125 ;
        RECT 80.365 199.095 81.275 199.110 ;
        RECT 80.355 199.090 81.275 199.095 ;
        RECT 80.350 199.080 81.275 199.090 ;
        RECT 81.465 199.085 81.800 199.335 ;
        RECT 80.345 199.070 81.275 199.080 ;
        RECT 80.335 199.065 81.275 199.070 ;
        RECT 80.325 199.055 81.275 199.065 ;
        RECT 80.315 199.050 81.275 199.055 ;
        RECT 80.315 199.045 80.650 199.050 ;
        RECT 80.300 199.040 80.650 199.045 ;
        RECT 80.285 199.030 80.650 199.040 ;
        RECT 80.260 199.025 80.650 199.030 ;
        RECT 79.485 199.020 80.650 199.025 ;
        RECT 79.485 198.985 80.620 199.020 ;
        RECT 79.485 198.960 80.585 198.985 ;
        RECT 79.485 198.930 80.555 198.960 ;
        RECT 79.485 198.900 80.535 198.930 ;
        RECT 79.485 198.870 80.515 198.900 ;
        RECT 79.485 198.860 80.445 198.870 ;
        RECT 79.485 198.850 80.420 198.860 ;
        RECT 79.485 198.835 80.400 198.850 ;
        RECT 79.485 198.820 80.380 198.835 ;
        RECT 79.590 198.810 80.375 198.820 ;
        RECT 79.590 198.775 80.360 198.810 ;
        RECT 77.905 198.405 78.860 198.625 ;
        RECT 78.575 197.945 78.860 198.405 ;
        RECT 79.145 197.945 79.420 198.645 ;
        RECT 79.590 198.525 80.345 198.775 ;
        RECT 81.015 198.600 81.275 199.050 ;
        RECT 81.970 198.925 82.140 199.475 ;
        RECT 83.265 199.525 83.595 200.155 ;
        RECT 84.645 199.525 84.975 200.155 ;
        RECT 82.310 199.085 82.645 199.355 ;
        RECT 83.265 198.925 83.515 199.525 ;
        RECT 83.685 199.085 84.015 199.335 ;
        RECT 84.225 199.085 84.555 199.335 ;
        RECT 84.725 198.925 84.975 199.525 ;
        RECT 80.015 197.945 80.495 198.285 ;
        RECT 81.875 197.945 82.205 198.925 ;
        RECT 83.265 197.945 83.595 198.925 ;
        RECT 84.645 197.945 84.975 198.925 ;
        RECT 52.905 196.455 53.235 197.435 ;
        RECT 56.125 196.455 56.455 197.435 ;
        RECT 69.485 196.735 69.760 197.435 ;
        RECT 70.355 197.095 70.835 197.435 ;
        RECT 52.905 195.855 53.155 196.455 ;
        RECT 53.325 196.045 53.655 196.295 ;
        RECT 56.125 195.855 56.375 196.455 ;
        RECT 56.545 196.045 56.875 196.295 ;
        RECT 52.905 195.225 53.235 195.855 ;
        RECT 56.125 195.225 56.455 195.855 ;
        RECT 69.485 195.705 69.655 196.735 ;
        RECT 69.930 196.605 70.685 196.855 ;
        RECT 69.930 196.570 70.700 196.605 ;
        RECT 69.930 196.560 70.715 196.570 ;
        RECT 69.825 196.545 70.720 196.560 ;
        RECT 69.825 196.530 70.740 196.545 ;
        RECT 69.825 196.520 70.760 196.530 ;
        RECT 69.825 196.510 70.785 196.520 ;
        RECT 69.825 196.480 70.855 196.510 ;
        RECT 69.825 196.450 70.875 196.480 ;
        RECT 69.825 196.420 70.895 196.450 ;
        RECT 69.825 196.395 70.925 196.420 ;
        RECT 69.825 196.360 70.960 196.395 ;
        RECT 69.825 196.355 70.990 196.360 ;
        RECT 69.825 195.960 70.055 196.355 ;
        RECT 70.600 196.350 70.990 196.355 ;
        RECT 70.625 196.340 70.990 196.350 ;
        RECT 70.640 196.335 70.990 196.340 ;
        RECT 70.655 196.330 70.990 196.335 ;
        RECT 71.355 196.330 71.615 196.780 ;
        RECT 70.655 196.325 71.615 196.330 ;
        RECT 70.665 196.315 71.615 196.325 ;
        RECT 70.675 196.310 71.615 196.315 ;
        RECT 70.685 196.300 71.615 196.310 ;
        RECT 70.690 196.290 71.615 196.300 ;
        RECT 70.695 196.285 71.615 196.290 ;
        RECT 70.705 196.270 71.615 196.285 ;
        RECT 70.710 196.255 71.615 196.270 ;
        RECT 70.720 196.230 71.615 196.255 ;
        RECT 70.225 195.760 70.555 196.185 ;
        RECT 69.485 195.225 69.745 195.705 ;
        RECT 70.335 195.275 70.555 195.760 ;
        RECT 70.725 196.160 71.615 196.230 ;
        RECT 71.795 196.545 72.125 197.395 ;
        RECT 72.735 196.965 72.985 197.385 ;
        RECT 73.775 196.965 74.025 197.385 ;
        RECT 72.735 196.795 74.025 196.965 ;
        RECT 74.205 196.965 74.535 197.395 ;
        RECT 74.205 196.795 74.660 196.965 ;
        RECT 78.865 196.815 79.400 197.435 ;
        RECT 70.725 195.435 70.895 196.160 ;
        RECT 71.065 195.605 71.615 195.990 ;
        RECT 71.795 195.780 71.985 196.545 ;
        RECT 72.725 196.295 72.940 196.625 ;
        RECT 72.155 195.965 72.465 196.295 ;
        RECT 72.635 195.965 72.940 196.295 ;
        RECT 73.115 195.965 73.400 196.625 ;
        RECT 73.595 195.965 73.860 196.625 ;
        RECT 74.075 195.965 74.320 196.625 ;
        RECT 72.295 195.795 72.465 195.965 ;
        RECT 74.490 195.795 74.660 196.795 ;
        RECT 77.490 196.635 77.880 196.810 ;
        RECT 77.490 196.465 78.915 196.635 ;
        RECT 70.725 195.265 71.615 195.435 ;
        RECT 71.795 195.270 72.125 195.780 ;
        RECT 72.295 195.625 74.660 195.795 ;
        RECT 77.365 195.735 77.720 196.295 ;
        RECT 73.675 195.285 74.005 195.625 ;
        RECT 77.890 195.565 78.060 196.465 ;
        RECT 78.230 195.735 78.495 196.295 ;
        RECT 78.745 195.965 78.915 196.465 ;
        RECT 79.085 195.795 79.400 196.815 ;
        RECT 108.105 196.455 108.435 197.435 ;
        RECT 107.685 196.045 108.015 196.295 ;
        RECT 108.185 195.855 108.435 196.455 ;
        RECT 77.890 195.235 78.170 195.565 ;
        RECT 78.785 195.225 79.400 195.795 ;
        RECT 108.105 195.225 108.435 195.855 ;
        RECT 109.050 196.415 109.305 197.295 ;
        RECT 110.630 197.055 110.800 197.345 ;
        RECT 110.000 196.885 110.800 197.055 ;
        RECT 111.390 197.095 112.260 197.435 ;
        RECT 109.050 195.765 109.260 196.415 ;
        RECT 110.000 196.295 110.170 196.885 ;
        RECT 111.390 196.715 111.560 197.095 ;
        RECT 112.495 196.975 112.665 197.435 ;
        RECT 113.500 197.005 113.670 197.345 ;
        RECT 114.405 197.005 114.575 197.345 ;
        RECT 110.340 196.545 111.560 196.715 ;
        RECT 111.730 196.635 112.190 196.925 ;
        RECT 112.495 196.805 113.055 196.975 ;
        RECT 113.500 196.835 114.575 197.005 ;
        RECT 114.745 197.105 115.425 197.435 ;
        RECT 115.640 197.105 115.890 197.435 ;
        RECT 112.885 196.665 113.055 196.805 ;
        RECT 111.730 196.625 112.695 196.635 ;
        RECT 111.390 196.455 111.560 196.545 ;
        RECT 112.020 196.465 112.695 196.625 ;
        RECT 109.430 196.265 110.170 196.295 ;
        RECT 109.430 195.965 110.345 196.265 ;
        RECT 110.020 195.790 110.345 195.965 ;
        RECT 109.050 195.235 109.305 195.765 ;
        RECT 110.025 195.435 110.345 195.790 ;
        RECT 110.515 196.005 111.055 196.375 ;
        RECT 111.390 196.285 111.795 196.455 ;
        RECT 110.515 195.605 110.755 196.005 ;
        RECT 111.235 195.835 111.455 196.115 ;
        RECT 110.925 195.665 111.455 195.835 ;
        RECT 110.925 195.435 111.095 195.665 ;
        RECT 110.025 195.265 111.095 195.435 ;
        RECT 111.625 195.505 111.795 196.285 ;
        RECT 111.965 195.675 112.315 196.295 ;
        RECT 112.485 195.675 112.695 196.465 ;
        RECT 112.885 196.495 114.385 196.665 ;
        RECT 112.885 195.805 113.055 196.495 ;
        RECT 114.745 196.325 114.915 197.105 ;
        RECT 115.720 196.975 115.890 197.105 ;
        RECT 113.225 196.155 114.915 196.325 ;
        RECT 115.085 196.545 115.550 196.935 ;
        RECT 115.720 196.805 116.115 196.975 ;
        RECT 113.225 195.975 113.395 196.155 ;
        RECT 111.625 195.225 112.575 195.505 ;
        RECT 112.885 195.415 113.145 195.805 ;
        RECT 113.565 195.735 114.355 195.985 ;
        RECT 112.795 195.245 113.145 195.415 ;
        RECT 114.560 195.445 114.730 196.155 ;
        RECT 115.085 195.955 115.255 196.545 ;
        RECT 114.900 195.735 115.255 195.955 ;
        RECT 115.425 195.735 115.775 196.355 ;
        RECT 115.945 195.445 116.115 196.805 ;
        RECT 116.480 196.635 116.805 197.420 ;
        RECT 116.285 195.585 116.745 196.635 ;
        RECT 114.560 195.275 115.415 195.445 ;
        RECT 115.620 195.275 116.115 195.445 ;
        RECT 116.975 195.315 117.145 197.435 ;
        RECT 117.815 196.935 118.070 197.435 ;
        RECT 117.320 196.765 118.070 196.935 ;
        RECT 117.320 195.775 117.550 196.765 ;
        RECT 117.720 195.945 118.070 196.595 ;
        RECT 117.320 195.605 118.070 195.775 ;
        RECT 117.815 195.315 118.070 195.605 ;
        RECT 43.730 194.335 43.985 194.625 ;
        RECT 43.730 194.165 44.480 194.335 ;
        RECT 43.730 193.345 44.080 193.995 ;
        RECT 44.250 193.175 44.480 194.165 ;
        RECT 43.730 193.005 44.480 193.175 ;
        RECT 43.730 192.505 43.985 193.005 ;
        RECT 44.655 192.505 44.825 194.625 ;
        RECT 45.685 194.495 46.180 194.665 ;
        RECT 46.385 194.495 47.240 194.665 ;
        RECT 45.055 193.305 45.515 194.355 ;
        RECT 44.995 192.520 45.320 193.305 ;
        RECT 45.685 193.135 45.855 194.495 ;
        RECT 46.025 193.585 46.375 194.205 ;
        RECT 46.545 193.985 46.900 194.205 ;
        RECT 46.545 193.395 46.715 193.985 ;
        RECT 47.070 193.785 47.240 194.495 ;
        RECT 48.655 194.525 49.005 194.695 ;
        RECT 47.445 193.955 48.235 194.205 ;
        RECT 48.655 194.135 48.915 194.525 ;
        RECT 49.225 194.435 50.175 194.715 ;
        RECT 48.405 193.785 48.575 193.965 ;
        RECT 45.685 192.965 46.080 193.135 ;
        RECT 46.250 193.005 46.715 193.395 ;
        RECT 46.885 193.615 48.575 193.785 ;
        RECT 45.910 192.835 46.080 192.965 ;
        RECT 46.885 192.835 47.055 193.615 ;
        RECT 48.745 193.445 48.915 194.135 ;
        RECT 47.415 193.275 48.915 193.445 ;
        RECT 49.105 193.475 49.315 194.265 ;
        RECT 49.485 193.645 49.835 194.265 ;
        RECT 50.005 193.655 50.175 194.435 ;
        RECT 50.705 194.505 51.775 194.675 ;
        RECT 50.705 194.275 50.875 194.505 ;
        RECT 50.345 194.105 50.875 194.275 ;
        RECT 50.345 193.825 50.565 194.105 ;
        RECT 51.045 193.935 51.285 194.335 ;
        RECT 50.005 193.485 50.410 193.655 ;
        RECT 50.745 193.565 51.285 193.935 ;
        RECT 51.455 194.150 51.775 194.505 ;
        RECT 52.495 194.175 52.750 194.705 ;
        RECT 51.455 193.975 51.780 194.150 ;
        RECT 51.455 193.675 52.370 193.975 ;
        RECT 51.630 193.645 52.370 193.675 ;
        RECT 49.105 193.315 49.780 193.475 ;
        RECT 50.240 193.395 50.410 193.485 ;
        RECT 49.105 193.305 50.070 193.315 ;
        RECT 48.745 193.135 48.915 193.275 ;
        RECT 45.910 192.505 46.160 192.835 ;
        RECT 46.375 192.505 47.055 192.835 ;
        RECT 47.225 192.935 48.300 193.105 ;
        RECT 48.745 192.965 49.305 193.135 ;
        RECT 49.610 193.015 50.070 193.305 ;
        RECT 50.240 193.225 51.460 193.395 ;
        RECT 47.225 192.595 47.395 192.935 ;
        RECT 48.130 192.595 48.300 192.935 ;
        RECT 49.135 192.505 49.305 192.965 ;
        RECT 50.240 192.845 50.410 193.225 ;
        RECT 51.630 193.055 51.800 193.645 ;
        RECT 52.540 193.525 52.750 194.175 ;
        RECT 49.540 192.505 50.410 192.845 ;
        RECT 51.000 192.885 51.800 193.055 ;
        RECT 51.000 192.595 51.170 192.885 ;
        RECT 52.495 192.645 52.750 193.525 ;
        RECT 52.930 194.175 53.185 194.705 ;
        RECT 53.905 194.505 54.975 194.675 ;
        RECT 52.930 193.525 53.140 194.175 ;
        RECT 53.905 194.150 54.225 194.505 ;
        RECT 53.900 193.975 54.225 194.150 ;
        RECT 53.310 193.675 54.225 193.975 ;
        RECT 54.395 193.935 54.635 194.335 ;
        RECT 54.805 194.275 54.975 194.505 ;
        RECT 55.505 194.435 56.455 194.715 ;
        RECT 56.675 194.525 57.025 194.695 ;
        RECT 54.805 194.105 55.335 194.275 ;
        RECT 53.310 193.645 54.050 193.675 ;
        RECT 52.930 192.645 53.185 193.525 ;
        RECT 53.880 193.055 54.050 193.645 ;
        RECT 54.395 193.565 54.935 193.935 ;
        RECT 55.115 193.825 55.335 194.105 ;
        RECT 55.505 193.655 55.675 194.435 ;
        RECT 55.270 193.485 55.675 193.655 ;
        RECT 55.845 193.645 56.195 194.265 ;
        RECT 55.270 193.395 55.440 193.485 ;
        RECT 56.365 193.475 56.575 194.265 ;
        RECT 54.220 193.225 55.440 193.395 ;
        RECT 55.900 193.315 56.575 193.475 ;
        RECT 53.880 192.885 54.680 193.055 ;
        RECT 54.510 192.595 54.680 192.885 ;
        RECT 55.270 192.845 55.440 193.225 ;
        RECT 55.610 193.305 56.575 193.315 ;
        RECT 56.765 194.135 57.025 194.525 ;
        RECT 58.440 194.495 59.295 194.665 ;
        RECT 59.500 194.495 59.995 194.665 ;
        RECT 56.765 193.445 56.935 194.135 ;
        RECT 57.105 193.785 57.275 193.965 ;
        RECT 57.445 193.955 58.235 194.205 ;
        RECT 58.440 193.785 58.610 194.495 ;
        RECT 58.780 193.985 59.135 194.205 ;
        RECT 57.105 193.615 58.795 193.785 ;
        RECT 55.610 193.015 56.070 193.305 ;
        RECT 56.765 193.275 58.265 193.445 ;
        RECT 56.765 193.135 56.935 193.275 ;
        RECT 56.375 192.965 56.935 193.135 ;
        RECT 55.270 192.505 56.140 192.845 ;
        RECT 56.375 192.505 56.545 192.965 ;
        RECT 57.380 192.935 58.455 193.105 ;
        RECT 57.380 192.595 57.550 192.935 ;
        RECT 58.285 192.595 58.455 192.935 ;
        RECT 58.625 192.835 58.795 193.615 ;
        RECT 58.965 193.395 59.135 193.985 ;
        RECT 59.305 193.585 59.655 194.205 ;
        RECT 58.965 193.005 59.430 193.395 ;
        RECT 59.825 193.135 59.995 194.495 ;
        RECT 60.165 193.305 60.625 194.355 ;
        RECT 59.600 192.965 59.995 193.135 ;
        RECT 59.600 192.835 59.770 192.965 ;
        RECT 58.625 192.505 59.305 192.835 ;
        RECT 59.520 192.505 59.770 192.835 ;
        RECT 60.360 192.520 60.685 193.305 ;
        RECT 60.855 192.505 61.025 194.625 ;
        RECT 61.695 194.335 61.950 194.625 ;
        RECT 61.200 194.165 61.950 194.335 ;
        RECT 61.200 193.175 61.430 194.165 ;
        RECT 66.245 194.085 66.575 194.715 ;
        RECT 61.600 193.345 61.950 193.995 ;
        RECT 66.245 193.485 66.495 194.085 ;
        RECT 72.675 194.065 73.005 194.485 ;
        RECT 73.185 194.315 73.445 194.715 ;
        RECT 74.115 194.315 74.285 194.665 ;
        RECT 73.185 194.145 74.850 194.315 ;
        RECT 75.020 194.210 75.295 194.555 ;
        RECT 72.755 193.975 73.005 194.065 ;
        RECT 74.680 193.975 74.850 194.145 ;
        RECT 66.665 193.645 66.995 193.895 ;
        RECT 72.250 193.645 72.585 193.895 ;
        RECT 72.755 193.645 73.470 193.975 ;
        RECT 73.685 193.645 74.510 193.975 ;
        RECT 74.680 193.645 74.955 193.975 ;
        RECT 61.200 193.005 61.950 193.175 ;
        RECT 61.695 192.505 61.950 193.005 ;
        RECT 66.245 192.505 66.575 193.485 ;
        RECT 72.755 193.085 72.925 193.645 ;
        RECT 73.185 193.185 73.515 193.475 ;
        RECT 73.685 193.355 73.930 193.645 ;
        RECT 74.680 193.475 74.850 193.645 ;
        RECT 75.125 193.475 75.295 194.210 ;
        RECT 74.190 193.305 74.850 193.475 ;
        RECT 74.190 193.185 74.360 193.305 ;
        RECT 73.185 193.015 74.360 193.185 ;
        RECT 72.745 192.515 74.360 192.845 ;
        RECT 75.020 192.505 75.295 193.475 ;
        RECT 75.465 194.210 75.740 194.555 ;
        RECT 76.475 194.315 76.645 194.665 ;
        RECT 77.315 194.315 77.575 194.715 ;
        RECT 75.465 193.475 75.635 194.210 ;
        RECT 75.910 194.145 77.575 194.315 ;
        RECT 75.910 193.975 76.080 194.145 ;
        RECT 77.755 194.065 78.085 194.485 ;
        RECT 84.940 194.075 85.185 194.680 ;
        RECT 77.755 193.975 78.005 194.065 ;
        RECT 75.805 193.645 76.080 193.975 ;
        RECT 76.250 193.645 77.075 193.975 ;
        RECT 77.290 193.645 78.005 193.975 ;
        RECT 84.665 193.905 85.895 194.075 ;
        RECT 78.175 193.645 78.510 193.895 ;
        RECT 75.910 193.475 76.080 193.645 ;
        RECT 75.465 192.505 75.740 193.475 ;
        RECT 75.910 193.305 76.570 193.475 ;
        RECT 76.830 193.355 77.075 193.645 ;
        RECT 76.400 193.185 76.570 193.305 ;
        RECT 77.245 193.185 77.575 193.475 ;
        RECT 76.400 193.015 77.575 193.185 ;
        RECT 77.835 193.085 78.005 193.645 ;
        RECT 84.665 193.095 85.005 193.905 ;
        RECT 85.175 193.340 85.925 193.530 ;
        RECT 76.400 192.515 78.015 192.845 ;
        RECT 84.665 192.685 85.180 193.095 ;
        RECT 85.755 192.675 85.925 193.340 ;
        RECT 86.095 193.355 86.285 194.715 ;
        RECT 86.455 193.865 86.730 194.715 ;
        RECT 86.920 194.350 87.450 194.715 ;
        RECT 87.275 194.315 87.450 194.350 ;
        RECT 86.455 193.695 86.735 193.865 ;
        RECT 86.455 193.555 86.730 193.695 ;
        RECT 86.935 193.355 87.105 194.155 ;
        RECT 86.095 193.185 87.105 193.355 ;
        RECT 87.275 194.145 88.205 194.315 ;
        RECT 88.375 194.145 88.630 194.715 ;
        RECT 87.275 193.015 87.445 194.145 ;
        RECT 88.035 193.975 88.205 194.145 ;
        RECT 86.320 192.845 87.445 193.015 ;
        RECT 87.615 193.645 87.810 193.975 ;
        RECT 88.035 193.645 88.290 193.975 ;
        RECT 87.615 192.675 87.785 193.645 ;
        RECT 88.460 193.475 88.630 194.145 ;
        RECT 85.755 192.505 87.785 192.675 ;
        RECT 88.295 192.505 88.630 193.475 ;
        RECT 90.165 194.085 90.495 194.715 ;
        RECT 91.655 194.335 91.825 194.715 ;
        RECT 91.655 194.165 92.320 194.335 ;
        RECT 92.515 194.210 92.775 194.715 ;
        RECT 90.165 193.485 90.415 194.085 ;
        RECT 90.585 193.645 90.915 193.895 ;
        RECT 91.585 193.615 91.915 193.985 ;
        RECT 92.150 193.910 92.320 194.165 ;
        RECT 92.150 193.580 92.435 193.910 ;
        RECT 90.165 192.505 90.495 193.485 ;
        RECT 92.150 193.435 92.320 193.580 ;
        RECT 91.655 193.265 92.320 193.435 ;
        RECT 92.605 193.410 92.775 194.210 ;
        RECT 96.605 194.085 96.935 194.715 ;
        RECT 96.185 193.645 96.515 193.895 ;
        RECT 96.685 193.485 96.935 194.085 ;
        RECT 91.655 192.505 91.825 193.265 ;
        RECT 92.505 192.505 92.775 193.410 ;
        RECT 96.605 192.505 96.935 193.485 ;
        RECT 97.550 194.175 97.805 194.705 ;
        RECT 98.525 194.505 99.595 194.675 ;
        RECT 97.550 193.525 97.760 194.175 ;
        RECT 98.525 194.150 98.845 194.505 ;
        RECT 98.520 193.975 98.845 194.150 ;
        RECT 97.930 193.675 98.845 193.975 ;
        RECT 99.015 193.935 99.255 194.335 ;
        RECT 99.425 194.275 99.595 194.505 ;
        RECT 100.125 194.435 101.075 194.715 ;
        RECT 101.295 194.525 101.645 194.695 ;
        RECT 99.425 194.105 99.955 194.275 ;
        RECT 97.930 193.645 98.670 193.675 ;
        RECT 97.550 192.645 97.805 193.525 ;
        RECT 98.500 193.055 98.670 193.645 ;
        RECT 99.015 193.565 99.555 193.935 ;
        RECT 99.735 193.825 99.955 194.105 ;
        RECT 100.125 193.655 100.295 194.435 ;
        RECT 99.890 193.485 100.295 193.655 ;
        RECT 100.465 193.645 100.815 194.265 ;
        RECT 99.890 193.395 100.060 193.485 ;
        RECT 100.985 193.475 101.195 194.265 ;
        RECT 98.840 193.225 100.060 193.395 ;
        RECT 100.520 193.315 101.195 193.475 ;
        RECT 98.500 192.885 99.300 193.055 ;
        RECT 99.130 192.595 99.300 192.885 ;
        RECT 99.890 192.845 100.060 193.225 ;
        RECT 100.230 193.305 101.195 193.315 ;
        RECT 101.385 194.135 101.645 194.525 ;
        RECT 103.060 194.495 103.915 194.665 ;
        RECT 104.120 194.495 104.615 194.665 ;
        RECT 101.385 193.445 101.555 194.135 ;
        RECT 101.725 193.785 101.895 193.965 ;
        RECT 102.065 193.955 102.855 194.205 ;
        RECT 103.060 193.785 103.230 194.495 ;
        RECT 103.400 193.985 103.755 194.205 ;
        RECT 101.725 193.615 103.415 193.785 ;
        RECT 100.230 193.015 100.690 193.305 ;
        RECT 101.385 193.275 102.885 193.445 ;
        RECT 101.385 193.135 101.555 193.275 ;
        RECT 100.995 192.965 101.555 193.135 ;
        RECT 99.890 192.505 100.760 192.845 ;
        RECT 100.995 192.505 101.165 192.965 ;
        RECT 102.000 192.935 103.075 193.105 ;
        RECT 102.000 192.595 102.170 192.935 ;
        RECT 102.905 192.595 103.075 192.935 ;
        RECT 103.245 192.835 103.415 193.615 ;
        RECT 103.585 193.395 103.755 193.985 ;
        RECT 103.925 193.585 104.275 194.205 ;
        RECT 103.585 193.005 104.050 193.395 ;
        RECT 104.445 193.135 104.615 194.495 ;
        RECT 104.785 193.305 105.245 194.355 ;
        RECT 104.220 192.965 104.615 193.135 ;
        RECT 104.220 192.835 104.390 192.965 ;
        RECT 103.245 192.505 103.925 192.835 ;
        RECT 104.140 192.505 104.390 192.835 ;
        RECT 104.980 192.520 105.305 193.305 ;
        RECT 105.475 192.505 105.645 194.625 ;
        RECT 106.315 194.335 106.570 194.625 ;
        RECT 105.820 194.165 106.570 194.335 ;
        RECT 105.820 193.175 106.050 194.165 ;
        RECT 106.745 194.145 107.130 194.715 ;
        RECT 108.145 194.255 108.425 194.715 ;
        RECT 106.220 193.345 106.570 193.995 ;
        RECT 106.745 193.475 107.025 194.145 ;
        RECT 107.300 194.085 108.425 194.255 ;
        RECT 107.300 193.975 107.750 194.085 ;
        RECT 107.195 193.645 107.750 193.975 ;
        RECT 108.615 193.915 109.015 194.715 ;
        RECT 109.855 194.255 110.140 194.715 ;
        RECT 105.820 193.005 106.570 193.175 ;
        RECT 106.315 192.505 106.570 193.005 ;
        RECT 106.745 192.505 107.130 193.475 ;
        RECT 107.300 193.185 107.750 193.645 ;
        RECT 107.920 193.355 109.015 193.915 ;
        RECT 107.300 192.965 108.425 193.185 ;
        RECT 108.145 192.505 108.425 192.965 ;
        RECT 108.615 192.505 109.015 193.355 ;
        RECT 109.185 194.085 110.140 194.255 ;
        RECT 109.185 193.185 109.395 194.085 ;
        RECT 110.700 194.075 110.945 194.680 ;
        RECT 109.565 193.355 110.255 193.915 ;
        RECT 110.425 193.905 111.655 194.075 ;
        RECT 109.185 192.965 110.140 193.185 ;
        RECT 109.855 192.505 110.140 192.965 ;
        RECT 110.425 193.095 110.765 193.905 ;
        RECT 110.935 193.340 111.685 193.530 ;
        RECT 110.425 192.685 110.940 193.095 ;
        RECT 111.515 192.675 111.685 193.340 ;
        RECT 111.855 193.355 112.045 194.715 ;
        RECT 112.215 193.865 112.490 194.715 ;
        RECT 112.680 194.350 113.210 194.715 ;
        RECT 113.035 194.315 113.210 194.350 ;
        RECT 112.215 193.695 112.495 193.865 ;
        RECT 112.215 193.555 112.490 193.695 ;
        RECT 112.695 193.355 112.865 194.155 ;
        RECT 111.855 193.185 112.865 193.355 ;
        RECT 113.035 194.145 113.965 194.315 ;
        RECT 114.135 194.145 114.390 194.715 ;
        RECT 113.035 193.015 113.205 194.145 ;
        RECT 113.795 193.975 113.965 194.145 ;
        RECT 112.080 192.845 113.205 193.015 ;
        RECT 113.375 193.645 113.570 193.975 ;
        RECT 113.795 193.645 114.050 193.975 ;
        RECT 113.375 192.675 113.545 193.645 ;
        RECT 114.220 193.475 114.390 194.145 ;
        RECT 111.515 192.505 113.545 192.675 ;
        RECT 114.055 192.505 114.390 193.475 ;
        RECT 115.465 194.085 115.795 194.715 ;
        RECT 115.465 193.485 115.715 194.085 ;
        RECT 115.885 193.645 116.215 193.895 ;
        RECT 115.465 192.505 115.795 193.485 ;
        RECT 37.750 190.975 38.005 191.855 ;
        RECT 39.330 191.615 39.500 191.905 ;
        RECT 38.700 191.445 39.500 191.615 ;
        RECT 40.090 191.655 40.960 191.995 ;
        RECT 37.750 190.325 37.960 190.975 ;
        RECT 38.700 190.855 38.870 191.445 ;
        RECT 40.090 191.275 40.260 191.655 ;
        RECT 41.195 191.535 41.365 191.995 ;
        RECT 42.200 191.565 42.370 191.905 ;
        RECT 43.105 191.565 43.275 191.905 ;
        RECT 39.040 191.105 40.260 191.275 ;
        RECT 40.430 191.195 40.890 191.485 ;
        RECT 41.195 191.365 41.755 191.535 ;
        RECT 42.200 191.395 43.275 191.565 ;
        RECT 43.445 191.665 44.125 191.995 ;
        RECT 44.340 191.665 44.590 191.995 ;
        RECT 41.585 191.225 41.755 191.365 ;
        RECT 40.430 191.185 41.395 191.195 ;
        RECT 40.090 191.015 40.260 191.105 ;
        RECT 40.720 191.025 41.395 191.185 ;
        RECT 38.130 190.825 38.870 190.855 ;
        RECT 38.130 190.525 39.045 190.825 ;
        RECT 38.720 190.350 39.045 190.525 ;
        RECT 37.750 189.795 38.005 190.325 ;
        RECT 38.725 189.995 39.045 190.350 ;
        RECT 39.215 190.565 39.755 190.935 ;
        RECT 40.090 190.845 40.495 191.015 ;
        RECT 39.215 190.165 39.455 190.565 ;
        RECT 39.935 190.395 40.155 190.675 ;
        RECT 39.625 190.225 40.155 190.395 ;
        RECT 39.625 189.995 39.795 190.225 ;
        RECT 38.725 189.825 39.795 189.995 ;
        RECT 40.325 190.065 40.495 190.845 ;
        RECT 40.665 190.235 41.015 190.855 ;
        RECT 41.185 190.235 41.395 191.025 ;
        RECT 41.585 191.055 43.085 191.225 ;
        RECT 41.585 190.365 41.755 191.055 ;
        RECT 43.445 190.885 43.615 191.665 ;
        RECT 44.420 191.535 44.590 191.665 ;
        RECT 41.925 190.715 43.615 190.885 ;
        RECT 43.785 191.105 44.250 191.495 ;
        RECT 44.420 191.365 44.815 191.535 ;
        RECT 41.925 190.535 42.095 190.715 ;
        RECT 40.325 189.785 41.275 190.065 ;
        RECT 41.585 189.975 41.845 190.365 ;
        RECT 42.265 190.295 43.055 190.545 ;
        RECT 41.495 189.805 41.845 189.975 ;
        RECT 43.260 190.005 43.430 190.715 ;
        RECT 43.785 190.515 43.955 191.105 ;
        RECT 43.600 190.295 43.955 190.515 ;
        RECT 44.125 190.295 44.475 190.915 ;
        RECT 44.645 190.005 44.815 191.365 ;
        RECT 45.180 191.195 45.505 191.980 ;
        RECT 44.985 190.145 45.445 191.195 ;
        RECT 43.260 189.835 44.115 190.005 ;
        RECT 44.320 189.835 44.815 190.005 ;
        RECT 45.675 189.875 45.845 191.995 ;
        RECT 46.515 191.495 46.770 191.995 ;
        RECT 46.020 191.325 46.770 191.495 ;
        RECT 46.020 190.335 46.250 191.325 ;
        RECT 46.420 190.505 46.770 191.155 ;
        RECT 51.545 191.090 51.815 191.995 ;
        RECT 52.495 191.235 52.665 191.995 ;
        RECT 54.015 191.825 56.045 191.995 ;
        RECT 46.020 190.165 46.770 190.335 ;
        RECT 46.515 189.875 46.770 190.165 ;
        RECT 51.545 190.290 51.715 191.090 ;
        RECT 52.000 191.065 52.665 191.235 ;
        RECT 52.925 191.405 53.440 191.815 ;
        RECT 52.000 190.920 52.170 191.065 ;
        RECT 51.885 190.590 52.170 190.920 ;
        RECT 52.000 190.335 52.170 190.590 ;
        RECT 52.405 190.515 52.735 190.885 ;
        RECT 52.925 190.595 53.265 191.405 ;
        RECT 54.015 191.160 54.185 191.825 ;
        RECT 54.580 191.485 55.705 191.655 ;
        RECT 53.435 190.970 54.185 191.160 ;
        RECT 54.355 191.145 55.365 191.315 ;
        RECT 52.925 190.425 54.155 190.595 ;
        RECT 51.545 189.785 51.805 190.290 ;
        RECT 52.000 190.165 52.665 190.335 ;
        RECT 52.495 189.785 52.665 190.165 ;
        RECT 53.200 189.820 53.445 190.425 ;
        RECT 54.355 189.785 54.545 191.145 ;
        RECT 54.715 190.125 54.990 190.945 ;
        RECT 55.195 190.345 55.365 191.145 ;
        RECT 55.535 190.355 55.705 191.485 ;
        RECT 55.875 190.855 56.045 191.825 ;
        RECT 56.555 191.025 56.890 191.995 ;
        RECT 58.075 191.235 58.245 191.995 ;
        RECT 58.075 191.065 58.740 191.235 ;
        RECT 58.925 191.090 59.195 191.995 ;
        RECT 62.130 191.495 62.385 191.995 ;
        RECT 62.130 191.325 62.880 191.495 ;
        RECT 55.875 190.525 56.070 190.855 ;
        RECT 56.295 190.525 56.550 190.855 ;
        RECT 56.295 190.355 56.465 190.525 ;
        RECT 56.720 190.355 56.890 191.025 ;
        RECT 58.570 190.920 58.740 191.065 ;
        RECT 58.005 190.515 58.335 190.885 ;
        RECT 58.570 190.590 58.855 190.920 ;
        RECT 55.535 190.185 56.465 190.355 ;
        RECT 55.535 190.150 55.710 190.185 ;
        RECT 54.715 189.955 54.995 190.125 ;
        RECT 54.715 189.785 54.990 189.955 ;
        RECT 55.180 189.785 55.710 190.150 ;
        RECT 56.635 189.785 56.890 190.355 ;
        RECT 58.570 190.335 58.740 190.590 ;
        RECT 58.075 190.165 58.740 190.335 ;
        RECT 59.025 190.290 59.195 191.090 ;
        RECT 62.130 190.505 62.480 191.155 ;
        RECT 62.650 190.335 62.880 191.325 ;
        RECT 58.075 189.785 58.245 190.165 ;
        RECT 58.935 189.785 59.195 190.290 ;
        RECT 62.130 190.165 62.880 190.335 ;
        RECT 62.130 189.875 62.385 190.165 ;
        RECT 63.055 189.875 63.225 191.995 ;
        RECT 63.395 191.195 63.720 191.980 ;
        RECT 64.310 191.665 64.560 191.995 ;
        RECT 64.775 191.665 65.455 191.995 ;
        RECT 64.310 191.535 64.480 191.665 ;
        RECT 64.085 191.365 64.480 191.535 ;
        RECT 63.455 190.145 63.915 191.195 ;
        RECT 64.085 190.005 64.255 191.365 ;
        RECT 64.650 191.105 65.115 191.495 ;
        RECT 64.425 190.295 64.775 190.915 ;
        RECT 64.945 190.515 65.115 191.105 ;
        RECT 65.285 190.885 65.455 191.665 ;
        RECT 65.625 191.565 65.795 191.905 ;
        RECT 66.530 191.565 66.700 191.905 ;
        RECT 65.625 191.395 66.700 191.565 ;
        RECT 67.535 191.535 67.705 191.995 ;
        RECT 67.940 191.655 68.810 191.995 ;
        RECT 67.145 191.365 67.705 191.535 ;
        RECT 67.145 191.225 67.315 191.365 ;
        RECT 65.815 191.055 67.315 191.225 ;
        RECT 68.010 191.195 68.470 191.485 ;
        RECT 65.285 190.715 66.975 190.885 ;
        RECT 64.945 190.295 65.300 190.515 ;
        RECT 65.470 190.005 65.640 190.715 ;
        RECT 65.845 190.295 66.635 190.545 ;
        RECT 66.805 190.535 66.975 190.715 ;
        RECT 67.145 190.365 67.315 191.055 ;
        RECT 64.085 189.835 64.580 190.005 ;
        RECT 64.785 189.835 65.640 190.005 ;
        RECT 67.055 189.975 67.315 190.365 ;
        RECT 67.505 191.185 68.470 191.195 ;
        RECT 68.640 191.275 68.810 191.655 ;
        RECT 69.400 191.615 69.570 191.905 ;
        RECT 69.400 191.445 70.200 191.615 ;
        RECT 67.505 191.025 68.180 191.185 ;
        RECT 68.640 191.105 69.860 191.275 ;
        RECT 67.505 190.235 67.715 191.025 ;
        RECT 68.640 191.015 68.810 191.105 ;
        RECT 67.885 190.235 68.235 190.855 ;
        RECT 68.405 190.845 68.810 191.015 ;
        RECT 68.405 190.065 68.575 190.845 ;
        RECT 68.745 190.395 68.965 190.675 ;
        RECT 69.145 190.565 69.685 190.935 ;
        RECT 70.030 190.855 70.200 191.445 ;
        RECT 70.895 190.975 71.150 191.855 ;
        RECT 71.815 191.655 72.195 191.825 ;
        RECT 71.815 191.485 71.985 191.655 ;
        RECT 73.575 191.485 73.905 191.995 ;
        RECT 70.030 190.825 70.770 190.855 ;
        RECT 68.745 190.225 69.275 190.395 ;
        RECT 67.055 189.805 67.405 189.975 ;
        RECT 67.625 189.785 68.575 190.065 ;
        RECT 69.105 189.995 69.275 190.225 ;
        RECT 69.445 190.165 69.685 190.565 ;
        RECT 69.855 190.525 70.770 190.825 ;
        RECT 69.855 190.350 70.180 190.525 ;
        RECT 69.855 189.995 70.175 190.350 ;
        RECT 70.940 190.325 71.150 190.975 ;
        RECT 69.105 189.825 70.175 189.995 ;
        RECT 70.895 189.795 71.150 190.325 ;
        RECT 71.325 191.285 71.985 191.485 ;
        RECT 72.155 191.315 74.375 191.485 ;
        RECT 71.325 190.355 71.495 191.285 ;
        RECT 72.155 191.115 72.325 191.315 ;
        RECT 71.665 190.945 72.325 191.115 ;
        RECT 72.495 190.975 74.035 191.145 ;
        RECT 71.665 190.525 71.835 190.945 ;
        RECT 72.495 190.775 72.665 190.975 ;
        RECT 72.065 190.605 72.665 190.775 ;
        RECT 72.835 190.605 73.530 190.805 ;
        RECT 73.790 190.525 74.035 190.975 ;
        RECT 72.155 190.355 73.065 190.435 ;
        RECT 74.205 190.355 74.375 191.315 ;
        RECT 76.885 191.195 77.215 191.995 ;
        RECT 77.755 191.195 78.085 191.995 ;
        RECT 76.385 190.525 76.625 191.195 ;
        RECT 76.805 191.025 78.085 191.195 ;
        RECT 86.420 191.185 86.675 191.855 ;
        RECT 87.320 191.445 87.650 191.955 ;
        RECT 76.805 190.355 76.975 191.025 ;
        RECT 77.145 190.525 77.455 190.855 ;
        RECT 77.625 190.525 78.005 190.855 ;
        RECT 78.205 190.525 78.490 190.855 ;
        RECT 77.250 190.355 77.455 190.525 ;
        RECT 71.325 189.875 71.645 190.355 ;
        RECT 71.815 190.265 73.065 190.355 ;
        RECT 71.815 190.185 72.325 190.265 ;
        RECT 71.815 189.785 72.045 190.185 ;
        RECT 72.735 189.785 73.065 190.265 ;
        RECT 73.910 189.810 74.375 190.355 ;
        RECT 76.385 189.785 77.080 190.355 ;
        RECT 77.250 189.830 77.600 190.355 ;
        RECT 77.790 189.830 78.005 190.525 ;
        RECT 86.420 190.325 86.600 191.185 ;
        RECT 87.320 190.855 87.570 191.445 ;
        RECT 87.920 191.295 88.090 191.905 ;
        RECT 88.820 191.615 89.060 191.905 ;
        RECT 89.860 191.695 90.490 191.945 ;
        RECT 89.860 191.615 90.030 191.695 ;
        RECT 91.460 191.615 91.630 191.905 ;
        RECT 92.430 191.780 93.260 191.950 ;
        RECT 88.820 191.445 90.030 191.615 ;
        RECT 86.770 190.525 87.570 190.855 ;
        RECT 86.420 190.125 86.675 190.325 ;
        RECT 86.335 189.955 86.675 190.125 ;
        RECT 86.420 189.795 86.675 189.955 ;
        RECT 87.320 189.875 87.570 190.525 ;
        RECT 87.770 191.275 88.090 191.295 ;
        RECT 87.770 191.105 89.690 191.275 ;
        RECT 87.770 190.210 87.960 191.105 ;
        RECT 89.860 190.935 90.030 191.445 ;
        RECT 90.200 191.185 90.720 191.495 ;
        RECT 88.130 190.765 90.030 190.935 ;
        RECT 88.130 190.705 88.460 190.765 ;
        RECT 88.610 190.535 88.940 190.595 ;
        RECT 88.280 190.265 88.940 190.535 ;
        RECT 87.770 189.880 88.090 190.210 ;
        RECT 89.130 190.005 89.300 190.765 ;
        RECT 90.200 190.595 90.380 191.005 ;
        RECT 89.470 190.425 89.800 190.545 ;
        RECT 90.550 190.425 90.720 191.185 ;
        RECT 89.470 190.255 90.720 190.425 ;
        RECT 90.890 191.365 92.260 191.615 ;
        RECT 90.890 190.595 91.080 191.365 ;
        RECT 92.010 191.105 92.260 191.365 ;
        RECT 91.250 190.935 91.500 191.095 ;
        RECT 92.430 190.935 92.600 191.780 ;
        RECT 93.495 191.495 93.665 191.995 ;
        RECT 92.770 191.105 93.270 191.485 ;
        RECT 93.495 191.325 94.190 191.495 ;
        RECT 91.250 190.765 92.600 190.935 ;
        RECT 92.180 190.725 92.600 190.765 ;
        RECT 90.890 190.255 91.310 190.595 ;
        RECT 91.600 190.265 92.010 190.595 ;
        RECT 89.130 189.835 89.980 190.005 ;
        RECT 91.060 189.825 91.310 190.255 ;
        RECT 92.180 189.995 92.350 190.725 ;
        RECT 92.520 190.175 92.870 190.545 ;
        RECT 93.050 190.235 93.270 191.105 ;
        RECT 93.440 190.535 93.850 191.155 ;
        RECT 94.020 190.355 94.190 191.325 ;
        RECT 93.495 190.165 94.190 190.355 ;
        RECT 92.180 189.795 93.195 189.995 ;
        RECT 93.495 189.835 93.665 190.165 ;
        RECT 94.380 189.875 94.605 191.995 ;
        RECT 95.275 191.495 95.445 191.995 ;
        RECT 98.635 191.825 100.665 191.995 ;
        RECT 94.780 191.325 95.445 191.495 ;
        RECT 97.545 191.405 98.060 191.815 ;
        RECT 94.780 190.335 95.010 191.325 ;
        RECT 95.180 190.505 95.530 191.155 ;
        RECT 97.545 190.595 97.885 191.405 ;
        RECT 98.635 191.160 98.805 191.825 ;
        RECT 99.200 191.485 100.325 191.655 ;
        RECT 98.055 190.970 98.805 191.160 ;
        RECT 98.975 191.145 99.985 191.315 ;
        RECT 97.545 190.425 98.775 190.595 ;
        RECT 94.780 190.165 95.445 190.335 ;
        RECT 95.275 189.875 95.445 190.165 ;
        RECT 97.820 189.820 98.065 190.425 ;
        RECT 98.975 189.785 99.165 191.145 ;
        RECT 99.335 190.125 99.610 190.945 ;
        RECT 99.815 190.345 99.985 191.145 ;
        RECT 100.155 190.355 100.325 191.485 ;
        RECT 100.495 190.855 100.665 191.825 ;
        RECT 101.175 191.025 101.510 191.995 ;
        RECT 102.695 191.235 102.865 191.995 ;
        RECT 102.695 191.065 103.360 191.235 ;
        RECT 103.545 191.090 103.815 191.995 ;
        RECT 107.375 191.825 109.405 191.995 ;
        RECT 100.495 190.525 100.690 190.855 ;
        RECT 100.915 190.525 101.170 190.855 ;
        RECT 100.915 190.355 101.085 190.525 ;
        RECT 101.340 190.355 101.510 191.025 ;
        RECT 103.190 190.920 103.360 191.065 ;
        RECT 102.625 190.515 102.955 190.885 ;
        RECT 103.190 190.590 103.475 190.920 ;
        RECT 100.155 190.185 101.085 190.355 ;
        RECT 100.155 190.150 100.330 190.185 ;
        RECT 99.335 189.955 99.615 190.125 ;
        RECT 99.335 189.785 99.610 189.955 ;
        RECT 99.800 189.785 100.330 190.150 ;
        RECT 101.255 189.785 101.510 190.355 ;
        RECT 103.190 190.335 103.360 190.590 ;
        RECT 102.695 190.165 103.360 190.335 ;
        RECT 103.645 190.290 103.815 191.090 ;
        RECT 106.285 191.405 106.800 191.815 ;
        RECT 106.285 190.595 106.625 191.405 ;
        RECT 107.375 191.160 107.545 191.825 ;
        RECT 107.940 191.485 109.065 191.655 ;
        RECT 106.795 190.970 107.545 191.160 ;
        RECT 107.715 191.145 108.725 191.315 ;
        RECT 106.285 190.425 107.515 190.595 ;
        RECT 102.695 189.785 102.865 190.165 ;
        RECT 103.555 189.785 103.815 190.290 ;
        RECT 106.560 189.820 106.805 190.425 ;
        RECT 107.715 189.785 107.905 191.145 ;
        RECT 108.075 190.805 108.350 190.945 ;
        RECT 108.075 190.635 108.355 190.805 ;
        RECT 108.075 189.785 108.350 190.635 ;
        RECT 108.555 190.345 108.725 191.145 ;
        RECT 108.895 190.355 109.065 191.485 ;
        RECT 109.235 190.855 109.405 191.825 ;
        RECT 109.915 191.025 110.250 191.995 ;
        RECT 109.235 190.525 109.430 190.855 ;
        RECT 109.655 190.525 109.910 190.855 ;
        RECT 109.655 190.355 109.825 190.525 ;
        RECT 110.080 190.355 110.250 191.025 ;
        RECT 108.895 190.185 109.825 190.355 ;
        RECT 108.895 190.150 109.070 190.185 ;
        RECT 108.540 189.785 109.070 190.150 ;
        RECT 109.995 189.785 110.250 190.355 ;
        RECT 110.430 190.975 110.685 191.855 ;
        RECT 112.010 191.615 112.180 191.905 ;
        RECT 111.380 191.445 112.180 191.615 ;
        RECT 112.770 191.655 113.640 191.995 ;
        RECT 110.430 190.325 110.640 190.975 ;
        RECT 111.380 190.855 111.550 191.445 ;
        RECT 112.770 191.275 112.940 191.655 ;
        RECT 113.875 191.535 114.045 191.995 ;
        RECT 114.880 191.565 115.050 191.905 ;
        RECT 115.785 191.565 115.955 191.905 ;
        RECT 111.720 191.105 112.940 191.275 ;
        RECT 113.110 191.195 113.570 191.485 ;
        RECT 113.875 191.365 114.435 191.535 ;
        RECT 114.880 191.395 115.955 191.565 ;
        RECT 116.125 191.665 116.805 191.995 ;
        RECT 117.020 191.665 117.270 191.995 ;
        RECT 114.265 191.225 114.435 191.365 ;
        RECT 113.110 191.185 114.075 191.195 ;
        RECT 112.770 191.015 112.940 191.105 ;
        RECT 113.400 191.025 114.075 191.185 ;
        RECT 110.810 190.825 111.550 190.855 ;
        RECT 110.810 190.525 111.725 190.825 ;
        RECT 111.400 190.350 111.725 190.525 ;
        RECT 110.430 189.795 110.685 190.325 ;
        RECT 111.405 189.995 111.725 190.350 ;
        RECT 111.895 190.565 112.435 190.935 ;
        RECT 112.770 190.845 113.175 191.015 ;
        RECT 111.895 190.165 112.135 190.565 ;
        RECT 112.615 190.395 112.835 190.675 ;
        RECT 112.305 190.225 112.835 190.395 ;
        RECT 112.305 189.995 112.475 190.225 ;
        RECT 111.405 189.825 112.475 189.995 ;
        RECT 113.005 190.065 113.175 190.845 ;
        RECT 113.345 190.235 113.695 190.855 ;
        RECT 113.865 190.235 114.075 191.025 ;
        RECT 114.265 191.055 115.765 191.225 ;
        RECT 114.265 190.365 114.435 191.055 ;
        RECT 116.125 190.885 116.295 191.665 ;
        RECT 117.100 191.535 117.270 191.665 ;
        RECT 114.605 190.715 116.295 190.885 ;
        RECT 116.465 191.105 116.930 191.495 ;
        RECT 117.100 191.365 117.495 191.535 ;
        RECT 114.605 190.535 114.775 190.715 ;
        RECT 113.005 189.785 113.955 190.065 ;
        RECT 114.265 189.975 114.525 190.365 ;
        RECT 114.945 190.295 115.735 190.545 ;
        RECT 114.175 189.805 114.525 189.975 ;
        RECT 115.940 190.005 116.110 190.715 ;
        RECT 116.465 190.515 116.635 191.105 ;
        RECT 116.280 190.295 116.635 190.515 ;
        RECT 116.805 190.295 117.155 190.915 ;
        RECT 117.325 190.005 117.495 191.365 ;
        RECT 117.860 191.195 118.185 191.980 ;
        RECT 117.665 190.145 118.125 191.195 ;
        RECT 115.940 189.835 116.795 190.005 ;
        RECT 117.000 189.835 117.495 190.005 ;
        RECT 118.355 189.875 118.525 191.995 ;
        RECT 119.195 191.495 119.450 191.995 ;
        RECT 118.700 191.325 119.450 191.495 ;
        RECT 118.700 190.335 118.930 191.325 ;
        RECT 119.100 190.505 119.450 191.155 ;
        RECT 118.700 190.165 119.450 190.335 ;
        RECT 119.195 189.875 119.450 190.165 ;
        RECT 29.445 188.645 29.775 189.275 ;
        RECT 34.965 188.645 35.295 189.275 ;
        RECT 35.995 188.895 36.165 189.275 ;
        RECT 35.995 188.725 36.660 188.895 ;
        RECT 36.855 188.770 37.115 189.275 ;
        RECT 29.445 188.045 29.695 188.645 ;
        RECT 29.865 188.205 30.195 188.455 ;
        RECT 34.545 188.205 34.875 188.455 ;
        RECT 35.045 188.045 35.295 188.645 ;
        RECT 35.925 188.175 36.255 188.545 ;
        RECT 36.490 188.470 36.660 188.725 ;
        RECT 29.445 187.065 29.775 188.045 ;
        RECT 34.965 187.065 35.295 188.045 ;
        RECT 36.490 188.140 36.775 188.470 ;
        RECT 36.490 187.995 36.660 188.140 ;
        RECT 35.995 187.825 36.660 187.995 ;
        RECT 36.945 187.970 37.115 188.770 ;
        RECT 37.835 188.895 38.005 189.185 ;
        RECT 37.835 188.725 38.500 188.895 ;
        RECT 35.995 187.065 36.165 187.825 ;
        RECT 36.845 187.065 37.115 187.970 ;
        RECT 37.750 187.905 38.100 188.555 ;
        RECT 38.270 187.735 38.500 188.725 ;
        RECT 37.835 187.565 38.500 187.735 ;
        RECT 37.835 187.065 38.005 187.565 ;
        RECT 38.675 187.065 38.900 189.185 ;
        RECT 39.615 188.895 39.785 189.225 ;
        RECT 40.085 189.065 41.100 189.265 ;
        RECT 39.090 188.705 39.785 188.895 ;
        RECT 39.090 187.735 39.260 188.705 ;
        RECT 39.430 187.905 39.840 188.525 ;
        RECT 40.010 187.955 40.230 188.825 ;
        RECT 40.410 188.515 40.760 188.885 ;
        RECT 40.930 188.335 41.100 189.065 ;
        RECT 41.970 188.805 42.220 189.235 ;
        RECT 43.300 189.055 44.150 189.225 ;
        RECT 41.270 188.465 41.680 188.795 ;
        RECT 41.970 188.465 42.390 188.805 ;
        RECT 40.680 188.295 41.100 188.335 ;
        RECT 40.680 188.125 42.030 188.295 ;
        RECT 39.090 187.565 39.785 187.735 ;
        RECT 40.010 187.575 40.510 187.955 ;
        RECT 39.615 187.065 39.785 187.565 ;
        RECT 40.680 187.280 40.850 188.125 ;
        RECT 41.780 187.965 42.030 188.125 ;
        RECT 41.020 187.695 41.270 187.955 ;
        RECT 42.200 187.695 42.390 188.465 ;
        RECT 41.020 187.445 42.390 187.695 ;
        RECT 42.560 188.635 43.810 188.805 ;
        RECT 42.560 187.875 42.730 188.635 ;
        RECT 43.480 188.515 43.810 188.635 ;
        RECT 42.900 188.055 43.080 188.465 ;
        RECT 43.980 188.295 44.150 189.055 ;
        RECT 45.190 188.850 45.510 189.180 ;
        RECT 44.340 188.525 45.000 188.795 ;
        RECT 44.340 188.465 44.670 188.525 ;
        RECT 44.820 188.295 45.150 188.355 ;
        RECT 43.250 188.125 45.150 188.295 ;
        RECT 42.560 187.565 43.080 187.875 ;
        RECT 43.250 187.615 43.420 188.125 ;
        RECT 45.320 187.955 45.510 188.850 ;
        RECT 43.590 187.785 45.510 187.955 ;
        RECT 45.190 187.765 45.510 187.785 ;
        RECT 45.710 188.535 45.960 189.185 ;
        RECT 46.605 188.735 46.860 189.265 ;
        RECT 45.710 188.205 46.510 188.535 ;
        RECT 43.250 187.445 44.460 187.615 ;
        RECT 40.020 187.110 40.850 187.280 ;
        RECT 41.650 187.155 41.820 187.445 ;
        RECT 43.250 187.365 43.420 187.445 ;
        RECT 42.790 187.115 43.420 187.365 ;
        RECT 44.220 187.155 44.460 187.445 ;
        RECT 45.190 187.155 45.360 187.765 ;
        RECT 45.710 187.615 45.960 188.205 ;
        RECT 46.680 187.875 46.860 188.735 ;
        RECT 47.680 188.635 47.925 189.240 ;
        RECT 45.630 187.105 45.960 187.615 ;
        RECT 46.605 187.405 46.860 187.875 ;
        RECT 47.405 188.465 48.635 188.635 ;
        RECT 47.405 187.655 47.745 188.465 ;
        RECT 47.915 187.900 48.665 188.090 ;
        RECT 46.605 187.235 46.945 187.405 ;
        RECT 47.405 187.245 47.920 187.655 ;
        RECT 48.495 187.235 48.665 187.900 ;
        RECT 48.835 187.915 49.025 189.275 ;
        RECT 49.195 188.425 49.470 189.275 ;
        RECT 49.660 188.910 50.190 189.275 ;
        RECT 50.015 188.875 50.190 188.910 ;
        RECT 49.195 188.255 49.475 188.425 ;
        RECT 49.195 188.115 49.470 188.255 ;
        RECT 49.675 187.915 49.845 188.715 ;
        RECT 48.835 187.745 49.845 187.915 ;
        RECT 50.015 188.705 50.945 188.875 ;
        RECT 51.115 188.705 51.370 189.275 ;
        RECT 50.015 187.575 50.185 188.705 ;
        RECT 50.775 188.535 50.945 188.705 ;
        RECT 49.060 187.405 50.185 187.575 ;
        RECT 50.355 188.205 50.550 188.535 ;
        RECT 50.775 188.205 51.030 188.535 ;
        RECT 50.355 187.235 50.525 188.205 ;
        RECT 51.200 188.035 51.370 188.705 ;
        RECT 51.660 188.815 51.945 189.275 ;
        RECT 51.660 188.645 52.615 188.815 ;
        RECT 46.605 187.205 46.860 187.235 ;
        RECT 48.495 187.065 50.525 187.235 ;
        RECT 51.035 187.065 51.370 188.035 ;
        RECT 51.545 187.915 52.235 188.475 ;
        RECT 52.405 187.745 52.615 188.645 ;
        RECT 51.660 187.525 52.615 187.745 ;
        RECT 52.785 188.475 53.185 189.275 ;
        RECT 53.375 188.815 53.655 189.275 ;
        RECT 53.375 188.645 54.500 188.815 ;
        RECT 54.670 188.705 55.055 189.275 ;
        RECT 54.050 188.535 54.500 188.645 ;
        RECT 52.785 187.915 53.880 188.475 ;
        RECT 54.050 188.205 54.605 188.535 ;
        RECT 51.660 187.065 51.945 187.525 ;
        RECT 52.785 187.065 53.185 187.915 ;
        RECT 54.050 187.745 54.500 188.205 ;
        RECT 54.775 188.035 55.055 188.705 ;
        RECT 68.680 188.815 68.965 189.275 ;
        RECT 68.680 188.645 69.635 188.815 ;
        RECT 53.375 187.525 54.500 187.745 ;
        RECT 53.375 187.065 53.655 187.525 ;
        RECT 54.670 187.065 55.055 188.035 ;
        RECT 68.565 187.915 69.255 188.475 ;
        RECT 69.425 187.745 69.635 188.645 ;
        RECT 68.680 187.525 69.635 187.745 ;
        RECT 69.805 188.475 70.205 189.275 ;
        RECT 70.395 188.815 70.675 189.275 ;
        RECT 70.395 188.645 71.520 188.815 ;
        RECT 71.690 188.705 72.075 189.275 ;
        RECT 71.070 188.535 71.520 188.645 ;
        RECT 69.805 187.915 70.900 188.475 ;
        RECT 71.070 188.205 71.625 188.535 ;
        RECT 68.680 187.065 68.965 187.525 ;
        RECT 69.805 187.065 70.205 187.915 ;
        RECT 71.070 187.745 71.520 188.205 ;
        RECT 71.795 188.035 72.075 188.705 ;
        RECT 79.520 188.735 79.775 189.265 ;
        RECT 79.520 188.085 79.700 188.735 ;
        RECT 80.420 188.535 80.670 189.185 ;
        RECT 79.870 188.205 80.670 188.535 ;
        RECT 70.395 187.525 71.520 187.745 ;
        RECT 70.395 187.065 70.675 187.525 ;
        RECT 71.690 187.065 72.075 188.035 ;
        RECT 79.435 187.915 79.700 188.085 ;
        RECT 79.520 187.875 79.700 187.915 ;
        RECT 79.520 187.205 79.775 187.875 ;
        RECT 80.420 187.615 80.670 188.205 ;
        RECT 80.870 188.850 81.190 189.180 ;
        RECT 82.230 189.055 83.080 189.225 ;
        RECT 80.870 187.955 81.060 188.850 ;
        RECT 81.380 188.525 82.040 188.795 ;
        RECT 81.710 188.465 82.040 188.525 ;
        RECT 81.230 188.295 81.560 188.355 ;
        RECT 82.230 188.295 82.400 189.055 ;
        RECT 84.160 188.805 84.410 189.235 ;
        RECT 82.570 188.635 83.820 188.805 ;
        RECT 82.570 188.515 82.900 188.635 ;
        RECT 81.230 188.125 83.130 188.295 ;
        RECT 80.870 187.785 82.790 187.955 ;
        RECT 80.870 187.765 81.190 187.785 ;
        RECT 80.420 187.105 80.750 187.615 ;
        RECT 81.020 187.155 81.190 187.765 ;
        RECT 82.960 187.615 83.130 188.125 ;
        RECT 83.300 188.055 83.480 188.465 ;
        RECT 83.650 187.875 83.820 188.635 ;
        RECT 81.920 187.445 83.130 187.615 ;
        RECT 83.300 187.565 83.820 187.875 ;
        RECT 83.990 188.465 84.410 188.805 ;
        RECT 85.280 189.065 86.295 189.265 ;
        RECT 84.700 188.465 85.110 188.795 ;
        RECT 83.990 187.695 84.180 188.465 ;
        RECT 85.280 188.335 85.450 189.065 ;
        RECT 86.595 188.895 86.765 189.225 ;
        RECT 85.620 188.515 85.970 188.885 ;
        RECT 85.280 188.295 85.700 188.335 ;
        RECT 84.350 188.125 85.700 188.295 ;
        RECT 84.350 187.965 84.600 188.125 ;
        RECT 85.110 187.695 85.360 187.955 ;
        RECT 83.990 187.445 85.360 187.695 ;
        RECT 81.920 187.155 82.160 187.445 ;
        RECT 82.960 187.365 83.130 187.445 ;
        RECT 82.960 187.115 83.590 187.365 ;
        RECT 84.560 187.155 84.730 187.445 ;
        RECT 85.530 187.280 85.700 188.125 ;
        RECT 86.150 187.955 86.370 188.825 ;
        RECT 86.595 188.705 87.290 188.895 ;
        RECT 85.870 187.575 86.370 187.955 ;
        RECT 86.540 187.905 86.950 188.525 ;
        RECT 87.120 187.735 87.290 188.705 ;
        RECT 86.595 187.565 87.290 187.735 ;
        RECT 85.530 187.110 86.360 187.280 ;
        RECT 86.595 187.065 86.765 187.565 ;
        RECT 87.480 187.065 87.705 189.185 ;
        RECT 88.375 188.895 88.545 189.185 ;
        RECT 87.880 188.725 88.545 188.895 ;
        RECT 87.880 187.735 88.110 188.725 ;
        RECT 89.705 188.645 90.035 189.275 ;
        RECT 90.645 188.770 90.905 189.275 ;
        RECT 91.595 188.895 91.765 189.275 ;
        RECT 88.280 187.905 88.630 188.555 ;
        RECT 89.705 188.045 89.955 188.645 ;
        RECT 90.125 188.205 90.455 188.455 ;
        RECT 87.880 187.565 88.545 187.735 ;
        RECT 88.375 187.065 88.545 187.565 ;
        RECT 89.705 187.065 90.035 188.045 ;
        RECT 90.645 187.970 90.815 188.770 ;
        RECT 91.100 188.725 91.765 188.895 ;
        RECT 94.900 188.815 95.185 189.275 ;
        RECT 91.100 188.470 91.270 188.725 ;
        RECT 94.900 188.645 95.855 188.815 ;
        RECT 90.985 188.140 91.270 188.470 ;
        RECT 91.505 188.175 91.835 188.545 ;
        RECT 91.100 187.995 91.270 188.140 ;
        RECT 90.645 187.065 90.915 187.970 ;
        RECT 91.100 187.825 91.765 187.995 ;
        RECT 94.785 187.915 95.475 188.475 ;
        RECT 91.595 187.065 91.765 187.825 ;
        RECT 95.645 187.745 95.855 188.645 ;
        RECT 94.900 187.525 95.855 187.745 ;
        RECT 96.025 188.475 96.425 189.275 ;
        RECT 96.615 188.815 96.895 189.275 ;
        RECT 96.615 188.645 97.740 188.815 ;
        RECT 97.910 188.705 98.295 189.275 ;
        RECT 97.290 188.535 97.740 188.645 ;
        RECT 96.025 187.915 97.120 188.475 ;
        RECT 97.290 188.205 97.845 188.535 ;
        RECT 94.900 187.065 95.185 187.525 ;
        RECT 96.025 187.065 96.425 187.915 ;
        RECT 97.290 187.745 97.740 188.205 ;
        RECT 98.015 188.035 98.295 188.705 ;
        RECT 96.615 187.525 97.740 187.745 ;
        RECT 96.615 187.065 96.895 187.525 ;
        RECT 97.910 187.065 98.295 188.035 ;
        RECT 98.470 188.735 98.725 189.265 ;
        RECT 99.445 189.065 100.515 189.235 ;
        RECT 98.470 188.085 98.680 188.735 ;
        RECT 99.445 188.710 99.765 189.065 ;
        RECT 99.440 188.535 99.765 188.710 ;
        RECT 98.850 188.235 99.765 188.535 ;
        RECT 99.935 188.495 100.175 188.895 ;
        RECT 100.345 188.835 100.515 189.065 ;
        RECT 101.045 188.995 101.995 189.275 ;
        RECT 102.215 189.085 102.565 189.255 ;
        RECT 100.345 188.665 100.875 188.835 ;
        RECT 98.850 188.205 99.590 188.235 ;
        RECT 98.470 187.205 98.725 188.085 ;
        RECT 99.420 187.615 99.590 188.205 ;
        RECT 99.935 188.125 100.475 188.495 ;
        RECT 100.655 188.385 100.875 188.665 ;
        RECT 101.045 188.215 101.215 188.995 ;
        RECT 100.810 188.045 101.215 188.215 ;
        RECT 101.385 188.205 101.735 188.825 ;
        RECT 100.810 187.955 100.980 188.045 ;
        RECT 101.905 188.035 102.115 188.825 ;
        RECT 99.760 187.785 100.980 187.955 ;
        RECT 101.440 187.875 102.115 188.035 ;
        RECT 99.420 187.445 100.220 187.615 ;
        RECT 100.050 187.155 100.220 187.445 ;
        RECT 100.810 187.405 100.980 187.785 ;
        RECT 101.150 187.865 102.115 187.875 ;
        RECT 102.305 188.695 102.565 189.085 ;
        RECT 103.980 189.055 104.835 189.225 ;
        RECT 105.040 189.055 105.535 189.225 ;
        RECT 102.305 188.005 102.475 188.695 ;
        RECT 102.645 188.345 102.815 188.525 ;
        RECT 102.985 188.515 103.775 188.765 ;
        RECT 103.980 188.345 104.150 189.055 ;
        RECT 104.320 188.545 104.675 188.765 ;
        RECT 102.645 188.175 104.335 188.345 ;
        RECT 101.150 187.575 101.610 187.865 ;
        RECT 102.305 187.835 103.805 188.005 ;
        RECT 102.305 187.695 102.475 187.835 ;
        RECT 101.915 187.525 102.475 187.695 ;
        RECT 100.810 187.065 101.680 187.405 ;
        RECT 101.915 187.065 102.085 187.525 ;
        RECT 102.920 187.495 103.995 187.665 ;
        RECT 102.920 187.155 103.090 187.495 ;
        RECT 103.825 187.155 103.995 187.495 ;
        RECT 104.165 187.395 104.335 188.175 ;
        RECT 104.505 187.955 104.675 188.545 ;
        RECT 104.845 188.145 105.195 188.765 ;
        RECT 104.505 187.565 104.970 187.955 ;
        RECT 105.365 187.695 105.535 189.055 ;
        RECT 105.705 187.865 106.165 188.915 ;
        RECT 105.140 187.525 105.535 187.695 ;
        RECT 105.140 187.395 105.310 187.525 ;
        RECT 104.165 187.065 104.845 187.395 ;
        RECT 105.060 187.065 105.310 187.395 ;
        RECT 105.900 187.080 106.225 187.865 ;
        RECT 106.395 187.065 106.565 189.185 ;
        RECT 107.235 188.895 107.490 189.185 ;
        RECT 106.740 188.725 107.490 188.895 ;
        RECT 113.275 188.895 113.445 189.275 ;
        RECT 113.275 188.725 113.940 188.895 ;
        RECT 114.135 188.770 114.395 189.275 ;
        RECT 106.740 187.735 106.970 188.725 ;
        RECT 107.140 187.905 107.490 188.555 ;
        RECT 113.205 188.175 113.535 188.545 ;
        RECT 113.770 188.470 113.940 188.725 ;
        RECT 113.770 188.140 114.055 188.470 ;
        RECT 113.770 187.995 113.940 188.140 ;
        RECT 113.275 187.825 113.940 187.995 ;
        RECT 114.225 187.970 114.395 188.770 ;
        RECT 116.035 188.895 116.205 189.275 ;
        RECT 116.035 188.725 116.700 188.895 ;
        RECT 116.895 188.770 117.155 189.275 ;
        RECT 115.965 188.175 116.295 188.545 ;
        RECT 116.530 188.470 116.700 188.725 ;
        RECT 116.530 188.140 116.815 188.470 ;
        RECT 116.530 187.995 116.700 188.140 ;
        RECT 106.740 187.565 107.490 187.735 ;
        RECT 107.235 187.065 107.490 187.565 ;
        RECT 113.275 187.065 113.445 187.825 ;
        RECT 114.125 187.065 114.395 187.970 ;
        RECT 116.035 187.825 116.700 187.995 ;
        RECT 116.985 187.970 117.155 188.770 ;
        RECT 116.035 187.065 116.205 187.825 ;
        RECT 116.885 187.065 117.155 187.970 ;
        RECT 25.790 186.055 26.045 186.555 ;
        RECT 25.790 185.885 26.540 186.055 ;
        RECT 25.790 185.065 26.140 185.715 ;
        RECT 26.310 184.895 26.540 185.885 ;
        RECT 25.790 184.725 26.540 184.895 ;
        RECT 25.790 184.435 26.045 184.725 ;
        RECT 26.715 184.435 26.885 186.555 ;
        RECT 27.055 185.755 27.380 186.540 ;
        RECT 27.970 186.225 28.220 186.555 ;
        RECT 28.435 186.225 29.115 186.555 ;
        RECT 27.970 186.095 28.140 186.225 ;
        RECT 27.745 185.925 28.140 186.095 ;
        RECT 27.115 184.705 27.575 185.755 ;
        RECT 27.745 184.565 27.915 185.925 ;
        RECT 28.310 185.665 28.775 186.055 ;
        RECT 28.085 184.855 28.435 185.475 ;
        RECT 28.605 185.075 28.775 185.665 ;
        RECT 28.945 185.445 29.115 186.225 ;
        RECT 29.285 186.125 29.455 186.465 ;
        RECT 30.190 186.125 30.360 186.465 ;
        RECT 29.285 185.955 30.360 186.125 ;
        RECT 31.195 186.095 31.365 186.555 ;
        RECT 31.600 186.215 32.470 186.555 ;
        RECT 30.805 185.925 31.365 186.095 ;
        RECT 30.805 185.785 30.975 185.925 ;
        RECT 29.475 185.615 30.975 185.785 ;
        RECT 31.670 185.755 32.130 186.045 ;
        RECT 28.945 185.275 30.635 185.445 ;
        RECT 28.605 184.855 28.960 185.075 ;
        RECT 29.130 184.565 29.300 185.275 ;
        RECT 29.505 184.855 30.295 185.105 ;
        RECT 30.465 185.095 30.635 185.275 ;
        RECT 30.805 184.925 30.975 185.615 ;
        RECT 27.745 184.395 28.240 184.565 ;
        RECT 28.445 184.395 29.300 184.565 ;
        RECT 30.715 184.535 30.975 184.925 ;
        RECT 31.165 185.745 32.130 185.755 ;
        RECT 32.300 185.835 32.470 186.215 ;
        RECT 33.060 186.175 33.230 186.465 ;
        RECT 33.060 186.005 33.860 186.175 ;
        RECT 31.165 185.585 31.840 185.745 ;
        RECT 32.300 185.665 33.520 185.835 ;
        RECT 31.165 184.795 31.375 185.585 ;
        RECT 32.300 185.575 32.470 185.665 ;
        RECT 31.545 184.795 31.895 185.415 ;
        RECT 32.065 185.405 32.470 185.575 ;
        RECT 32.065 184.625 32.235 185.405 ;
        RECT 32.405 184.955 32.625 185.235 ;
        RECT 32.805 185.125 33.345 185.495 ;
        RECT 33.690 185.415 33.860 186.005 ;
        RECT 34.555 185.535 34.810 186.415 ;
        RECT 38.185 185.575 38.515 186.555 ;
        RECT 33.690 185.385 34.430 185.415 ;
        RECT 32.405 184.785 32.935 184.955 ;
        RECT 30.715 184.365 31.065 184.535 ;
        RECT 31.285 184.345 32.235 184.625 ;
        RECT 32.765 184.555 32.935 184.785 ;
        RECT 33.105 184.725 33.345 185.125 ;
        RECT 33.515 185.085 34.430 185.385 ;
        RECT 33.515 184.910 33.840 185.085 ;
        RECT 33.515 184.555 33.835 184.910 ;
        RECT 34.600 184.885 34.810 185.535 ;
        RECT 37.765 185.165 38.095 185.415 ;
        RECT 38.265 184.975 38.515 185.575 ;
        RECT 32.765 184.385 33.835 184.555 ;
        RECT 34.555 184.355 34.810 184.885 ;
        RECT 38.185 184.345 38.515 184.975 ;
        RECT 39.130 185.585 39.465 186.555 ;
        RECT 39.975 186.385 42.005 186.555 ;
        RECT 39.130 184.915 39.300 185.585 ;
        RECT 39.975 185.415 40.145 186.385 ;
        RECT 39.470 185.085 39.725 185.415 ;
        RECT 39.950 185.085 40.145 185.415 ;
        RECT 40.315 186.045 41.440 186.215 ;
        RECT 39.555 184.915 39.725 185.085 ;
        RECT 40.315 184.915 40.485 186.045 ;
        RECT 39.130 184.345 39.385 184.915 ;
        RECT 39.555 184.745 40.485 184.915 ;
        RECT 40.655 185.705 41.665 185.875 ;
        RECT 40.655 184.905 40.825 185.705 ;
        RECT 40.310 184.710 40.485 184.745 ;
        RECT 40.310 184.345 40.840 184.710 ;
        RECT 41.030 184.685 41.305 185.505 ;
        RECT 41.025 184.515 41.305 184.685 ;
        RECT 41.030 184.345 41.305 184.515 ;
        RECT 41.475 184.345 41.665 185.705 ;
        RECT 41.835 185.720 42.005 186.385 ;
        RECT 42.580 185.965 43.095 186.375 ;
        RECT 41.835 185.530 42.585 185.720 ;
        RECT 42.755 185.155 43.095 185.965 ;
        RECT 41.865 184.985 43.095 185.155 ;
        RECT 44.190 185.585 44.525 186.555 ;
        RECT 45.035 186.385 47.065 186.555 ;
        RECT 42.575 184.380 42.820 184.985 ;
        RECT 44.190 184.915 44.360 185.585 ;
        RECT 45.035 185.415 45.205 186.385 ;
        RECT 44.530 185.085 44.785 185.415 ;
        RECT 45.010 185.085 45.205 185.415 ;
        RECT 45.375 186.045 46.500 186.215 ;
        RECT 44.615 184.915 44.785 185.085 ;
        RECT 45.375 184.915 45.545 186.045 ;
        RECT 44.190 184.345 44.445 184.915 ;
        RECT 44.615 184.745 45.545 184.915 ;
        RECT 45.715 185.705 46.725 185.875 ;
        RECT 45.715 184.905 45.885 185.705 ;
        RECT 45.370 184.710 45.545 184.745 ;
        RECT 45.370 184.345 45.900 184.710 ;
        RECT 46.090 184.685 46.365 185.505 ;
        RECT 46.085 184.515 46.365 184.685 ;
        RECT 46.090 184.345 46.365 184.515 ;
        RECT 46.535 184.345 46.725 185.705 ;
        RECT 46.895 185.720 47.065 186.385 ;
        RECT 47.640 185.965 48.155 186.375 ;
        RECT 46.895 185.530 47.645 185.720 ;
        RECT 47.815 185.155 48.155 185.965 ;
        RECT 46.925 184.985 48.155 185.155 ;
        RECT 49.225 185.575 49.555 186.555 ;
        RECT 47.635 184.380 47.880 184.985 ;
        RECT 49.225 184.975 49.475 185.575 ;
        RECT 50.630 185.535 50.885 186.415 ;
        RECT 52.210 186.175 52.380 186.465 ;
        RECT 51.580 186.005 52.380 186.175 ;
        RECT 52.970 186.215 53.840 186.555 ;
        RECT 49.645 185.165 49.975 185.415 ;
        RECT 49.225 184.345 49.555 184.975 ;
        RECT 50.630 184.885 50.840 185.535 ;
        RECT 51.580 185.415 51.750 186.005 ;
        RECT 52.970 185.835 53.140 186.215 ;
        RECT 54.075 186.095 54.245 186.555 ;
        RECT 55.080 186.125 55.250 186.465 ;
        RECT 55.985 186.125 56.155 186.465 ;
        RECT 51.920 185.665 53.140 185.835 ;
        RECT 53.310 185.755 53.770 186.045 ;
        RECT 54.075 185.925 54.635 186.095 ;
        RECT 55.080 185.955 56.155 186.125 ;
        RECT 56.325 186.225 57.005 186.555 ;
        RECT 57.220 186.225 57.470 186.555 ;
        RECT 54.465 185.785 54.635 185.925 ;
        RECT 53.310 185.745 54.275 185.755 ;
        RECT 52.970 185.575 53.140 185.665 ;
        RECT 53.600 185.585 54.275 185.745 ;
        RECT 51.010 185.385 51.750 185.415 ;
        RECT 51.010 185.085 51.925 185.385 ;
        RECT 51.600 184.910 51.925 185.085 ;
        RECT 50.630 184.355 50.885 184.885 ;
        RECT 51.605 184.555 51.925 184.910 ;
        RECT 52.095 185.125 52.635 185.495 ;
        RECT 52.970 185.405 53.375 185.575 ;
        RECT 52.095 184.725 52.335 185.125 ;
        RECT 52.815 184.955 53.035 185.235 ;
        RECT 52.505 184.785 53.035 184.955 ;
        RECT 52.505 184.555 52.675 184.785 ;
        RECT 51.605 184.385 52.675 184.555 ;
        RECT 53.205 184.625 53.375 185.405 ;
        RECT 53.545 184.795 53.895 185.415 ;
        RECT 54.065 184.795 54.275 185.585 ;
        RECT 54.465 185.615 55.965 185.785 ;
        RECT 54.465 184.925 54.635 185.615 ;
        RECT 56.325 185.445 56.495 186.225 ;
        RECT 57.300 186.095 57.470 186.225 ;
        RECT 54.805 185.275 56.495 185.445 ;
        RECT 56.665 185.665 57.130 186.055 ;
        RECT 57.300 185.925 57.695 186.095 ;
        RECT 54.805 185.095 54.975 185.275 ;
        RECT 53.205 184.345 54.155 184.625 ;
        RECT 54.465 184.535 54.725 184.925 ;
        RECT 55.145 184.855 55.935 185.105 ;
        RECT 54.375 184.365 54.725 184.535 ;
        RECT 56.140 184.565 56.310 185.275 ;
        RECT 56.665 185.075 56.835 185.665 ;
        RECT 56.480 184.855 56.835 185.075 ;
        RECT 57.005 184.855 57.355 185.475 ;
        RECT 57.525 184.565 57.695 185.925 ;
        RECT 58.060 185.755 58.385 186.540 ;
        RECT 57.865 184.705 58.325 185.755 ;
        RECT 56.140 184.395 56.995 184.565 ;
        RECT 57.200 184.395 57.695 184.565 ;
        RECT 58.555 184.435 58.725 186.555 ;
        RECT 59.395 186.055 59.650 186.555 ;
        RECT 58.900 185.885 59.650 186.055 ;
        RECT 79.720 186.095 80.005 186.555 ;
        RECT 58.900 184.895 59.130 185.885 ;
        RECT 79.720 185.875 80.675 186.095 ;
        RECT 59.300 185.065 59.650 185.715 ;
        RECT 79.605 185.145 80.295 185.705 ;
        RECT 80.465 184.975 80.675 185.875 ;
        RECT 58.900 184.725 59.650 184.895 ;
        RECT 59.395 184.435 59.650 184.725 ;
        RECT 79.720 184.805 80.675 184.975 ;
        RECT 80.845 185.705 81.245 186.555 ;
        RECT 81.435 186.095 81.715 186.555 ;
        RECT 81.435 185.875 82.560 186.095 ;
        RECT 80.845 185.145 81.940 185.705 ;
        RECT 82.110 185.415 82.560 185.875 ;
        RECT 82.730 185.585 83.115 186.555 ;
        RECT 86.215 186.385 88.245 186.555 ;
        RECT 79.720 184.345 80.005 184.805 ;
        RECT 80.845 184.345 81.245 185.145 ;
        RECT 82.110 185.085 82.665 185.415 ;
        RECT 82.110 184.975 82.560 185.085 ;
        RECT 81.435 184.805 82.560 184.975 ;
        RECT 82.835 184.915 83.115 185.585 ;
        RECT 85.125 185.965 85.640 186.375 ;
        RECT 85.125 185.155 85.465 185.965 ;
        RECT 86.215 185.720 86.385 186.385 ;
        RECT 86.780 186.045 87.905 186.215 ;
        RECT 85.635 185.530 86.385 185.720 ;
        RECT 86.555 185.705 87.565 185.875 ;
        RECT 85.125 184.985 86.355 185.155 ;
        RECT 81.435 184.345 81.715 184.805 ;
        RECT 82.730 184.345 83.115 184.915 ;
        RECT 85.400 184.380 85.645 184.985 ;
        RECT 86.555 184.345 86.745 185.705 ;
        RECT 86.915 185.025 87.190 185.505 ;
        RECT 86.915 184.855 87.195 185.025 ;
        RECT 87.395 184.905 87.565 185.705 ;
        RECT 87.735 184.915 87.905 186.045 ;
        RECT 88.075 185.415 88.245 186.385 ;
        RECT 88.755 185.585 89.090 186.555 ;
        RECT 88.075 185.085 88.270 185.415 ;
        RECT 88.495 185.085 88.750 185.415 ;
        RECT 88.495 184.915 88.665 185.085 ;
        RECT 88.920 184.915 89.090 185.585 ;
        RECT 86.915 184.345 87.190 184.855 ;
        RECT 87.735 184.745 88.665 184.915 ;
        RECT 87.735 184.710 87.910 184.745 ;
        RECT 87.380 184.345 87.910 184.710 ;
        RECT 88.835 184.345 89.090 184.915 ;
        RECT 89.705 185.575 90.035 186.555 ;
        RECT 92.600 186.095 92.885 186.555 ;
        RECT 92.600 185.875 93.555 186.095 ;
        RECT 89.705 184.975 89.955 185.575 ;
        RECT 90.125 185.165 90.455 185.415 ;
        RECT 92.485 185.145 93.175 185.705 ;
        RECT 93.345 184.975 93.555 185.875 ;
        RECT 89.705 184.345 90.035 184.975 ;
        RECT 92.600 184.805 93.555 184.975 ;
        RECT 93.725 185.705 94.125 186.555 ;
        RECT 94.315 186.095 94.595 186.555 ;
        RECT 94.315 185.875 95.440 186.095 ;
        RECT 93.725 185.145 94.820 185.705 ;
        RECT 94.990 185.415 95.440 185.875 ;
        RECT 95.610 185.585 95.995 186.555 ;
        RECT 97.255 186.385 99.285 186.555 ;
        RECT 92.600 184.345 92.885 184.805 ;
        RECT 93.725 184.345 94.125 185.145 ;
        RECT 94.990 185.085 95.545 185.415 ;
        RECT 94.990 184.975 95.440 185.085 ;
        RECT 94.315 184.805 95.440 184.975 ;
        RECT 95.715 184.915 95.995 185.585 ;
        RECT 96.165 185.965 96.680 186.375 ;
        RECT 96.165 185.155 96.505 185.965 ;
        RECT 97.255 185.720 97.425 186.385 ;
        RECT 97.820 186.045 98.945 186.215 ;
        RECT 96.675 185.530 97.425 185.720 ;
        RECT 97.595 185.705 98.605 185.875 ;
        RECT 96.165 184.985 97.395 185.155 ;
        RECT 94.315 184.345 94.595 184.805 ;
        RECT 95.610 184.345 95.995 184.915 ;
        RECT 96.440 184.380 96.685 184.985 ;
        RECT 97.595 184.345 97.785 185.705 ;
        RECT 97.955 185.025 98.230 185.505 ;
        RECT 97.955 184.855 98.235 185.025 ;
        RECT 98.435 184.905 98.605 185.705 ;
        RECT 98.775 184.915 98.945 186.045 ;
        RECT 99.115 185.415 99.285 186.385 ;
        RECT 99.795 185.585 100.130 186.555 ;
        RECT 100.395 185.795 100.565 186.555 ;
        RECT 100.395 185.625 101.060 185.795 ;
        RECT 101.245 185.650 101.515 186.555 ;
        RECT 99.115 185.085 99.310 185.415 ;
        RECT 99.535 185.085 99.790 185.415 ;
        RECT 99.535 184.915 99.705 185.085 ;
        RECT 99.960 184.915 100.130 185.585 ;
        RECT 100.890 185.480 101.060 185.625 ;
        RECT 100.325 185.075 100.655 185.445 ;
        RECT 100.890 185.150 101.175 185.480 ;
        RECT 97.955 184.345 98.230 184.855 ;
        RECT 98.775 184.745 99.705 184.915 ;
        RECT 98.775 184.710 98.950 184.745 ;
        RECT 98.420 184.345 98.950 184.710 ;
        RECT 99.875 184.345 100.130 184.915 ;
        RECT 100.890 184.895 101.060 185.150 ;
        RECT 100.395 184.725 101.060 184.895 ;
        RECT 101.345 184.850 101.515 185.650 ;
        RECT 100.395 184.345 100.565 184.725 ;
        RECT 101.255 184.345 101.515 184.850 ;
        RECT 102.585 185.575 102.915 186.555 ;
        RECT 107.780 186.095 108.065 186.555 ;
        RECT 107.780 185.875 108.735 186.095 ;
        RECT 102.585 184.975 102.835 185.575 ;
        RECT 103.005 185.165 103.335 185.415 ;
        RECT 107.665 185.145 108.355 185.705 ;
        RECT 108.525 184.975 108.735 185.875 ;
        RECT 102.585 184.345 102.915 184.975 ;
        RECT 107.780 184.805 108.735 184.975 ;
        RECT 108.905 185.705 109.305 186.555 ;
        RECT 109.495 186.095 109.775 186.555 ;
        RECT 109.495 185.875 110.620 186.095 ;
        RECT 108.905 185.145 110.000 185.705 ;
        RECT 110.170 185.415 110.620 185.875 ;
        RECT 110.790 185.585 111.175 186.555 ;
        RECT 107.780 184.345 108.065 184.805 ;
        RECT 108.905 184.345 109.305 185.145 ;
        RECT 110.170 185.085 110.725 185.415 ;
        RECT 110.170 184.975 110.620 185.085 ;
        RECT 109.495 184.805 110.620 184.975 ;
        RECT 110.895 184.915 111.175 185.585 ;
        RECT 109.495 184.345 109.775 184.805 ;
        RECT 110.790 184.345 111.175 184.915 ;
        RECT 22.195 183.455 22.365 183.835 ;
        RECT 22.195 183.285 22.860 183.455 ;
        RECT 23.055 183.330 23.315 183.835 ;
        RECT 22.125 182.735 22.455 183.105 ;
        RECT 22.690 183.030 22.860 183.285 ;
        RECT 22.690 182.700 22.975 183.030 ;
        RECT 22.690 182.555 22.860 182.700 ;
        RECT 22.195 182.385 22.860 182.555 ;
        RECT 23.145 182.530 23.315 183.330 ;
        RECT 22.195 181.625 22.365 182.385 ;
        RECT 23.045 181.625 23.315 182.530 ;
        RECT 23.485 183.265 23.870 183.835 ;
        RECT 24.885 183.375 25.165 183.835 ;
        RECT 23.485 182.595 23.765 183.265 ;
        RECT 24.040 183.205 25.165 183.375 ;
        RECT 24.040 183.095 24.490 183.205 ;
        RECT 23.935 182.765 24.490 183.095 ;
        RECT 25.355 183.035 25.755 183.835 ;
        RECT 26.595 183.375 26.880 183.835 ;
        RECT 23.485 181.625 23.870 182.595 ;
        RECT 24.040 182.305 24.490 182.765 ;
        RECT 24.660 182.475 25.755 183.035 ;
        RECT 24.040 182.085 25.165 182.305 ;
        RECT 24.885 181.625 25.165 182.085 ;
        RECT 25.355 181.625 25.755 182.475 ;
        RECT 25.925 183.205 26.880 183.375 ;
        RECT 27.280 183.375 27.565 183.835 ;
        RECT 27.280 183.205 28.235 183.375 ;
        RECT 25.925 182.305 26.135 183.205 ;
        RECT 26.305 182.475 26.995 183.035 ;
        RECT 27.165 182.475 27.855 183.035 ;
        RECT 28.025 182.305 28.235 183.205 ;
        RECT 25.925 182.085 26.880 182.305 ;
        RECT 26.595 181.625 26.880 182.085 ;
        RECT 27.280 182.085 28.235 182.305 ;
        RECT 28.405 183.035 28.805 183.835 ;
        RECT 28.995 183.375 29.275 183.835 ;
        RECT 28.995 183.205 30.120 183.375 ;
        RECT 30.290 183.265 30.675 183.835 ;
        RECT 29.670 183.095 30.120 183.205 ;
        RECT 28.405 182.475 29.500 183.035 ;
        RECT 29.670 182.765 30.225 183.095 ;
        RECT 27.280 181.625 27.565 182.085 ;
        RECT 28.405 181.625 28.805 182.475 ;
        RECT 29.670 182.305 30.120 182.765 ;
        RECT 30.395 182.595 30.675 183.265 ;
        RECT 28.995 182.085 30.120 182.305 ;
        RECT 28.995 181.625 29.275 182.085 ;
        RECT 30.290 181.625 30.675 182.595 ;
        RECT 30.850 183.265 31.105 183.835 ;
        RECT 32.030 183.470 32.560 183.835 ;
        RECT 32.030 183.435 32.205 183.470 ;
        RECT 31.275 183.265 32.205 183.435 ;
        RECT 32.750 183.325 33.025 183.835 ;
        RECT 30.850 182.595 31.020 183.265 ;
        RECT 31.275 183.095 31.445 183.265 ;
        RECT 31.190 182.765 31.445 183.095 ;
        RECT 31.670 182.765 31.865 183.095 ;
        RECT 30.850 181.625 31.185 182.595 ;
        RECT 31.695 181.795 31.865 182.765 ;
        RECT 32.035 182.135 32.205 183.265 ;
        RECT 32.375 182.475 32.545 183.275 ;
        RECT 32.745 183.155 33.025 183.325 ;
        RECT 32.750 182.675 33.025 183.155 ;
        RECT 33.195 182.475 33.385 183.835 ;
        RECT 34.295 183.195 34.540 183.800 ;
        RECT 37.860 183.375 38.145 183.835 ;
        RECT 37.860 183.205 38.815 183.375 ;
        RECT 33.585 183.025 34.815 183.195 ;
        RECT 32.375 182.305 33.385 182.475 ;
        RECT 33.555 182.460 34.305 182.650 ;
        RECT 32.035 181.965 33.160 182.135 ;
        RECT 33.555 181.795 33.725 182.460 ;
        RECT 34.475 182.215 34.815 183.025 ;
        RECT 37.745 182.475 38.435 183.035 ;
        RECT 38.605 182.305 38.815 183.205 ;
        RECT 34.300 181.805 34.815 182.215 ;
        RECT 37.860 182.085 38.815 182.305 ;
        RECT 38.985 183.035 39.385 183.835 ;
        RECT 39.575 183.375 39.855 183.835 ;
        RECT 39.575 183.205 40.700 183.375 ;
        RECT 40.870 183.265 41.255 183.835 ;
        RECT 41.975 183.455 42.145 183.835 ;
        RECT 41.975 183.285 42.640 183.455 ;
        RECT 42.835 183.330 43.095 183.835 ;
        RECT 40.250 183.095 40.700 183.205 ;
        RECT 38.985 182.475 40.080 183.035 ;
        RECT 40.250 182.765 40.805 183.095 ;
        RECT 31.695 181.625 33.725 181.795 ;
        RECT 37.860 181.625 38.145 182.085 ;
        RECT 38.985 181.625 39.385 182.475 ;
        RECT 40.250 182.305 40.700 182.765 ;
        RECT 40.975 182.595 41.255 183.265 ;
        RECT 41.905 182.735 42.235 183.105 ;
        RECT 42.470 183.030 42.640 183.285 ;
        RECT 39.575 182.085 40.700 182.305 ;
        RECT 39.575 181.625 39.855 182.085 ;
        RECT 40.870 181.625 41.255 182.595 ;
        RECT 42.470 182.700 42.755 183.030 ;
        RECT 42.470 182.555 42.640 182.700 ;
        RECT 41.975 182.385 42.640 182.555 ;
        RECT 42.925 182.530 43.095 183.330 ;
        RECT 43.380 183.375 43.665 183.835 ;
        RECT 43.380 183.205 44.335 183.375 ;
        RECT 41.975 181.625 42.145 182.385 ;
        RECT 42.825 181.625 43.095 182.530 ;
        RECT 43.265 182.475 43.955 183.035 ;
        RECT 44.125 182.305 44.335 183.205 ;
        RECT 43.380 182.085 44.335 182.305 ;
        RECT 44.505 183.035 44.905 183.835 ;
        RECT 45.095 183.375 45.375 183.835 ;
        RECT 45.095 183.205 46.220 183.375 ;
        RECT 46.390 183.265 46.775 183.835 ;
        RECT 45.770 183.095 46.220 183.205 ;
        RECT 44.505 182.475 45.600 183.035 ;
        RECT 45.770 182.765 46.325 183.095 ;
        RECT 43.380 181.625 43.665 182.085 ;
        RECT 44.505 181.625 44.905 182.475 ;
        RECT 45.770 182.305 46.220 182.765 ;
        RECT 46.495 182.595 46.775 183.265 ;
        RECT 47.060 183.375 47.345 183.835 ;
        RECT 47.060 183.205 48.015 183.375 ;
        RECT 45.095 182.085 46.220 182.305 ;
        RECT 45.095 181.625 45.375 182.085 ;
        RECT 46.390 181.625 46.775 182.595 ;
        RECT 46.945 182.475 47.635 183.035 ;
        RECT 47.805 182.305 48.015 183.205 ;
        RECT 47.060 182.085 48.015 182.305 ;
        RECT 48.185 183.035 48.585 183.835 ;
        RECT 48.775 183.375 49.055 183.835 ;
        RECT 48.775 183.205 49.900 183.375 ;
        RECT 50.070 183.265 50.455 183.835 ;
        RECT 49.450 183.095 49.900 183.205 ;
        RECT 48.185 182.475 49.280 183.035 ;
        RECT 49.450 182.765 50.005 183.095 ;
        RECT 47.060 181.625 47.345 182.085 ;
        RECT 48.185 181.625 48.585 182.475 ;
        RECT 49.450 182.305 49.900 182.765 ;
        RECT 50.175 182.595 50.455 183.265 ;
        RECT 48.775 182.085 49.900 182.305 ;
        RECT 48.775 181.625 49.055 182.085 ;
        RECT 50.070 181.625 50.455 182.595 ;
        RECT 50.630 183.265 50.885 183.835 ;
        RECT 51.810 183.470 52.340 183.835 ;
        RECT 51.810 183.435 51.985 183.470 ;
        RECT 51.055 183.265 51.985 183.435 ;
        RECT 50.630 182.595 50.800 183.265 ;
        RECT 51.055 183.095 51.225 183.265 ;
        RECT 50.970 182.765 51.225 183.095 ;
        RECT 51.450 182.765 51.645 183.095 ;
        RECT 50.630 181.625 50.965 182.595 ;
        RECT 51.475 181.795 51.645 182.765 ;
        RECT 51.815 182.135 51.985 183.265 ;
        RECT 52.155 182.475 52.325 183.275 ;
        RECT 52.530 182.985 52.805 183.835 ;
        RECT 52.525 182.815 52.805 182.985 ;
        RECT 52.530 182.675 52.805 182.815 ;
        RECT 52.975 182.475 53.165 183.835 ;
        RECT 54.075 183.195 54.320 183.800 ;
        RECT 55.665 183.205 55.995 183.835 ;
        RECT 56.720 183.375 57.005 183.835 ;
        RECT 56.720 183.205 57.675 183.375 ;
        RECT 53.365 183.025 54.595 183.195 ;
        RECT 52.155 182.305 53.165 182.475 ;
        RECT 53.335 182.460 54.085 182.650 ;
        RECT 51.815 181.965 52.940 182.135 ;
        RECT 53.335 181.795 53.505 182.460 ;
        RECT 54.255 182.215 54.595 183.025 ;
        RECT 55.245 182.765 55.575 183.015 ;
        RECT 55.745 182.605 55.995 183.205 ;
        RECT 54.080 181.805 54.595 182.215 ;
        RECT 51.475 181.625 53.505 181.795 ;
        RECT 55.665 181.625 55.995 182.605 ;
        RECT 56.605 182.475 57.295 183.035 ;
        RECT 57.465 182.305 57.675 183.205 ;
        RECT 56.720 182.085 57.675 182.305 ;
        RECT 57.845 183.035 58.245 183.835 ;
        RECT 58.435 183.375 58.715 183.835 ;
        RECT 58.435 183.205 59.560 183.375 ;
        RECT 59.730 183.265 60.115 183.835 ;
        RECT 60.375 183.455 60.545 183.835 ;
        RECT 60.375 183.285 61.040 183.455 ;
        RECT 61.235 183.330 61.495 183.835 ;
        RECT 59.110 183.095 59.560 183.205 ;
        RECT 57.845 182.475 58.940 183.035 ;
        RECT 59.110 182.765 59.665 183.095 ;
        RECT 56.720 181.625 57.005 182.085 ;
        RECT 57.845 181.625 58.245 182.475 ;
        RECT 59.110 182.305 59.560 182.765 ;
        RECT 59.835 182.595 60.115 183.265 ;
        RECT 60.305 182.735 60.635 183.105 ;
        RECT 60.870 183.030 61.040 183.285 ;
        RECT 58.435 182.085 59.560 182.305 ;
        RECT 58.435 181.625 58.715 182.085 ;
        RECT 59.730 181.625 60.115 182.595 ;
        RECT 60.870 182.700 61.155 183.030 ;
        RECT 60.870 182.555 61.040 182.700 ;
        RECT 60.375 182.385 61.040 182.555 ;
        RECT 61.325 182.530 61.495 183.330 ;
        RECT 60.375 181.625 60.545 182.385 ;
        RECT 61.225 181.625 61.495 182.530 ;
        RECT 61.665 183.330 61.925 183.835 ;
        RECT 62.615 183.455 62.785 183.835 ;
        RECT 61.665 182.530 61.835 183.330 ;
        RECT 62.120 183.285 62.785 183.455 ;
        RECT 73.015 183.435 73.215 183.790 ;
        RECT 73.885 183.435 74.085 183.780 ;
        RECT 62.120 183.030 62.290 183.285 ;
        RECT 72.245 183.265 74.085 183.435 ;
        RECT 74.820 183.435 74.990 183.685 ;
        RECT 74.820 183.265 75.295 183.435 ;
        RECT 62.005 182.700 62.290 183.030 ;
        RECT 62.525 182.735 62.855 183.105 ;
        RECT 62.120 182.555 62.290 182.700 ;
        RECT 61.665 181.625 61.935 182.530 ;
        RECT 62.120 182.385 62.785 182.555 ;
        RECT 62.615 181.625 62.785 182.385 ;
        RECT 72.245 181.640 72.505 183.265 ;
        RECT 72.685 182.295 72.905 183.095 ;
        RECT 73.145 182.475 73.445 183.095 ;
        RECT 73.615 182.475 73.945 183.095 ;
        RECT 74.115 182.475 74.435 183.095 ;
        RECT 74.605 182.475 74.955 183.095 ;
        RECT 75.125 182.295 75.295 183.265 ;
        RECT 76.130 183.225 76.630 183.835 ;
        RECT 75.925 182.765 76.275 183.015 ;
        RECT 76.460 182.595 76.630 183.225 ;
        RECT 77.260 183.355 77.590 183.835 ;
        RECT 78.155 183.355 78.485 183.835 ;
        RECT 77.260 183.185 78.485 183.355 ;
        RECT 79.095 183.205 79.435 183.835 ;
        RECT 76.800 182.815 77.130 183.015 ;
        RECT 77.300 182.815 77.630 183.015 ;
        RECT 77.800 182.815 78.220 183.015 ;
        RECT 78.395 182.845 79.090 183.015 ;
        RECT 78.395 182.595 78.565 182.845 ;
        RECT 79.260 182.595 79.435 183.205 ;
        RECT 72.685 182.085 75.295 182.295 ;
        RECT 76.130 182.425 78.565 182.595 ;
        RECT 76.130 181.625 76.460 182.425 ;
        RECT 77.260 181.625 77.590 182.425 ;
        RECT 79.095 181.625 79.435 182.595 ;
        RECT 79.610 183.295 79.865 183.825 ;
        RECT 80.585 183.625 81.655 183.795 ;
        RECT 79.610 182.645 79.820 183.295 ;
        RECT 80.585 183.270 80.905 183.625 ;
        RECT 80.580 183.095 80.905 183.270 ;
        RECT 79.990 182.795 80.905 183.095 ;
        RECT 81.075 183.055 81.315 183.455 ;
        RECT 81.485 183.395 81.655 183.625 ;
        RECT 82.185 183.555 83.135 183.835 ;
        RECT 83.355 183.645 83.705 183.815 ;
        RECT 81.485 183.225 82.015 183.395 ;
        RECT 79.990 182.765 80.730 182.795 ;
        RECT 79.610 181.765 79.865 182.645 ;
        RECT 80.560 182.175 80.730 182.765 ;
        RECT 81.075 182.685 81.615 183.055 ;
        RECT 81.795 182.945 82.015 183.225 ;
        RECT 82.185 182.775 82.355 183.555 ;
        RECT 81.950 182.605 82.355 182.775 ;
        RECT 82.525 182.765 82.875 183.385 ;
        RECT 81.950 182.515 82.120 182.605 ;
        RECT 83.045 182.595 83.255 183.385 ;
        RECT 80.900 182.345 82.120 182.515 ;
        RECT 82.580 182.435 83.255 182.595 ;
        RECT 80.560 182.005 81.360 182.175 ;
        RECT 81.190 181.715 81.360 182.005 ;
        RECT 81.950 181.965 82.120 182.345 ;
        RECT 82.290 182.425 83.255 182.435 ;
        RECT 83.445 183.255 83.705 183.645 ;
        RECT 85.120 183.615 85.975 183.785 ;
        RECT 86.180 183.615 86.675 183.785 ;
        RECT 83.445 182.565 83.615 183.255 ;
        RECT 83.785 182.905 83.955 183.085 ;
        RECT 84.125 183.075 84.915 183.325 ;
        RECT 85.120 182.905 85.290 183.615 ;
        RECT 85.460 183.105 85.815 183.325 ;
        RECT 83.785 182.735 85.475 182.905 ;
        RECT 82.290 182.135 82.750 182.425 ;
        RECT 83.445 182.395 84.945 182.565 ;
        RECT 83.445 182.255 83.615 182.395 ;
        RECT 83.055 182.085 83.615 182.255 ;
        RECT 81.950 181.625 82.820 181.965 ;
        RECT 83.055 181.625 83.225 182.085 ;
        RECT 84.060 182.055 85.135 182.225 ;
        RECT 84.060 181.715 84.230 182.055 ;
        RECT 84.965 181.715 85.135 182.055 ;
        RECT 85.305 181.955 85.475 182.735 ;
        RECT 85.645 182.515 85.815 183.105 ;
        RECT 85.985 182.705 86.335 183.325 ;
        RECT 85.645 182.125 86.110 182.515 ;
        RECT 86.505 182.255 86.675 183.615 ;
        RECT 86.845 182.425 87.305 183.475 ;
        RECT 86.280 182.085 86.675 182.255 ;
        RECT 86.280 181.955 86.450 182.085 ;
        RECT 85.305 181.625 85.985 181.955 ;
        RECT 86.200 181.625 86.450 181.955 ;
        RECT 87.040 181.640 87.365 182.425 ;
        RECT 87.535 181.625 87.705 183.745 ;
        RECT 88.375 183.455 88.630 183.745 ;
        RECT 87.880 183.285 88.630 183.455 ;
        RECT 90.185 183.330 90.445 183.835 ;
        RECT 91.135 183.455 91.305 183.835 ;
        RECT 87.880 182.295 88.110 183.285 ;
        RECT 88.280 182.465 88.630 183.115 ;
        RECT 90.185 182.530 90.355 183.330 ;
        RECT 90.640 183.285 91.305 183.455 ;
        RECT 92.490 183.295 92.745 183.825 ;
        RECT 93.465 183.625 94.535 183.795 ;
        RECT 90.640 183.030 90.810 183.285 ;
        RECT 90.525 182.700 90.810 183.030 ;
        RECT 91.045 182.735 91.375 183.105 ;
        RECT 90.640 182.555 90.810 182.700 ;
        RECT 92.490 182.645 92.700 183.295 ;
        RECT 93.465 183.270 93.785 183.625 ;
        RECT 93.460 183.095 93.785 183.270 ;
        RECT 92.870 182.795 93.785 183.095 ;
        RECT 93.955 183.055 94.195 183.455 ;
        RECT 94.365 183.395 94.535 183.625 ;
        RECT 95.065 183.555 96.015 183.835 ;
        RECT 96.235 183.645 96.585 183.815 ;
        RECT 94.365 183.225 94.895 183.395 ;
        RECT 92.870 182.765 93.610 182.795 ;
        RECT 87.880 182.125 88.630 182.295 ;
        RECT 88.375 181.625 88.630 182.125 ;
        RECT 90.185 181.625 90.455 182.530 ;
        RECT 90.640 182.385 91.305 182.555 ;
        RECT 91.135 181.625 91.305 182.385 ;
        RECT 92.490 181.765 92.745 182.645 ;
        RECT 93.440 182.175 93.610 182.765 ;
        RECT 93.955 182.685 94.495 183.055 ;
        RECT 94.675 182.945 94.895 183.225 ;
        RECT 95.065 182.775 95.235 183.555 ;
        RECT 94.830 182.605 95.235 182.775 ;
        RECT 95.405 182.765 95.755 183.385 ;
        RECT 94.830 182.515 95.000 182.605 ;
        RECT 95.925 182.595 96.135 183.385 ;
        RECT 93.780 182.345 95.000 182.515 ;
        RECT 95.460 182.435 96.135 182.595 ;
        RECT 93.440 182.005 94.240 182.175 ;
        RECT 94.070 181.715 94.240 182.005 ;
        RECT 94.830 181.965 95.000 182.345 ;
        RECT 95.170 182.425 96.135 182.435 ;
        RECT 96.325 183.255 96.585 183.645 ;
        RECT 98.000 183.615 98.855 183.785 ;
        RECT 99.060 183.615 99.555 183.785 ;
        RECT 96.325 182.565 96.495 183.255 ;
        RECT 96.665 182.905 96.835 183.085 ;
        RECT 97.005 183.075 97.795 183.325 ;
        RECT 98.000 182.905 98.170 183.615 ;
        RECT 98.340 183.105 98.695 183.325 ;
        RECT 96.665 182.735 98.355 182.905 ;
        RECT 95.170 182.135 95.630 182.425 ;
        RECT 96.325 182.395 97.825 182.565 ;
        RECT 96.325 182.255 96.495 182.395 ;
        RECT 95.935 182.085 96.495 182.255 ;
        RECT 94.830 181.625 95.700 181.965 ;
        RECT 95.935 181.625 96.105 182.085 ;
        RECT 96.940 182.055 98.015 182.225 ;
        RECT 96.940 181.715 97.110 182.055 ;
        RECT 97.845 181.715 98.015 182.055 ;
        RECT 98.185 181.955 98.355 182.735 ;
        RECT 98.525 182.515 98.695 183.105 ;
        RECT 98.865 182.705 99.215 183.325 ;
        RECT 98.525 182.125 98.990 182.515 ;
        RECT 99.385 182.255 99.555 183.615 ;
        RECT 99.725 182.425 100.185 183.475 ;
        RECT 99.160 182.085 99.555 182.255 ;
        RECT 99.160 181.955 99.330 182.085 ;
        RECT 98.185 181.625 98.865 181.955 ;
        RECT 99.080 181.625 99.330 181.955 ;
        RECT 99.920 181.640 100.245 182.425 ;
        RECT 100.415 181.625 100.585 183.745 ;
        RECT 101.255 183.455 101.510 183.745 ;
        RECT 100.760 183.285 101.510 183.455 ;
        RECT 100.760 182.295 100.990 183.285 ;
        RECT 102.610 183.265 102.865 183.835 ;
        RECT 103.790 183.470 104.320 183.835 ;
        RECT 103.790 183.435 103.965 183.470 ;
        RECT 103.035 183.265 103.965 183.435 ;
        RECT 101.160 182.465 101.510 183.115 ;
        RECT 102.610 182.595 102.780 183.265 ;
        RECT 103.035 183.095 103.205 183.265 ;
        RECT 102.950 182.765 103.205 183.095 ;
        RECT 103.430 182.765 103.625 183.095 ;
        RECT 100.760 182.125 101.510 182.295 ;
        RECT 101.255 181.625 101.510 182.125 ;
        RECT 102.610 181.625 102.945 182.595 ;
        RECT 103.455 181.795 103.625 182.765 ;
        RECT 103.795 182.135 103.965 183.265 ;
        RECT 104.135 182.475 104.305 183.275 ;
        RECT 104.510 182.985 104.785 183.835 ;
        RECT 104.505 182.815 104.785 182.985 ;
        RECT 104.510 182.675 104.785 182.815 ;
        RECT 104.955 182.475 105.145 183.835 ;
        RECT 106.055 183.195 106.300 183.800 ;
        RECT 106.745 183.265 107.130 183.835 ;
        RECT 108.145 183.375 108.425 183.835 ;
        RECT 105.345 183.025 106.575 183.195 ;
        RECT 104.135 182.305 105.145 182.475 ;
        RECT 105.315 182.460 106.065 182.650 ;
        RECT 103.795 181.965 104.920 182.135 ;
        RECT 105.315 181.795 105.485 182.460 ;
        RECT 106.235 182.215 106.575 183.025 ;
        RECT 106.060 181.805 106.575 182.215 ;
        RECT 106.745 182.595 107.025 183.265 ;
        RECT 107.300 183.205 108.425 183.375 ;
        RECT 107.300 183.095 107.750 183.205 ;
        RECT 107.195 182.765 107.750 183.095 ;
        RECT 108.615 183.035 109.015 183.835 ;
        RECT 109.855 183.375 110.140 183.835 ;
        RECT 103.455 181.625 105.485 181.795 ;
        RECT 106.745 181.625 107.130 182.595 ;
        RECT 107.300 182.305 107.750 182.765 ;
        RECT 107.920 182.475 109.015 183.035 ;
        RECT 107.300 182.085 108.425 182.305 ;
        RECT 108.145 181.625 108.425 182.085 ;
        RECT 108.615 181.625 109.015 182.475 ;
        RECT 109.185 183.205 110.140 183.375 ;
        RECT 109.185 182.305 109.395 183.205 ;
        RECT 110.700 183.195 110.945 183.800 ;
        RECT 109.565 182.475 110.255 183.035 ;
        RECT 110.425 183.025 111.655 183.195 ;
        RECT 109.185 182.085 110.140 182.305 ;
        RECT 109.855 181.625 110.140 182.085 ;
        RECT 110.425 182.215 110.765 183.025 ;
        RECT 110.935 182.460 111.685 182.650 ;
        RECT 110.425 181.805 110.940 182.215 ;
        RECT 111.515 181.795 111.685 182.460 ;
        RECT 111.855 182.475 112.045 183.835 ;
        RECT 112.215 182.985 112.490 183.835 ;
        RECT 112.680 183.470 113.210 183.835 ;
        RECT 113.035 183.435 113.210 183.470 ;
        RECT 112.215 182.815 112.495 182.985 ;
        RECT 112.215 182.675 112.490 182.815 ;
        RECT 112.695 182.475 112.865 183.275 ;
        RECT 111.855 182.305 112.865 182.475 ;
        RECT 113.035 183.265 113.965 183.435 ;
        RECT 114.135 183.265 114.390 183.835 ;
        RECT 113.035 182.135 113.205 183.265 ;
        RECT 113.795 183.095 113.965 183.265 ;
        RECT 112.080 181.965 113.205 182.135 ;
        RECT 113.375 182.765 113.570 183.095 ;
        RECT 113.795 182.765 114.050 183.095 ;
        RECT 113.375 181.795 113.545 182.765 ;
        RECT 114.220 182.595 114.390 183.265 ;
        RECT 111.515 181.625 113.545 181.795 ;
        RECT 114.055 181.625 114.390 182.595 ;
        RECT 115.490 183.295 115.745 183.825 ;
        RECT 116.465 183.625 117.535 183.795 ;
        RECT 115.490 182.645 115.700 183.295 ;
        RECT 116.465 183.270 116.785 183.625 ;
        RECT 116.460 183.095 116.785 183.270 ;
        RECT 115.870 182.795 116.785 183.095 ;
        RECT 116.955 183.055 117.195 183.455 ;
        RECT 117.365 183.395 117.535 183.625 ;
        RECT 118.065 183.555 119.015 183.835 ;
        RECT 119.235 183.645 119.585 183.815 ;
        RECT 117.365 183.225 117.895 183.395 ;
        RECT 115.870 182.765 116.610 182.795 ;
        RECT 115.490 181.765 115.745 182.645 ;
        RECT 116.440 182.175 116.610 182.765 ;
        RECT 116.955 182.685 117.495 183.055 ;
        RECT 117.675 182.945 117.895 183.225 ;
        RECT 118.065 182.775 118.235 183.555 ;
        RECT 117.830 182.605 118.235 182.775 ;
        RECT 118.405 182.765 118.755 183.385 ;
        RECT 117.830 182.515 118.000 182.605 ;
        RECT 118.925 182.595 119.135 183.385 ;
        RECT 116.780 182.345 118.000 182.515 ;
        RECT 118.460 182.435 119.135 182.595 ;
        RECT 116.440 182.005 117.240 182.175 ;
        RECT 117.070 181.715 117.240 182.005 ;
        RECT 117.830 181.965 118.000 182.345 ;
        RECT 118.170 182.425 119.135 182.435 ;
        RECT 119.325 183.255 119.585 183.645 ;
        RECT 121.000 183.615 121.855 183.785 ;
        RECT 122.060 183.615 122.555 183.785 ;
        RECT 119.325 182.565 119.495 183.255 ;
        RECT 119.665 182.905 119.835 183.085 ;
        RECT 120.005 183.075 120.795 183.325 ;
        RECT 121.000 182.905 121.170 183.615 ;
        RECT 121.340 183.105 121.695 183.325 ;
        RECT 119.665 182.735 121.355 182.905 ;
        RECT 118.170 182.135 118.630 182.425 ;
        RECT 119.325 182.395 120.825 182.565 ;
        RECT 119.325 182.255 119.495 182.395 ;
        RECT 118.935 182.085 119.495 182.255 ;
        RECT 117.830 181.625 118.700 181.965 ;
        RECT 118.935 181.625 119.105 182.085 ;
        RECT 119.940 182.055 121.015 182.225 ;
        RECT 119.940 181.715 120.110 182.055 ;
        RECT 120.845 181.715 121.015 182.055 ;
        RECT 121.185 181.955 121.355 182.735 ;
        RECT 121.525 182.515 121.695 183.105 ;
        RECT 121.865 182.705 122.215 183.325 ;
        RECT 121.525 182.125 121.990 182.515 ;
        RECT 122.385 182.255 122.555 183.615 ;
        RECT 122.725 182.425 123.185 183.475 ;
        RECT 122.160 182.085 122.555 182.255 ;
        RECT 122.160 181.955 122.330 182.085 ;
        RECT 121.185 181.625 121.865 181.955 ;
        RECT 122.080 181.625 122.330 181.955 ;
        RECT 122.920 181.640 123.245 182.425 ;
        RECT 123.415 181.625 123.585 183.745 ;
        RECT 124.255 183.455 124.510 183.745 ;
        RECT 123.760 183.285 124.510 183.455 ;
        RECT 123.760 182.295 123.990 183.285 ;
        RECT 124.160 182.465 124.510 183.115 ;
        RECT 123.760 182.125 124.510 182.295 ;
        RECT 124.255 181.625 124.510 182.125 ;
        RECT 24.870 180.615 25.125 181.115 ;
        RECT 24.870 180.445 25.620 180.615 ;
        RECT 24.870 179.625 25.220 180.275 ;
        RECT 25.390 179.455 25.620 180.445 ;
        RECT 24.870 179.285 25.620 179.455 ;
        RECT 24.870 178.995 25.125 179.285 ;
        RECT 25.795 178.995 25.965 181.115 ;
        RECT 26.135 180.315 26.460 181.100 ;
        RECT 27.050 180.785 27.300 181.115 ;
        RECT 27.515 180.785 28.195 181.115 ;
        RECT 27.050 180.655 27.220 180.785 ;
        RECT 26.825 180.485 27.220 180.655 ;
        RECT 26.195 179.265 26.655 180.315 ;
        RECT 26.825 179.125 26.995 180.485 ;
        RECT 27.390 180.225 27.855 180.615 ;
        RECT 27.165 179.415 27.515 180.035 ;
        RECT 27.685 179.635 27.855 180.225 ;
        RECT 28.025 180.005 28.195 180.785 ;
        RECT 28.365 180.685 28.535 181.025 ;
        RECT 29.270 180.685 29.440 181.025 ;
        RECT 28.365 180.515 29.440 180.685 ;
        RECT 30.275 180.655 30.445 181.115 ;
        RECT 30.680 180.775 31.550 181.115 ;
        RECT 29.885 180.485 30.445 180.655 ;
        RECT 29.885 180.345 30.055 180.485 ;
        RECT 28.555 180.175 30.055 180.345 ;
        RECT 30.750 180.315 31.210 180.605 ;
        RECT 28.025 179.835 29.715 180.005 ;
        RECT 27.685 179.415 28.040 179.635 ;
        RECT 28.210 179.125 28.380 179.835 ;
        RECT 28.585 179.415 29.375 179.665 ;
        RECT 29.545 179.655 29.715 179.835 ;
        RECT 29.885 179.485 30.055 180.175 ;
        RECT 26.825 178.955 27.320 179.125 ;
        RECT 27.525 178.955 28.380 179.125 ;
        RECT 29.795 179.095 30.055 179.485 ;
        RECT 30.245 180.305 31.210 180.315 ;
        RECT 31.380 180.395 31.550 180.775 ;
        RECT 32.140 180.735 32.310 181.025 ;
        RECT 32.140 180.565 32.940 180.735 ;
        RECT 30.245 180.145 30.920 180.305 ;
        RECT 31.380 180.225 32.600 180.395 ;
        RECT 30.245 179.355 30.455 180.145 ;
        RECT 31.380 180.135 31.550 180.225 ;
        RECT 30.625 179.355 30.975 179.975 ;
        RECT 31.145 179.965 31.550 180.135 ;
        RECT 31.145 179.185 31.315 179.965 ;
        RECT 31.485 179.515 31.705 179.795 ;
        RECT 31.885 179.685 32.425 180.055 ;
        RECT 32.770 179.975 32.940 180.565 ;
        RECT 33.635 180.095 33.890 180.975 ;
        RECT 34.640 180.655 34.925 181.115 ;
        RECT 34.640 180.435 35.595 180.655 ;
        RECT 32.770 179.945 33.510 179.975 ;
        RECT 31.485 179.345 32.015 179.515 ;
        RECT 29.795 178.925 30.145 179.095 ;
        RECT 30.365 178.905 31.315 179.185 ;
        RECT 31.845 179.115 32.015 179.345 ;
        RECT 32.185 179.285 32.425 179.685 ;
        RECT 32.595 179.645 33.510 179.945 ;
        RECT 32.595 179.470 32.920 179.645 ;
        RECT 32.595 179.115 32.915 179.470 ;
        RECT 33.680 179.445 33.890 180.095 ;
        RECT 34.525 179.705 35.215 180.265 ;
        RECT 35.385 179.535 35.595 180.435 ;
        RECT 31.845 178.945 32.915 179.115 ;
        RECT 33.635 178.915 33.890 179.445 ;
        RECT 34.640 179.365 35.595 179.535 ;
        RECT 35.765 180.265 36.165 181.115 ;
        RECT 36.355 180.655 36.635 181.115 ;
        RECT 36.355 180.435 37.480 180.655 ;
        RECT 35.765 179.705 36.860 180.265 ;
        RECT 37.030 179.975 37.480 180.435 ;
        RECT 37.650 180.145 38.035 181.115 ;
        RECT 34.640 178.905 34.925 179.365 ;
        RECT 35.765 178.905 36.165 179.705 ;
        RECT 37.030 179.645 37.585 179.975 ;
        RECT 37.030 179.535 37.480 179.645 ;
        RECT 36.355 179.365 37.480 179.535 ;
        RECT 37.755 179.475 38.035 180.145 ;
        RECT 36.355 178.905 36.635 179.365 ;
        RECT 37.650 178.905 38.035 179.475 ;
        RECT 38.665 180.210 38.935 181.115 ;
        RECT 39.615 180.355 39.785 181.115 ;
        RECT 46.600 180.655 46.885 181.115 ;
        RECT 46.600 180.435 47.555 180.655 ;
        RECT 38.665 179.410 38.835 180.210 ;
        RECT 39.120 180.185 39.785 180.355 ;
        RECT 39.120 180.040 39.290 180.185 ;
        RECT 39.005 179.710 39.290 180.040 ;
        RECT 39.120 179.455 39.290 179.710 ;
        RECT 39.525 179.635 39.855 180.005 ;
        RECT 46.485 179.705 47.175 180.265 ;
        RECT 47.345 179.535 47.555 180.435 ;
        RECT 38.665 178.905 38.925 179.410 ;
        RECT 39.120 179.285 39.785 179.455 ;
        RECT 39.615 178.905 39.785 179.285 ;
        RECT 46.600 179.365 47.555 179.535 ;
        RECT 47.725 180.265 48.125 181.115 ;
        RECT 48.315 180.655 48.595 181.115 ;
        RECT 48.315 180.435 49.440 180.655 ;
        RECT 47.725 179.705 48.820 180.265 ;
        RECT 48.990 179.975 49.440 180.435 ;
        RECT 49.610 180.145 49.995 181.115 ;
        RECT 51.660 180.655 51.945 181.115 ;
        RECT 51.660 180.435 52.615 180.655 ;
        RECT 46.600 178.905 46.885 179.365 ;
        RECT 47.725 178.905 48.125 179.705 ;
        RECT 48.990 179.645 49.545 179.975 ;
        RECT 48.990 179.535 49.440 179.645 ;
        RECT 48.315 179.365 49.440 179.535 ;
        RECT 49.715 179.475 49.995 180.145 ;
        RECT 51.545 179.705 52.235 180.265 ;
        RECT 52.405 179.535 52.615 180.435 ;
        RECT 48.315 178.905 48.595 179.365 ;
        RECT 49.610 178.905 49.995 179.475 ;
        RECT 51.660 179.365 52.615 179.535 ;
        RECT 52.785 180.265 53.185 181.115 ;
        RECT 53.375 180.655 53.655 181.115 ;
        RECT 53.375 180.435 54.500 180.655 ;
        RECT 52.785 179.705 53.880 180.265 ;
        RECT 54.050 179.975 54.500 180.435 ;
        RECT 54.670 180.145 55.055 181.115 ;
        RECT 51.660 178.905 51.945 179.365 ;
        RECT 52.785 178.905 53.185 179.705 ;
        RECT 54.050 179.645 54.605 179.975 ;
        RECT 54.050 179.535 54.500 179.645 ;
        RECT 53.375 179.365 54.500 179.535 ;
        RECT 54.775 179.475 55.055 180.145 ;
        RECT 53.375 178.905 53.655 179.365 ;
        RECT 54.670 178.905 55.055 179.475 ;
        RECT 55.230 180.095 55.485 180.975 ;
        RECT 56.810 180.735 56.980 181.025 ;
        RECT 56.180 180.565 56.980 180.735 ;
        RECT 57.570 180.775 58.440 181.115 ;
        RECT 55.230 179.445 55.440 180.095 ;
        RECT 56.180 179.975 56.350 180.565 ;
        RECT 57.570 180.395 57.740 180.775 ;
        RECT 58.675 180.655 58.845 181.115 ;
        RECT 59.680 180.685 59.850 181.025 ;
        RECT 60.585 180.685 60.755 181.025 ;
        RECT 56.520 180.225 57.740 180.395 ;
        RECT 57.910 180.315 58.370 180.605 ;
        RECT 58.675 180.485 59.235 180.655 ;
        RECT 59.680 180.515 60.755 180.685 ;
        RECT 60.925 180.785 61.605 181.115 ;
        RECT 61.820 180.785 62.070 181.115 ;
        RECT 59.065 180.345 59.235 180.485 ;
        RECT 57.910 180.305 58.875 180.315 ;
        RECT 57.570 180.135 57.740 180.225 ;
        RECT 58.200 180.145 58.875 180.305 ;
        RECT 55.610 179.945 56.350 179.975 ;
        RECT 55.610 179.645 56.525 179.945 ;
        RECT 56.200 179.470 56.525 179.645 ;
        RECT 55.230 178.915 55.485 179.445 ;
        RECT 56.205 179.115 56.525 179.470 ;
        RECT 56.695 179.685 57.235 180.055 ;
        RECT 57.570 179.965 57.975 180.135 ;
        RECT 56.695 179.285 56.935 179.685 ;
        RECT 57.415 179.515 57.635 179.795 ;
        RECT 57.105 179.345 57.635 179.515 ;
        RECT 57.105 179.115 57.275 179.345 ;
        RECT 56.205 178.945 57.275 179.115 ;
        RECT 57.805 179.185 57.975 179.965 ;
        RECT 58.145 179.355 58.495 179.975 ;
        RECT 58.665 179.355 58.875 180.145 ;
        RECT 59.065 180.175 60.565 180.345 ;
        RECT 59.065 179.485 59.235 180.175 ;
        RECT 60.925 180.005 61.095 180.785 ;
        RECT 61.900 180.655 62.070 180.785 ;
        RECT 59.405 179.835 61.095 180.005 ;
        RECT 61.265 180.225 61.730 180.615 ;
        RECT 61.900 180.485 62.295 180.655 ;
        RECT 59.405 179.655 59.575 179.835 ;
        RECT 57.805 178.905 58.755 179.185 ;
        RECT 59.065 179.095 59.325 179.485 ;
        RECT 59.745 179.415 60.535 179.665 ;
        RECT 58.975 178.925 59.325 179.095 ;
        RECT 60.740 179.125 60.910 179.835 ;
        RECT 61.265 179.635 61.435 180.225 ;
        RECT 61.080 179.415 61.435 179.635 ;
        RECT 61.605 179.415 61.955 180.035 ;
        RECT 62.125 179.125 62.295 180.485 ;
        RECT 62.660 180.315 62.985 181.100 ;
        RECT 62.465 179.265 62.925 180.315 ;
        RECT 60.740 178.955 61.595 179.125 ;
        RECT 61.800 178.955 62.295 179.125 ;
        RECT 63.155 178.995 63.325 181.115 ;
        RECT 63.995 180.615 64.250 181.115 ;
        RECT 63.500 180.445 64.250 180.615 ;
        RECT 63.500 179.455 63.730 180.445 ;
        RECT 63.900 179.625 64.250 180.275 ;
        RECT 65.325 180.135 65.655 181.115 ;
        RECT 66.705 180.210 66.960 181.115 ;
        RECT 67.675 180.355 67.845 181.115 ;
        RECT 65.325 179.535 65.575 180.135 ;
        RECT 65.745 179.725 66.075 179.975 ;
        RECT 63.500 179.285 64.250 179.455 ;
        RECT 63.995 178.995 64.250 179.285 ;
        RECT 65.325 178.905 65.655 179.535 ;
        RECT 66.705 179.480 66.875 180.210 ;
        RECT 67.130 180.185 67.845 180.355 ;
        RECT 67.130 179.975 67.300 180.185 ;
        RECT 67.045 179.645 67.300 179.975 ;
        RECT 66.705 178.905 66.960 179.480 ;
        RECT 67.130 179.455 67.300 179.645 ;
        RECT 67.580 179.635 67.935 180.005 ;
        RECT 68.105 179.475 68.365 181.100 ;
        RECT 68.545 180.445 71.155 180.655 ;
        RECT 68.545 179.645 68.765 180.445 ;
        RECT 69.005 179.645 69.305 180.265 ;
        RECT 69.475 179.645 69.805 180.265 ;
        RECT 69.975 179.645 70.295 180.265 ;
        RECT 70.465 179.645 70.815 180.265 ;
        RECT 70.985 179.475 71.155 180.445 ;
        RECT 67.130 179.285 67.845 179.455 ;
        RECT 68.105 179.305 69.945 179.475 ;
        RECT 67.675 178.905 67.845 179.285 ;
        RECT 68.875 178.950 69.075 179.305 ;
        RECT 69.745 178.960 69.945 179.305 ;
        RECT 70.680 179.305 71.155 179.475 ;
        RECT 70.680 179.055 70.850 179.305 ;
        RECT 71.325 178.905 71.585 181.115 ;
        RECT 72.510 180.735 72.680 181.115 ;
        RECT 73.465 180.735 73.635 181.115 ;
        RECT 74.425 180.735 74.615 181.115 ;
        RECT 75.495 180.785 75.755 181.115 ;
        RECT 71.755 180.565 73.705 180.735 ;
        RECT 71.755 179.645 71.925 180.565 ;
        RECT 72.295 179.975 72.490 180.285 ;
        RECT 72.760 179.975 72.945 180.285 ;
        RECT 72.235 179.645 72.490 179.975 ;
        RECT 72.715 179.645 72.945 179.975 ;
        RECT 72.295 179.070 72.490 179.645 ;
        RECT 72.760 179.065 72.945 179.645 ;
        RECT 73.195 179.075 73.365 179.975 ;
        RECT 73.535 179.575 73.705 180.565 ;
        RECT 73.875 180.565 74.615 180.735 ;
        RECT 73.875 180.055 74.045 180.565 ;
        RECT 74.215 180.225 74.795 180.395 ;
        RECT 75.065 180.275 75.415 180.605 ;
        RECT 74.625 180.105 74.795 180.225 ;
        RECT 75.585 180.105 75.755 180.785 ;
        RECT 73.875 179.885 74.445 180.055 ;
        RECT 74.625 179.935 75.755 180.105 ;
        RECT 73.535 179.245 74.085 179.575 ;
        RECT 74.275 179.405 74.445 179.885 ;
        RECT 74.615 179.595 75.235 179.765 ;
        RECT 75.025 179.415 75.235 179.595 ;
        RECT 74.275 179.075 74.675 179.405 ;
        RECT 75.585 179.235 75.755 179.935 ;
        RECT 76.385 179.475 76.645 181.100 ;
        RECT 80.695 180.945 82.725 181.115 ;
        RECT 76.825 180.445 79.435 180.655 ;
        RECT 76.825 179.645 77.045 180.445 ;
        RECT 77.285 179.645 77.585 180.265 ;
        RECT 77.755 179.645 78.085 180.265 ;
        RECT 78.255 179.645 78.575 180.265 ;
        RECT 78.745 179.645 79.095 180.265 ;
        RECT 79.265 179.475 79.435 180.445 ;
        RECT 79.605 180.525 80.120 180.935 ;
        RECT 79.605 179.715 79.945 180.525 ;
        RECT 80.695 180.280 80.865 180.945 ;
        RECT 81.260 180.605 82.385 180.775 ;
        RECT 80.115 180.090 80.865 180.280 ;
        RECT 81.035 180.265 82.045 180.435 ;
        RECT 79.605 179.545 80.835 179.715 ;
        RECT 76.385 179.305 78.225 179.475 ;
        RECT 73.195 178.905 74.675 179.075 ;
        RECT 75.495 178.905 75.755 179.235 ;
        RECT 77.155 178.950 77.355 179.305 ;
        RECT 78.025 178.960 78.225 179.305 ;
        RECT 78.960 179.305 79.435 179.475 ;
        RECT 78.960 179.055 79.130 179.305 ;
        RECT 79.880 178.940 80.125 179.545 ;
        RECT 81.035 178.905 81.225 180.265 ;
        RECT 81.395 179.245 81.670 180.065 ;
        RECT 81.875 179.465 82.045 180.265 ;
        RECT 82.215 179.475 82.385 180.605 ;
        RECT 82.555 179.975 82.725 180.945 ;
        RECT 83.235 180.145 83.570 181.115 ;
        RECT 82.555 179.645 82.750 179.975 ;
        RECT 82.975 179.645 83.230 179.975 ;
        RECT 82.975 179.475 83.145 179.645 ;
        RECT 83.400 179.475 83.570 180.145 ;
        RECT 84.230 179.975 84.475 181.115 ;
        RECT 85.090 179.975 85.340 181.110 ;
        RECT 85.940 180.385 86.200 181.110 ;
        RECT 86.800 180.385 87.060 181.110 ;
        RECT 87.660 180.385 87.920 181.110 ;
        RECT 88.520 180.385 88.780 181.110 ;
        RECT 89.365 180.385 89.625 181.110 ;
        RECT 90.225 180.385 90.485 181.110 ;
        RECT 91.085 180.385 91.345 181.110 ;
        RECT 85.940 180.370 91.345 180.385 ;
        RECT 91.955 180.370 92.245 181.110 ;
        RECT 94.440 180.655 94.725 181.115 ;
        RECT 94.440 180.435 95.395 180.655 ;
        RECT 85.940 180.145 92.685 180.370 ;
        RECT 82.215 179.305 83.145 179.475 ;
        RECT 82.215 179.270 82.390 179.305 ;
        RECT 81.395 179.075 81.675 179.245 ;
        RECT 81.395 178.905 81.670 179.075 ;
        RECT 81.860 178.905 82.390 179.270 ;
        RECT 83.315 178.905 83.570 179.475 ;
        RECT 83.745 179.415 84.060 179.975 ;
        RECT 84.230 179.725 91.350 179.975 ;
        RECT 84.230 178.915 84.480 179.725 ;
        RECT 85.090 178.915 85.340 179.725 ;
        RECT 91.520 179.555 92.685 180.145 ;
        RECT 94.325 179.705 95.015 180.265 ;
        RECT 85.940 179.385 92.685 179.555 ;
        RECT 95.185 179.535 95.395 180.435 ;
        RECT 85.940 178.930 86.200 179.385 ;
        RECT 86.800 178.930 87.060 179.385 ;
        RECT 87.660 178.930 87.920 179.385 ;
        RECT 88.505 178.930 88.780 179.385 ;
        RECT 89.365 178.930 89.625 179.385 ;
        RECT 90.225 178.930 90.485 179.385 ;
        RECT 91.085 178.930 91.345 179.385 ;
        RECT 91.955 178.930 92.215 179.385 ;
        RECT 94.440 179.365 95.395 179.535 ;
        RECT 95.565 180.265 95.965 181.115 ;
        RECT 96.155 180.655 96.435 181.115 ;
        RECT 96.155 180.435 97.280 180.655 ;
        RECT 95.565 179.705 96.660 180.265 ;
        RECT 96.830 179.975 97.280 180.435 ;
        RECT 97.450 180.145 97.835 181.115 ;
        RECT 98.120 180.655 98.405 181.115 ;
        RECT 98.120 180.435 99.075 180.655 ;
        RECT 94.440 178.905 94.725 179.365 ;
        RECT 95.565 178.905 95.965 179.705 ;
        RECT 96.830 179.645 97.385 179.975 ;
        RECT 96.830 179.535 97.280 179.645 ;
        RECT 96.155 179.365 97.280 179.535 ;
        RECT 97.555 179.475 97.835 180.145 ;
        RECT 98.005 179.705 98.695 180.265 ;
        RECT 98.865 179.535 99.075 180.435 ;
        RECT 96.155 178.905 96.435 179.365 ;
        RECT 97.450 178.905 97.835 179.475 ;
        RECT 98.120 179.365 99.075 179.535 ;
        RECT 99.245 180.265 99.645 181.115 ;
        RECT 99.835 180.655 100.115 181.115 ;
        RECT 99.835 180.435 100.960 180.655 ;
        RECT 99.245 179.705 100.340 180.265 ;
        RECT 100.510 179.975 100.960 180.435 ;
        RECT 101.130 180.145 101.515 181.115 ;
        RECT 98.120 178.905 98.405 179.365 ;
        RECT 99.245 178.905 99.645 179.705 ;
        RECT 100.510 179.645 101.065 179.975 ;
        RECT 100.510 179.535 100.960 179.645 ;
        RECT 99.835 179.365 100.960 179.535 ;
        RECT 101.235 179.475 101.515 180.145 ;
        RECT 99.835 178.905 100.115 179.365 ;
        RECT 101.130 178.905 101.515 179.475 ;
        RECT 102.145 180.210 102.415 181.115 ;
        RECT 103.095 180.355 103.265 181.115 ;
        RECT 102.145 179.410 102.315 180.210 ;
        RECT 102.600 180.185 103.265 180.355 ;
        RECT 102.600 180.040 102.770 180.185 ;
        RECT 102.485 179.710 102.770 180.040 ;
        RECT 103.985 180.145 104.325 181.115 ;
        RECT 105.830 180.315 106.160 181.115 ;
        RECT 106.960 180.315 107.290 181.115 ;
        RECT 108.755 180.945 110.785 181.115 ;
        RECT 104.855 180.145 107.290 180.315 ;
        RECT 107.665 180.525 108.180 180.935 ;
        RECT 102.600 179.455 102.770 179.710 ;
        RECT 103.005 179.635 103.335 180.005 ;
        RECT 103.985 179.535 104.160 180.145 ;
        RECT 104.855 179.895 105.025 180.145 ;
        RECT 104.330 179.725 105.025 179.895 ;
        RECT 105.200 179.725 105.620 179.925 ;
        RECT 105.790 179.725 106.120 179.925 ;
        RECT 106.290 179.725 106.620 179.925 ;
        RECT 102.145 178.905 102.405 179.410 ;
        RECT 102.600 179.285 103.265 179.455 ;
        RECT 103.095 178.905 103.265 179.285 ;
        RECT 103.985 178.905 104.325 179.535 ;
        RECT 104.935 179.385 106.160 179.555 ;
        RECT 104.935 178.905 105.265 179.385 ;
        RECT 105.830 178.905 106.160 179.385 ;
        RECT 106.790 179.515 106.960 180.145 ;
        RECT 107.145 179.725 107.495 179.975 ;
        RECT 107.665 179.715 108.005 180.525 ;
        RECT 108.755 180.280 108.925 180.945 ;
        RECT 109.320 180.605 110.445 180.775 ;
        RECT 108.175 180.090 108.925 180.280 ;
        RECT 109.095 180.265 110.105 180.435 ;
        RECT 107.665 179.545 108.895 179.715 ;
        RECT 106.790 178.905 107.290 179.515 ;
        RECT 107.940 178.940 108.185 179.545 ;
        RECT 109.095 178.905 109.285 180.265 ;
        RECT 109.455 179.245 109.730 180.065 ;
        RECT 109.935 179.465 110.105 180.265 ;
        RECT 110.275 179.475 110.445 180.605 ;
        RECT 110.615 179.975 110.785 180.945 ;
        RECT 111.295 180.145 111.630 181.115 ;
        RECT 110.615 179.645 110.810 179.975 ;
        RECT 111.035 179.645 111.290 179.975 ;
        RECT 111.035 179.475 111.205 179.645 ;
        RECT 111.460 179.475 111.630 180.145 ;
        RECT 110.275 179.305 111.205 179.475 ;
        RECT 110.275 179.270 110.450 179.305 ;
        RECT 109.455 179.075 109.735 179.245 ;
        RECT 109.455 178.905 109.730 179.075 ;
        RECT 109.920 178.905 110.450 179.270 ;
        RECT 111.375 178.905 111.630 179.475 ;
        RECT 111.810 180.095 112.065 180.975 ;
        RECT 113.390 180.735 113.560 181.025 ;
        RECT 112.760 180.565 113.560 180.735 ;
        RECT 114.150 180.775 115.020 181.115 ;
        RECT 111.810 179.445 112.020 180.095 ;
        RECT 112.760 179.975 112.930 180.565 ;
        RECT 114.150 180.395 114.320 180.775 ;
        RECT 115.255 180.655 115.425 181.115 ;
        RECT 116.260 180.685 116.430 181.025 ;
        RECT 117.165 180.685 117.335 181.025 ;
        RECT 113.100 180.225 114.320 180.395 ;
        RECT 114.490 180.315 114.950 180.605 ;
        RECT 115.255 180.485 115.815 180.655 ;
        RECT 116.260 180.515 117.335 180.685 ;
        RECT 117.505 180.785 118.185 181.115 ;
        RECT 118.400 180.785 118.650 181.115 ;
        RECT 115.645 180.345 115.815 180.485 ;
        RECT 114.490 180.305 115.455 180.315 ;
        RECT 114.150 180.135 114.320 180.225 ;
        RECT 114.780 180.145 115.455 180.305 ;
        RECT 112.190 179.945 112.930 179.975 ;
        RECT 112.190 179.645 113.105 179.945 ;
        RECT 112.780 179.470 113.105 179.645 ;
        RECT 111.810 178.915 112.065 179.445 ;
        RECT 112.785 179.115 113.105 179.470 ;
        RECT 113.275 179.685 113.815 180.055 ;
        RECT 114.150 179.965 114.555 180.135 ;
        RECT 113.275 179.285 113.515 179.685 ;
        RECT 113.995 179.515 114.215 179.795 ;
        RECT 113.685 179.345 114.215 179.515 ;
        RECT 113.685 179.115 113.855 179.345 ;
        RECT 112.785 178.945 113.855 179.115 ;
        RECT 114.385 179.185 114.555 179.965 ;
        RECT 114.725 179.355 115.075 179.975 ;
        RECT 115.245 179.355 115.455 180.145 ;
        RECT 115.645 180.175 117.145 180.345 ;
        RECT 115.645 179.485 115.815 180.175 ;
        RECT 117.505 180.005 117.675 180.785 ;
        RECT 118.480 180.655 118.650 180.785 ;
        RECT 115.985 179.835 117.675 180.005 ;
        RECT 117.845 180.225 118.310 180.615 ;
        RECT 118.480 180.485 118.875 180.655 ;
        RECT 115.985 179.655 116.155 179.835 ;
        RECT 114.385 178.905 115.335 179.185 ;
        RECT 115.645 179.095 115.905 179.485 ;
        RECT 116.325 179.415 117.115 179.665 ;
        RECT 115.555 178.925 115.905 179.095 ;
        RECT 117.320 179.125 117.490 179.835 ;
        RECT 117.845 179.635 118.015 180.225 ;
        RECT 117.660 179.415 118.015 179.635 ;
        RECT 118.185 179.415 118.535 180.035 ;
        RECT 118.705 179.125 118.875 180.485 ;
        RECT 119.240 180.315 119.565 181.100 ;
        RECT 119.045 179.265 119.505 180.315 ;
        RECT 117.320 178.955 118.175 179.125 ;
        RECT 118.380 178.955 118.875 179.125 ;
        RECT 119.735 178.995 119.905 181.115 ;
        RECT 120.575 180.615 120.830 181.115 ;
        RECT 120.080 180.445 120.830 180.615 ;
        RECT 120.080 179.455 120.310 180.445 ;
        RECT 120.480 179.625 120.830 180.275 ;
        RECT 121.005 180.210 121.275 181.115 ;
        RECT 121.955 180.355 122.125 181.115 ;
        RECT 120.080 179.285 120.830 179.455 ;
        RECT 120.575 178.995 120.830 179.285 ;
        RECT 121.005 179.410 121.175 180.210 ;
        RECT 121.460 180.185 122.125 180.355 ;
        RECT 122.475 180.355 122.645 181.115 ;
        RECT 122.475 180.185 123.140 180.355 ;
        RECT 123.325 180.210 123.595 181.115 ;
        RECT 121.460 180.040 121.630 180.185 ;
        RECT 121.345 179.710 121.630 180.040 ;
        RECT 122.970 180.040 123.140 180.185 ;
        RECT 121.460 179.455 121.630 179.710 ;
        RECT 121.865 179.635 122.195 180.005 ;
        RECT 122.405 179.635 122.735 180.005 ;
        RECT 122.970 179.710 123.255 180.040 ;
        RECT 122.970 179.455 123.140 179.710 ;
        RECT 121.005 178.905 121.265 179.410 ;
        RECT 121.460 179.285 122.125 179.455 ;
        RECT 121.955 178.905 122.125 179.285 ;
        RECT 122.475 179.285 123.140 179.455 ;
        RECT 123.425 179.410 123.595 180.210 ;
        RECT 122.475 178.905 122.645 179.285 ;
        RECT 123.335 178.905 123.595 179.410 ;
        RECT 25.765 177.765 26.095 178.395 ;
        RECT 26.705 177.890 26.965 178.395 ;
        RECT 27.655 178.015 27.825 178.395 ;
        RECT 25.765 177.165 26.015 177.765 ;
        RECT 26.185 177.325 26.515 177.575 ;
        RECT 25.765 176.185 26.095 177.165 ;
        RECT 26.705 177.090 26.875 177.890 ;
        RECT 27.160 177.845 27.825 178.015 ;
        RECT 28.090 177.855 28.345 178.385 ;
        RECT 29.065 178.185 30.135 178.355 ;
        RECT 27.160 177.590 27.330 177.845 ;
        RECT 27.045 177.260 27.330 177.590 ;
        RECT 27.565 177.295 27.895 177.665 ;
        RECT 27.160 177.115 27.330 177.260 ;
        RECT 28.090 177.205 28.300 177.855 ;
        RECT 29.065 177.830 29.385 178.185 ;
        RECT 29.060 177.655 29.385 177.830 ;
        RECT 28.470 177.355 29.385 177.655 ;
        RECT 29.555 177.615 29.795 178.015 ;
        RECT 29.965 177.955 30.135 178.185 ;
        RECT 30.665 178.115 31.615 178.395 ;
        RECT 31.835 178.205 32.185 178.375 ;
        RECT 29.965 177.785 30.495 177.955 ;
        RECT 28.470 177.325 29.210 177.355 ;
        RECT 26.705 176.185 26.975 177.090 ;
        RECT 27.160 176.945 27.825 177.115 ;
        RECT 27.655 176.185 27.825 176.945 ;
        RECT 28.090 176.325 28.345 177.205 ;
        RECT 29.040 176.735 29.210 177.325 ;
        RECT 29.555 177.245 30.095 177.615 ;
        RECT 30.275 177.505 30.495 177.785 ;
        RECT 30.665 177.335 30.835 178.115 ;
        RECT 30.430 177.165 30.835 177.335 ;
        RECT 31.005 177.325 31.355 177.945 ;
        RECT 30.430 177.075 30.600 177.165 ;
        RECT 31.525 177.155 31.735 177.945 ;
        RECT 29.380 176.905 30.600 177.075 ;
        RECT 31.060 176.995 31.735 177.155 ;
        RECT 29.040 176.565 29.840 176.735 ;
        RECT 29.670 176.275 29.840 176.565 ;
        RECT 30.430 176.525 30.600 176.905 ;
        RECT 30.770 176.985 31.735 176.995 ;
        RECT 31.925 177.815 32.185 178.205 ;
        RECT 33.600 178.175 34.455 178.345 ;
        RECT 34.660 178.175 35.155 178.345 ;
        RECT 31.925 177.125 32.095 177.815 ;
        RECT 32.265 177.465 32.435 177.645 ;
        RECT 32.605 177.635 33.395 177.885 ;
        RECT 33.600 177.465 33.770 178.175 ;
        RECT 33.940 177.665 34.295 177.885 ;
        RECT 32.265 177.295 33.955 177.465 ;
        RECT 30.770 176.695 31.230 176.985 ;
        RECT 31.925 176.955 33.425 177.125 ;
        RECT 31.925 176.815 32.095 176.955 ;
        RECT 31.535 176.645 32.095 176.815 ;
        RECT 30.430 176.185 31.300 176.525 ;
        RECT 31.535 176.185 31.705 176.645 ;
        RECT 32.540 176.615 33.615 176.785 ;
        RECT 32.540 176.275 32.710 176.615 ;
        RECT 33.445 176.275 33.615 176.615 ;
        RECT 33.785 176.515 33.955 177.295 ;
        RECT 34.125 177.075 34.295 177.665 ;
        RECT 34.465 177.265 34.815 177.885 ;
        RECT 34.125 176.685 34.590 177.075 ;
        RECT 34.985 176.815 35.155 178.175 ;
        RECT 35.325 176.985 35.785 178.035 ;
        RECT 34.760 176.645 35.155 176.815 ;
        RECT 34.760 176.515 34.930 176.645 ;
        RECT 33.785 176.185 34.465 176.515 ;
        RECT 34.680 176.185 34.930 176.515 ;
        RECT 35.520 176.200 35.845 176.985 ;
        RECT 36.015 176.185 36.185 178.305 ;
        RECT 36.855 178.015 37.110 178.305 ;
        RECT 36.360 177.845 37.110 178.015 ;
        RECT 36.360 176.855 36.590 177.845 ;
        RECT 37.750 177.825 38.005 178.395 ;
        RECT 38.930 178.030 39.460 178.395 ;
        RECT 39.650 178.225 39.925 178.395 ;
        RECT 39.645 178.055 39.925 178.225 ;
        RECT 38.930 177.995 39.105 178.030 ;
        RECT 38.175 177.825 39.105 177.995 ;
        RECT 36.760 177.025 37.110 177.675 ;
        RECT 37.750 177.155 37.920 177.825 ;
        RECT 38.175 177.655 38.345 177.825 ;
        RECT 38.090 177.325 38.345 177.655 ;
        RECT 38.570 177.325 38.765 177.655 ;
        RECT 36.360 176.685 37.110 176.855 ;
        RECT 36.855 176.185 37.110 176.685 ;
        RECT 37.750 176.185 38.085 177.155 ;
        RECT 38.595 176.355 38.765 177.325 ;
        RECT 38.935 176.695 39.105 177.825 ;
        RECT 39.275 177.035 39.445 177.835 ;
        RECT 39.650 177.235 39.925 178.055 ;
        RECT 40.095 177.035 40.285 178.395 ;
        RECT 41.195 177.755 41.440 178.360 ;
        RECT 43.930 177.785 44.430 178.395 ;
        RECT 40.485 177.585 41.715 177.755 ;
        RECT 39.275 176.865 40.285 177.035 ;
        RECT 40.455 177.020 41.205 177.210 ;
        RECT 38.935 176.525 40.060 176.695 ;
        RECT 40.455 176.355 40.625 177.020 ;
        RECT 41.375 176.775 41.715 177.585 ;
        RECT 43.725 177.325 44.075 177.575 ;
        RECT 44.260 177.155 44.430 177.785 ;
        RECT 45.060 177.915 45.390 178.395 ;
        RECT 45.955 177.915 46.285 178.395 ;
        RECT 45.060 177.745 46.285 177.915 ;
        RECT 46.895 177.765 47.235 178.395 ;
        RECT 44.600 177.375 44.930 177.575 ;
        RECT 45.100 177.375 45.430 177.575 ;
        RECT 45.600 177.375 46.020 177.575 ;
        RECT 46.195 177.405 46.890 177.575 ;
        RECT 46.195 177.155 46.365 177.405 ;
        RECT 47.060 177.155 47.235 177.765 ;
        RECT 41.200 176.365 41.715 176.775 ;
        RECT 43.930 176.985 46.365 177.155 ;
        RECT 38.595 176.185 40.625 176.355 ;
        RECT 43.930 176.185 44.260 176.985 ;
        RECT 45.060 176.185 45.390 176.985 ;
        RECT 46.895 176.185 47.235 177.155 ;
        RECT 47.865 177.765 48.205 178.395 ;
        RECT 48.815 177.915 49.145 178.395 ;
        RECT 49.710 177.915 50.040 178.395 ;
        RECT 47.865 177.155 48.040 177.765 ;
        RECT 48.815 177.745 50.040 177.915 ;
        RECT 50.670 177.785 51.170 178.395 ;
        RECT 48.210 177.405 48.905 177.575 ;
        RECT 48.735 177.155 48.905 177.405 ;
        RECT 49.080 177.375 49.500 177.575 ;
        RECT 49.670 177.375 50.000 177.575 ;
        RECT 50.170 177.375 50.500 177.575 ;
        RECT 50.670 177.155 50.840 177.785 ;
        RECT 51.545 177.765 51.885 178.395 ;
        RECT 52.495 177.915 52.825 178.395 ;
        RECT 53.390 177.915 53.720 178.395 ;
        RECT 51.025 177.325 51.375 177.575 ;
        RECT 51.545 177.155 51.720 177.765 ;
        RECT 52.495 177.745 53.720 177.915 ;
        RECT 54.350 177.785 54.850 178.395 ;
        RECT 51.890 177.405 52.585 177.575 ;
        RECT 52.415 177.155 52.585 177.405 ;
        RECT 52.760 177.375 53.180 177.575 ;
        RECT 53.350 177.375 53.680 177.575 ;
        RECT 53.850 177.375 54.180 177.575 ;
        RECT 54.350 177.155 54.520 177.785 ;
        RECT 55.960 177.755 56.205 178.360 ;
        RECT 55.685 177.585 56.915 177.755 ;
        RECT 54.705 177.325 55.055 177.575 ;
        RECT 47.865 176.185 48.205 177.155 ;
        RECT 48.735 176.985 51.170 177.155 ;
        RECT 49.710 176.185 50.040 176.985 ;
        RECT 50.840 176.185 51.170 176.985 ;
        RECT 51.545 176.185 51.885 177.155 ;
        RECT 52.415 176.985 54.850 177.155 ;
        RECT 53.390 176.185 53.720 176.985 ;
        RECT 54.520 176.185 54.850 176.985 ;
        RECT 55.685 176.775 56.025 177.585 ;
        RECT 56.195 177.020 56.945 177.210 ;
        RECT 55.685 176.365 56.200 176.775 ;
        RECT 56.775 176.355 56.945 177.020 ;
        RECT 57.115 177.035 57.305 178.395 ;
        RECT 57.475 177.545 57.750 178.395 ;
        RECT 57.940 178.030 58.470 178.395 ;
        RECT 58.295 177.995 58.470 178.030 ;
        RECT 57.475 177.375 57.755 177.545 ;
        RECT 57.475 177.235 57.750 177.375 ;
        RECT 57.955 177.035 58.125 177.835 ;
        RECT 57.115 176.865 58.125 177.035 ;
        RECT 58.295 177.825 59.225 177.995 ;
        RECT 59.395 177.825 59.650 178.395 ;
        RECT 60.795 177.915 61.055 178.305 ;
        RECT 61.655 177.915 61.950 178.305 ;
        RECT 62.575 178.065 62.875 178.395 ;
        RECT 58.295 176.695 58.465 177.825 ;
        RECT 59.055 177.655 59.225 177.825 ;
        RECT 57.340 176.525 58.465 176.695 ;
        RECT 58.635 177.325 58.830 177.655 ;
        RECT 59.055 177.325 59.310 177.655 ;
        RECT 58.635 176.355 58.805 177.325 ;
        RECT 59.480 177.155 59.650 177.825 ;
        RECT 56.775 176.185 58.805 176.355 ;
        RECT 59.315 176.185 59.650 177.155 ;
        RECT 60.300 177.745 61.950 177.915 ;
        RECT 60.300 177.235 60.705 177.745 ;
        RECT 60.875 177.405 62.015 177.575 ;
        RECT 60.300 177.065 61.055 177.235 ;
        RECT 60.795 176.815 61.055 177.065 ;
        RECT 61.845 177.155 62.015 177.405 ;
        RECT 62.185 177.325 62.535 177.895 ;
        RECT 62.705 177.155 62.875 178.065 ;
        RECT 61.845 176.985 62.875 177.155 ;
        RECT 60.795 176.645 61.915 176.815 ;
        RECT 60.795 176.185 61.055 176.645 ;
        RECT 61.655 176.185 61.915 176.645 ;
        RECT 62.565 176.185 62.875 176.985 ;
        RECT 64.405 177.820 64.660 178.395 ;
        RECT 65.375 178.015 65.545 178.395 ;
        RECT 64.830 177.845 65.545 178.015 ;
        RECT 64.405 177.090 64.575 177.820 ;
        RECT 64.830 177.655 65.000 177.845 ;
        RECT 66.245 177.820 66.500 178.395 ;
        RECT 67.215 178.015 67.385 178.395 ;
        RECT 66.670 177.845 67.385 178.015 ;
        RECT 68.115 178.035 68.445 178.395 ;
        RECT 69.145 178.035 69.475 178.395 ;
        RECT 64.745 177.325 65.000 177.655 ;
        RECT 64.830 177.115 65.000 177.325 ;
        RECT 65.280 177.295 65.635 177.665 ;
        RECT 64.405 176.185 64.660 177.090 ;
        RECT 64.830 176.945 65.545 177.115 ;
        RECT 65.375 176.185 65.545 176.945 ;
        RECT 66.245 177.090 66.415 177.820 ;
        RECT 66.670 177.655 66.840 177.845 ;
        RECT 68.115 177.825 69.475 178.035 ;
        RECT 69.985 177.805 70.695 178.395 ;
        RECT 71.635 177.995 71.835 178.350 ;
        RECT 72.505 177.995 72.705 178.340 ;
        RECT 70.465 177.715 70.695 177.805 ;
        RECT 66.585 177.325 66.840 177.655 ;
        RECT 66.670 177.115 66.840 177.325 ;
        RECT 67.120 177.295 67.475 177.665 ;
        RECT 68.105 177.325 68.415 177.655 ;
        RECT 68.625 177.325 69.000 177.655 ;
        RECT 69.320 177.325 69.815 177.655 ;
        RECT 66.245 176.185 66.500 177.090 ;
        RECT 66.670 176.945 67.385 177.115 ;
        RECT 67.215 176.185 67.385 176.945 ;
        RECT 68.625 176.355 68.795 177.325 ;
        RECT 68.965 176.835 69.295 177.055 ;
        RECT 69.490 177.035 69.815 177.325 ;
        RECT 69.990 177.035 70.320 177.575 ;
        RECT 70.490 176.835 70.695 177.715 ;
        RECT 68.965 176.605 70.695 176.835 ;
        RECT 68.965 176.205 69.295 176.605 ;
        RECT 69.995 176.185 70.695 176.605 ;
        RECT 70.865 177.825 72.705 177.995 ;
        RECT 73.440 177.995 73.610 178.245 ;
        RECT 73.440 177.825 73.915 177.995 ;
        RECT 70.865 176.200 71.125 177.825 ;
        RECT 71.305 176.855 71.525 177.655 ;
        RECT 71.765 177.035 72.065 177.655 ;
        RECT 72.235 177.035 72.565 177.655 ;
        RECT 72.735 177.035 73.055 177.655 ;
        RECT 73.225 177.035 73.575 177.655 ;
        RECT 73.745 176.855 73.915 177.825 ;
        RECT 74.290 177.785 74.790 178.395 ;
        RECT 74.085 177.325 74.435 177.575 ;
        RECT 74.620 177.155 74.790 177.785 ;
        RECT 75.420 177.915 75.750 178.395 ;
        RECT 76.315 177.915 76.645 178.395 ;
        RECT 75.420 177.745 76.645 177.915 ;
        RECT 77.255 177.765 77.595 178.395 ;
        RECT 82.495 178.390 82.665 178.395 ;
        RECT 83.335 178.390 83.505 178.395 ;
        RECT 84.175 178.390 84.425 178.395 ;
        RECT 78.215 177.915 78.545 178.390 ;
        RECT 79.055 177.915 79.385 178.390 ;
        RECT 79.895 177.915 80.225 178.390 ;
        RECT 80.735 177.915 81.065 178.390 ;
        RECT 81.575 177.915 81.905 178.390 ;
        RECT 82.415 177.915 82.745 178.390 ;
        RECT 83.255 177.915 83.585 178.390 ;
        RECT 84.095 177.915 84.425 178.390 ;
        RECT 84.935 177.915 85.265 178.390 ;
        RECT 85.775 177.915 86.105 178.390 ;
        RECT 86.615 177.915 86.945 178.390 ;
        RECT 87.455 177.915 87.785 178.390 ;
        RECT 88.295 177.915 88.625 178.390 ;
        RECT 74.960 177.375 75.290 177.575 ;
        RECT 75.460 177.375 75.790 177.575 ;
        RECT 75.960 177.375 76.380 177.575 ;
        RECT 76.555 177.405 77.250 177.575 ;
        RECT 76.555 177.155 76.725 177.405 ;
        RECT 77.420 177.155 77.595 177.765 ;
        RECT 71.305 176.645 73.915 176.855 ;
        RECT 74.290 176.985 76.725 177.155 ;
        RECT 74.290 176.185 74.620 176.985 ;
        RECT 75.420 176.185 75.750 176.985 ;
        RECT 77.255 176.185 77.595 177.155 ;
        RECT 77.765 177.745 84.425 177.915 ;
        RECT 84.595 177.745 86.945 177.915 ;
        RECT 87.115 177.745 88.625 177.915 ;
        RECT 96.145 177.765 96.475 178.395 ;
        RECT 98.925 177.765 99.265 178.395 ;
        RECT 99.875 177.915 100.205 178.395 ;
        RECT 100.770 177.915 101.100 178.395 ;
        RECT 77.765 177.205 78.040 177.745 ;
        RECT 84.595 177.575 84.770 177.745 ;
        RECT 87.115 177.575 87.285 177.745 ;
        RECT 78.210 177.375 84.770 177.575 ;
        RECT 84.975 177.375 87.285 177.575 ;
        RECT 87.455 177.375 88.630 177.575 ;
        RECT 84.595 177.205 84.770 177.375 ;
        RECT 87.115 177.205 87.285 177.375 ;
        RECT 77.765 177.035 84.425 177.205 ;
        RECT 84.595 177.035 86.945 177.205 ;
        RECT 87.115 177.035 88.625 177.205 ;
        RECT 78.215 176.185 78.545 177.035 ;
        RECT 79.055 176.185 79.385 177.035 ;
        RECT 79.895 176.185 80.225 177.035 ;
        RECT 80.735 176.185 81.065 177.035 ;
        RECT 81.575 176.185 81.905 177.035 ;
        RECT 82.415 176.185 82.745 177.035 ;
        RECT 83.255 176.185 83.585 177.035 ;
        RECT 84.095 176.185 84.425 177.035 ;
        RECT 84.935 176.185 85.265 177.035 ;
        RECT 85.775 176.185 86.105 177.035 ;
        RECT 86.615 176.185 86.945 177.035 ;
        RECT 87.455 176.185 87.785 177.035 ;
        RECT 88.295 176.185 88.625 177.035 ;
        RECT 96.145 177.165 96.395 177.765 ;
        RECT 96.565 177.325 96.895 177.575 ;
        RECT 96.145 176.185 96.475 177.165 ;
        RECT 98.925 177.155 99.100 177.765 ;
        RECT 99.875 177.745 101.100 177.915 ;
        RECT 101.730 177.785 102.230 178.395 ;
        RECT 99.270 177.405 99.965 177.575 ;
        RECT 100.140 177.545 100.560 177.575 ;
        RECT 99.795 177.155 99.965 177.405 ;
        RECT 100.135 177.375 100.560 177.545 ;
        RECT 100.730 177.375 101.060 177.575 ;
        RECT 101.230 177.375 101.560 177.575 ;
        RECT 101.730 177.155 101.900 177.785 ;
        RECT 105.365 177.765 105.705 178.395 ;
        RECT 106.315 177.915 106.645 178.395 ;
        RECT 107.210 177.915 107.540 178.395 ;
        RECT 102.085 177.325 102.435 177.575 ;
        RECT 105.365 177.155 105.540 177.765 ;
        RECT 106.315 177.745 107.540 177.915 ;
        RECT 108.170 177.785 108.670 178.395 ;
        RECT 109.045 177.825 109.430 178.395 ;
        RECT 110.445 177.935 110.725 178.395 ;
        RECT 105.710 177.405 106.405 177.575 ;
        RECT 106.235 177.155 106.405 177.405 ;
        RECT 106.580 177.375 107.000 177.575 ;
        RECT 107.170 177.375 107.500 177.575 ;
        RECT 107.670 177.375 108.000 177.575 ;
        RECT 108.170 177.155 108.340 177.785 ;
        RECT 108.525 177.325 108.875 177.575 ;
        RECT 109.045 177.155 109.325 177.825 ;
        RECT 109.600 177.765 110.725 177.935 ;
        RECT 109.600 177.655 110.050 177.765 ;
        RECT 109.495 177.325 110.050 177.655 ;
        RECT 110.915 177.595 111.315 178.395 ;
        RECT 112.155 177.935 112.440 178.395 ;
        RECT 98.925 176.185 99.265 177.155 ;
        RECT 99.795 176.985 102.230 177.155 ;
        RECT 100.770 176.185 101.100 176.985 ;
        RECT 101.900 176.185 102.230 176.985 ;
        RECT 105.365 176.185 105.705 177.155 ;
        RECT 106.235 176.985 108.670 177.155 ;
        RECT 107.210 176.185 107.540 176.985 ;
        RECT 108.340 176.185 108.670 176.985 ;
        RECT 109.045 176.185 109.430 177.155 ;
        RECT 109.600 176.865 110.050 177.325 ;
        RECT 110.220 177.035 111.315 177.595 ;
        RECT 109.600 176.645 110.725 176.865 ;
        RECT 110.445 176.185 110.725 176.645 ;
        RECT 110.915 176.185 111.315 177.035 ;
        RECT 111.485 177.765 112.440 177.935 ;
        RECT 113.625 177.765 113.955 178.395 ;
        RECT 117.305 177.765 117.635 178.395 ;
        RECT 111.485 176.865 111.695 177.765 ;
        RECT 111.865 177.035 112.555 177.595 ;
        RECT 113.205 177.325 113.535 177.575 ;
        RECT 113.705 177.165 113.955 177.765 ;
        RECT 116.885 177.325 117.215 177.575 ;
        RECT 117.385 177.165 117.635 177.765 ;
        RECT 111.485 176.645 112.440 176.865 ;
        RECT 112.155 176.185 112.440 176.645 ;
        RECT 113.625 176.185 113.955 177.165 ;
        RECT 117.305 176.185 117.635 177.165 ;
        RECT 26.225 174.695 26.555 175.675 ;
        RECT 27.280 175.215 27.565 175.675 ;
        RECT 27.280 174.995 28.235 175.215 ;
        RECT 26.225 174.095 26.475 174.695 ;
        RECT 26.645 174.285 26.975 174.535 ;
        RECT 27.165 174.265 27.855 174.825 ;
        RECT 28.025 174.095 28.235 174.995 ;
        RECT 26.225 173.465 26.555 174.095 ;
        RECT 27.280 173.925 28.235 174.095 ;
        RECT 28.405 174.825 28.805 175.675 ;
        RECT 28.995 175.215 29.275 175.675 ;
        RECT 28.995 174.995 30.120 175.215 ;
        RECT 28.405 174.265 29.500 174.825 ;
        RECT 29.670 174.535 30.120 174.995 ;
        RECT 30.290 174.705 30.675 175.675 ;
        RECT 27.280 173.465 27.565 173.925 ;
        RECT 28.405 173.465 28.805 174.265 ;
        RECT 29.670 174.205 30.225 174.535 ;
        RECT 29.670 174.095 30.120 174.205 ;
        RECT 28.995 173.925 30.120 174.095 ;
        RECT 30.395 174.035 30.675 174.705 ;
        RECT 28.995 173.465 29.275 173.925 ;
        RECT 30.290 173.465 30.675 174.035 ;
        RECT 31.310 174.705 31.645 175.675 ;
        RECT 32.155 175.505 34.185 175.675 ;
        RECT 31.310 174.035 31.480 174.705 ;
        RECT 32.155 174.535 32.325 175.505 ;
        RECT 31.650 174.205 31.905 174.535 ;
        RECT 32.130 174.205 32.325 174.535 ;
        RECT 32.495 175.165 33.620 175.335 ;
        RECT 31.735 174.035 31.905 174.205 ;
        RECT 32.495 174.035 32.665 175.165 ;
        RECT 31.310 173.465 31.565 174.035 ;
        RECT 31.735 173.865 32.665 174.035 ;
        RECT 32.835 174.825 33.845 174.995 ;
        RECT 32.835 174.025 33.005 174.825 ;
        RECT 33.210 174.485 33.485 174.625 ;
        RECT 33.205 174.315 33.485 174.485 ;
        RECT 32.490 173.830 32.665 173.865 ;
        RECT 32.490 173.465 33.020 173.830 ;
        RECT 33.210 173.465 33.485 174.315 ;
        RECT 33.655 173.465 33.845 174.825 ;
        RECT 34.015 174.840 34.185 175.505 ;
        RECT 34.760 175.085 35.275 175.495 ;
        RECT 34.015 174.650 34.765 174.840 ;
        RECT 34.935 174.275 35.275 175.085 ;
        RECT 35.650 174.875 35.980 175.675 ;
        RECT 36.780 174.875 37.110 175.675 ;
        RECT 35.650 174.705 38.085 174.875 ;
        RECT 38.615 174.705 38.955 175.675 ;
        RECT 35.445 174.285 35.795 174.535 ;
        RECT 34.045 174.105 35.275 174.275 ;
        RECT 34.755 173.500 35.000 174.105 ;
        RECT 35.980 174.075 36.150 174.705 ;
        RECT 36.320 174.285 36.650 174.485 ;
        RECT 36.820 174.285 37.150 174.485 ;
        RECT 37.320 174.285 37.740 174.485 ;
        RECT 37.915 174.455 38.085 174.705 ;
        RECT 37.915 174.285 38.610 174.455 ;
        RECT 35.650 173.465 36.150 174.075 ;
        RECT 36.780 173.945 38.005 174.115 ;
        RECT 38.780 174.095 38.955 174.705 ;
        RECT 36.780 173.465 37.110 173.945 ;
        RECT 37.675 173.465 38.005 173.945 ;
        RECT 38.615 173.465 38.955 174.095 ;
        RECT 39.125 174.705 39.465 175.675 ;
        RECT 40.970 174.875 41.300 175.675 ;
        RECT 42.100 174.875 42.430 175.675 ;
        RECT 39.995 174.705 42.430 174.875 ;
        RECT 43.010 174.875 43.340 175.675 ;
        RECT 44.140 174.875 44.470 175.675 ;
        RECT 43.010 174.705 45.445 174.875 ;
        RECT 45.975 174.705 46.315 175.675 ;
        RECT 39.125 174.145 39.300 174.705 ;
        RECT 39.995 174.455 40.165 174.705 ;
        RECT 39.470 174.285 40.165 174.455 ;
        RECT 40.340 174.285 40.760 174.485 ;
        RECT 40.930 174.285 41.260 174.485 ;
        RECT 41.430 174.285 41.760 174.485 ;
        RECT 39.125 174.095 39.355 174.145 ;
        RECT 39.125 173.465 39.465 174.095 ;
        RECT 40.075 173.945 41.300 174.115 ;
        RECT 40.075 173.465 40.405 173.945 ;
        RECT 40.970 173.465 41.300 173.945 ;
        RECT 41.930 174.075 42.100 174.705 ;
        RECT 42.285 174.285 42.635 174.535 ;
        RECT 42.805 174.285 43.155 174.535 ;
        RECT 43.340 174.075 43.510 174.705 ;
        RECT 43.680 174.285 44.010 174.485 ;
        RECT 44.180 174.285 44.510 174.485 ;
        RECT 44.680 174.285 45.100 174.485 ;
        RECT 45.275 174.455 45.445 174.705 ;
        RECT 45.275 174.285 45.970 174.455 ;
        RECT 46.140 174.145 46.315 174.705 ;
        RECT 41.930 173.465 42.430 174.075 ;
        RECT 43.010 173.465 43.510 174.075 ;
        RECT 44.140 173.945 45.365 174.115 ;
        RECT 46.085 174.095 46.315 174.145 ;
        RECT 44.140 173.465 44.470 173.945 ;
        RECT 45.035 173.465 45.365 173.945 ;
        RECT 45.975 173.465 46.315 174.095 ;
        RECT 46.485 174.705 46.825 175.675 ;
        RECT 48.330 174.875 48.660 175.675 ;
        RECT 49.460 174.875 49.790 175.675 ;
        RECT 52.120 175.215 52.405 175.675 ;
        RECT 52.120 174.995 53.075 175.215 ;
        RECT 47.355 174.705 49.790 174.875 ;
        RECT 46.485 174.145 46.660 174.705 ;
        RECT 47.355 174.455 47.525 174.705 ;
        RECT 46.830 174.285 47.525 174.455 ;
        RECT 47.700 174.285 48.120 174.485 ;
        RECT 48.290 174.285 48.620 174.485 ;
        RECT 48.790 174.285 49.120 174.485 ;
        RECT 46.485 174.095 46.715 174.145 ;
        RECT 46.485 173.465 46.825 174.095 ;
        RECT 47.435 173.945 48.660 174.115 ;
        RECT 47.435 173.465 47.765 173.945 ;
        RECT 48.330 173.465 48.660 173.945 ;
        RECT 49.290 174.075 49.460 174.705 ;
        RECT 49.645 174.285 49.995 174.535 ;
        RECT 52.005 174.265 52.695 174.825 ;
        RECT 52.865 174.095 53.075 174.995 ;
        RECT 49.290 173.465 49.790 174.075 ;
        RECT 52.120 173.925 53.075 174.095 ;
        RECT 53.245 174.825 53.645 175.675 ;
        RECT 53.835 175.215 54.115 175.675 ;
        RECT 53.835 174.995 54.960 175.215 ;
        RECT 53.245 174.265 54.340 174.825 ;
        RECT 54.510 174.535 54.960 174.995 ;
        RECT 55.130 174.705 55.515 175.675 ;
        RECT 57.695 175.505 59.725 175.675 ;
        RECT 52.120 173.465 52.405 173.925 ;
        RECT 53.245 173.465 53.645 174.265 ;
        RECT 54.510 174.205 55.065 174.535 ;
        RECT 54.510 174.095 54.960 174.205 ;
        RECT 53.835 173.925 54.960 174.095 ;
        RECT 55.235 174.035 55.515 174.705 ;
        RECT 56.605 175.085 57.120 175.495 ;
        RECT 56.605 174.275 56.945 175.085 ;
        RECT 57.695 174.840 57.865 175.505 ;
        RECT 58.260 175.165 59.385 175.335 ;
        RECT 57.115 174.650 57.865 174.840 ;
        RECT 58.035 174.825 59.045 174.995 ;
        RECT 56.605 174.105 57.835 174.275 ;
        RECT 53.835 173.465 54.115 173.925 ;
        RECT 55.130 173.465 55.515 174.035 ;
        RECT 56.880 173.500 57.125 174.105 ;
        RECT 58.035 173.465 58.225 174.825 ;
        RECT 58.395 174.145 58.670 174.625 ;
        RECT 58.395 173.975 58.675 174.145 ;
        RECT 58.875 174.025 59.045 174.825 ;
        RECT 59.215 174.035 59.385 175.165 ;
        RECT 59.555 174.535 59.725 175.505 ;
        RECT 60.235 174.705 60.570 175.675 ;
        RECT 59.555 174.205 59.750 174.535 ;
        RECT 59.975 174.205 60.230 174.535 ;
        RECT 59.975 174.035 60.145 174.205 ;
        RECT 60.400 174.035 60.570 174.705 ;
        RECT 58.395 173.465 58.670 173.975 ;
        RECT 59.215 173.865 60.145 174.035 ;
        RECT 59.215 173.830 59.390 173.865 ;
        RECT 58.860 173.465 59.390 173.830 ;
        RECT 60.315 173.465 60.570 174.035 ;
        RECT 62.585 174.770 62.855 175.675 ;
        RECT 63.535 174.915 63.705 175.675 ;
        RECT 62.585 173.970 62.755 174.770 ;
        RECT 63.040 174.745 63.705 174.915 ;
        RECT 68.115 174.865 68.445 175.675 ;
        RECT 63.040 174.600 63.210 174.745 ;
        RECT 68.115 174.695 68.830 174.865 ;
        RECT 62.925 174.270 63.210 174.600 ;
        RECT 63.040 174.015 63.210 174.270 ;
        RECT 63.445 174.195 63.775 174.565 ;
        RECT 68.110 174.285 68.490 174.525 ;
        RECT 68.660 174.455 68.830 174.695 ;
        RECT 69.035 174.825 69.205 175.675 ;
        RECT 69.875 174.825 70.045 175.675 ;
        RECT 69.035 174.655 70.045 174.825 ;
        RECT 68.660 174.285 69.160 174.455 ;
        RECT 68.660 174.115 68.830 174.285 ;
        RECT 69.550 174.115 70.045 174.655 ;
        RECT 62.585 173.465 62.845 173.970 ;
        RECT 63.040 173.845 63.705 174.015 ;
        RECT 63.535 173.465 63.705 173.845 ;
        RECT 68.195 173.945 68.830 174.115 ;
        RECT 69.035 173.945 70.045 174.115 ;
        RECT 68.195 173.465 68.365 173.945 ;
        RECT 69.035 173.465 69.205 173.945 ;
        RECT 69.875 173.465 70.045 173.945 ;
        RECT 71.765 174.770 72.020 175.675 ;
        RECT 72.735 174.915 72.905 175.675 ;
        RECT 71.765 174.040 71.935 174.770 ;
        RECT 72.190 174.745 72.905 174.915 ;
        RECT 73.255 174.915 73.425 175.675 ;
        RECT 73.255 174.745 73.970 174.915 ;
        RECT 74.140 174.770 74.395 175.675 ;
        RECT 72.190 174.535 72.360 174.745 ;
        RECT 72.105 174.205 72.360 174.535 ;
        RECT 71.765 173.465 72.020 174.040 ;
        RECT 72.190 174.015 72.360 174.205 ;
        RECT 72.640 174.195 72.995 174.565 ;
        RECT 73.165 174.195 73.520 174.565 ;
        RECT 73.800 174.535 73.970 174.745 ;
        RECT 73.800 174.205 74.055 174.535 ;
        RECT 73.800 174.015 73.970 174.205 ;
        RECT 74.225 174.040 74.395 174.770 ;
        RECT 77.510 174.875 77.840 175.675 ;
        RECT 78.640 174.875 78.970 175.675 ;
        RECT 77.510 174.705 79.945 174.875 ;
        RECT 80.475 174.705 80.815 175.675 ;
        RECT 77.305 174.285 77.655 174.535 ;
        RECT 77.840 174.075 78.010 174.705 ;
        RECT 78.180 174.285 78.510 174.485 ;
        RECT 78.680 174.285 79.010 174.485 ;
        RECT 79.180 174.285 79.600 174.485 ;
        RECT 79.775 174.455 79.945 174.705 ;
        RECT 79.775 174.285 80.470 174.455 ;
        RECT 80.640 174.145 80.815 174.705 ;
        RECT 72.190 173.845 72.905 174.015 ;
        RECT 72.735 173.465 72.905 173.845 ;
        RECT 73.255 173.845 73.970 174.015 ;
        RECT 73.255 173.465 73.425 173.845 ;
        RECT 74.140 173.465 74.395 174.040 ;
        RECT 77.510 173.465 78.010 174.075 ;
        RECT 78.640 173.945 79.865 174.115 ;
        RECT 80.585 174.095 80.815 174.145 ;
        RECT 78.640 173.465 78.970 173.945 ;
        RECT 79.535 173.465 79.865 173.945 ;
        RECT 80.475 173.465 80.815 174.095 ;
        RECT 80.985 174.705 81.325 175.675 ;
        RECT 82.830 174.875 83.160 175.675 ;
        RECT 83.960 174.875 84.290 175.675 ;
        RECT 81.855 174.705 84.290 174.875 ;
        RECT 84.665 174.705 85.050 175.675 ;
        RECT 86.065 175.215 86.345 175.675 ;
        RECT 85.220 174.995 86.345 175.215 ;
        RECT 80.985 174.145 81.160 174.705 ;
        RECT 81.855 174.455 82.025 174.705 ;
        RECT 81.330 174.285 82.025 174.455 ;
        RECT 82.200 174.285 82.620 174.485 ;
        RECT 82.790 174.285 83.120 174.485 ;
        RECT 83.290 174.285 83.620 174.485 ;
        RECT 80.985 174.095 81.215 174.145 ;
        RECT 80.985 173.465 81.325 174.095 ;
        RECT 81.935 173.945 83.160 174.115 ;
        RECT 81.935 173.465 82.265 173.945 ;
        RECT 82.830 173.465 83.160 173.945 ;
        RECT 83.790 174.075 83.960 174.705 ;
        RECT 84.145 174.285 84.495 174.535 ;
        RECT 83.790 173.465 84.290 174.075 ;
        RECT 84.665 174.035 84.945 174.705 ;
        RECT 85.220 174.535 85.670 174.995 ;
        RECT 86.535 174.825 86.935 175.675 ;
        RECT 87.775 175.215 88.060 175.675 ;
        RECT 85.115 174.205 85.670 174.535 ;
        RECT 85.840 174.265 86.935 174.825 ;
        RECT 85.220 174.095 85.670 174.205 ;
        RECT 84.665 173.465 85.050 174.035 ;
        RECT 85.220 173.925 86.345 174.095 ;
        RECT 86.065 173.465 86.345 173.925 ;
        RECT 86.535 173.465 86.935 174.265 ;
        RECT 87.105 174.995 88.060 175.215 ;
        RECT 87.105 174.095 87.315 174.995 ;
        RECT 88.345 174.875 88.655 175.675 ;
        RECT 89.305 175.215 89.565 175.675 ;
        RECT 90.165 175.215 90.425 175.675 ;
        RECT 89.305 175.045 90.425 175.215 ;
        RECT 87.485 174.265 88.175 174.825 ;
        RECT 88.345 174.705 89.375 174.875 ;
        RECT 87.105 173.925 88.060 174.095 ;
        RECT 87.775 173.465 88.060 173.925 ;
        RECT 88.345 173.795 88.515 174.705 ;
        RECT 88.685 173.965 89.035 174.535 ;
        RECT 89.205 174.455 89.375 174.705 ;
        RECT 90.165 174.795 90.425 175.045 ;
        RECT 90.165 174.625 90.920 174.795 ;
        RECT 89.205 174.285 90.345 174.455 ;
        RECT 90.515 174.115 90.920 174.625 ;
        RECT 102.630 174.535 102.875 175.675 ;
        RECT 103.490 174.535 103.740 175.670 ;
        RECT 104.340 174.945 104.600 175.670 ;
        RECT 105.200 174.945 105.460 175.670 ;
        RECT 106.060 174.945 106.320 175.670 ;
        RECT 106.920 174.945 107.180 175.670 ;
        RECT 107.765 174.945 108.025 175.670 ;
        RECT 108.625 174.945 108.885 175.670 ;
        RECT 109.485 174.945 109.745 175.670 ;
        RECT 104.340 174.930 109.745 174.945 ;
        RECT 110.355 174.930 110.645 175.670 ;
        RECT 104.340 174.705 111.085 174.930 ;
        RECT 89.270 173.945 90.920 174.115 ;
        RECT 102.145 173.975 102.460 174.535 ;
        RECT 102.630 174.285 109.750 174.535 ;
        RECT 88.345 173.465 88.645 173.795 ;
        RECT 89.270 173.555 89.565 173.945 ;
        RECT 90.165 173.555 90.425 173.945 ;
        RECT 102.630 173.475 102.880 174.285 ;
        RECT 103.490 173.475 103.740 174.285 ;
        RECT 109.920 174.145 111.085 174.705 ;
        RECT 111.345 174.705 111.685 175.675 ;
        RECT 113.190 174.875 113.520 175.675 ;
        RECT 114.320 174.875 114.650 175.675 ;
        RECT 112.215 174.705 114.650 174.875 ;
        RECT 115.230 174.875 115.560 175.675 ;
        RECT 116.360 174.875 116.690 175.675 ;
        RECT 115.230 174.705 117.665 174.875 ;
        RECT 118.195 174.705 118.535 175.675 ;
        RECT 111.345 174.655 111.575 174.705 ;
        RECT 109.920 174.115 111.115 174.145 ;
        RECT 104.340 173.975 111.115 174.115 ;
        RECT 111.345 174.095 111.520 174.655 ;
        RECT 112.215 174.455 112.385 174.705 ;
        RECT 111.690 174.285 112.385 174.455 ;
        RECT 112.555 174.315 112.980 174.485 ;
        RECT 112.560 174.285 112.980 174.315 ;
        RECT 113.150 174.285 113.480 174.485 ;
        RECT 113.650 174.285 113.980 174.485 ;
        RECT 104.340 173.945 111.085 173.975 ;
        RECT 104.340 173.490 104.600 173.945 ;
        RECT 105.200 173.490 105.460 173.945 ;
        RECT 106.060 173.490 106.320 173.945 ;
        RECT 106.905 173.490 107.180 173.945 ;
        RECT 107.765 173.490 108.025 173.945 ;
        RECT 108.625 173.490 108.885 173.945 ;
        RECT 109.485 173.490 109.745 173.945 ;
        RECT 110.355 173.490 110.615 173.945 ;
        RECT 111.345 173.465 111.685 174.095 ;
        RECT 112.295 173.945 113.520 174.115 ;
        RECT 112.295 173.465 112.625 173.945 ;
        RECT 113.190 173.465 113.520 173.945 ;
        RECT 114.150 174.075 114.320 174.705 ;
        RECT 114.505 174.285 114.855 174.535 ;
        RECT 115.025 174.285 115.375 174.535 ;
        RECT 115.560 174.075 115.730 174.705 ;
        RECT 115.900 174.285 116.230 174.485 ;
        RECT 116.400 174.285 116.730 174.485 ;
        RECT 116.900 174.285 117.320 174.485 ;
        RECT 117.495 174.455 117.665 174.705 ;
        RECT 117.495 174.285 118.190 174.455 ;
        RECT 114.150 173.465 114.650 174.075 ;
        RECT 115.230 173.465 115.730 174.075 ;
        RECT 116.360 173.945 117.585 174.115 ;
        RECT 118.360 174.095 118.535 174.705 ;
        RECT 116.360 173.465 116.690 173.945 ;
        RECT 117.255 173.465 117.585 173.945 ;
        RECT 118.195 173.465 118.535 174.095 ;
        RECT 119.145 174.695 119.475 175.675 ;
        RECT 119.145 174.095 119.395 174.695 ;
        RECT 119.565 174.285 119.895 174.535 ;
        RECT 119.145 173.465 119.475 174.095 ;
        RECT 33.810 172.345 34.310 172.955 ;
        RECT 33.605 171.885 33.955 172.135 ;
        RECT 34.140 171.715 34.310 172.345 ;
        RECT 34.940 172.475 35.270 172.955 ;
        RECT 35.835 172.475 36.165 172.955 ;
        RECT 34.940 172.305 36.165 172.475 ;
        RECT 36.775 172.325 37.115 172.955 ;
        RECT 34.480 171.935 34.810 172.135 ;
        RECT 34.980 171.935 35.310 172.135 ;
        RECT 35.480 171.935 35.900 172.135 ;
        RECT 36.075 171.965 36.770 172.135 ;
        RECT 36.075 171.715 36.245 171.965 ;
        RECT 36.940 171.715 37.115 172.325 ;
        RECT 33.810 171.545 36.245 171.715 ;
        RECT 33.810 170.745 34.140 171.545 ;
        RECT 34.940 170.745 35.270 171.545 ;
        RECT 36.775 170.745 37.115 171.715 ;
        RECT 38.205 172.325 38.545 172.955 ;
        RECT 39.155 172.475 39.485 172.955 ;
        RECT 40.050 172.475 40.380 172.955 ;
        RECT 38.205 171.715 38.380 172.325 ;
        RECT 39.155 172.305 40.380 172.475 ;
        RECT 41.010 172.345 41.510 172.955 ;
        RECT 45.205 172.475 45.465 172.930 ;
        RECT 46.075 172.475 46.335 172.930 ;
        RECT 46.935 172.475 47.195 172.930 ;
        RECT 47.795 172.475 48.055 172.930 ;
        RECT 48.640 172.475 48.915 172.930 ;
        RECT 49.500 172.475 49.760 172.930 ;
        RECT 50.360 172.475 50.620 172.930 ;
        RECT 51.220 172.475 51.480 172.930 ;
        RECT 38.550 171.965 39.245 172.135 ;
        RECT 39.075 171.715 39.245 171.965 ;
        RECT 39.420 171.935 39.840 172.135 ;
        RECT 40.010 171.935 40.340 172.135 ;
        RECT 40.510 171.935 40.840 172.135 ;
        RECT 41.010 171.715 41.180 172.345 ;
        RECT 44.735 172.305 51.480 172.475 ;
        RECT 41.365 171.885 41.715 172.135 ;
        RECT 44.735 171.715 45.900 172.305 ;
        RECT 52.080 172.135 52.330 172.945 ;
        RECT 52.940 172.135 53.190 172.945 ;
        RECT 46.070 171.885 53.190 172.135 ;
        RECT 53.360 171.885 53.675 172.445 ;
        RECT 53.850 172.415 54.105 172.945 ;
        RECT 54.825 172.745 55.895 172.915 ;
        RECT 38.205 170.745 38.545 171.715 ;
        RECT 39.075 171.545 41.510 171.715 ;
        RECT 40.050 170.745 40.380 171.545 ;
        RECT 41.180 170.745 41.510 171.545 ;
        RECT 44.735 171.490 51.480 171.715 ;
        RECT 45.175 170.750 45.465 171.490 ;
        RECT 46.075 171.475 51.480 171.490 ;
        RECT 46.075 170.750 46.335 171.475 ;
        RECT 46.935 170.750 47.195 171.475 ;
        RECT 47.795 170.750 48.055 171.475 ;
        RECT 48.640 170.750 48.900 171.475 ;
        RECT 49.500 170.750 49.760 171.475 ;
        RECT 50.360 170.750 50.620 171.475 ;
        RECT 51.220 170.750 51.480 171.475 ;
        RECT 52.080 170.750 52.330 171.885 ;
        RECT 52.945 170.745 53.190 171.885 ;
        RECT 53.850 171.765 54.060 172.415 ;
        RECT 54.825 172.390 55.145 172.745 ;
        RECT 54.820 172.215 55.145 172.390 ;
        RECT 54.230 171.915 55.145 172.215 ;
        RECT 55.315 172.175 55.555 172.575 ;
        RECT 55.725 172.515 55.895 172.745 ;
        RECT 56.425 172.675 57.375 172.955 ;
        RECT 57.595 172.765 57.945 172.935 ;
        RECT 55.725 172.345 56.255 172.515 ;
        RECT 54.230 171.885 54.970 171.915 ;
        RECT 53.850 170.885 54.105 171.765 ;
        RECT 54.800 171.295 54.970 171.885 ;
        RECT 55.315 171.805 55.855 172.175 ;
        RECT 56.035 172.065 56.255 172.345 ;
        RECT 56.425 171.895 56.595 172.675 ;
        RECT 56.190 171.725 56.595 171.895 ;
        RECT 56.765 171.885 57.115 172.505 ;
        RECT 56.190 171.635 56.360 171.725 ;
        RECT 57.285 171.715 57.495 172.505 ;
        RECT 55.140 171.465 56.360 171.635 ;
        RECT 56.820 171.555 57.495 171.715 ;
        RECT 54.800 171.125 55.600 171.295 ;
        RECT 55.430 170.835 55.600 171.125 ;
        RECT 56.190 171.085 56.360 171.465 ;
        RECT 56.530 171.545 57.495 171.555 ;
        RECT 57.685 172.375 57.945 172.765 ;
        RECT 59.360 172.735 60.215 172.905 ;
        RECT 60.420 172.735 60.915 172.905 ;
        RECT 57.685 171.685 57.855 172.375 ;
        RECT 58.025 172.025 58.195 172.205 ;
        RECT 58.365 172.195 59.155 172.445 ;
        RECT 59.360 172.025 59.530 172.735 ;
        RECT 59.700 172.225 60.055 172.445 ;
        RECT 58.025 171.855 59.715 172.025 ;
        RECT 56.530 171.255 56.990 171.545 ;
        RECT 57.685 171.515 59.185 171.685 ;
        RECT 57.685 171.375 57.855 171.515 ;
        RECT 57.295 171.205 57.855 171.375 ;
        RECT 56.190 170.745 57.060 171.085 ;
        RECT 57.295 170.745 57.465 171.205 ;
        RECT 58.300 171.175 59.375 171.345 ;
        RECT 58.300 170.835 58.470 171.175 ;
        RECT 59.205 170.835 59.375 171.175 ;
        RECT 59.545 171.075 59.715 171.855 ;
        RECT 59.885 171.635 60.055 172.225 ;
        RECT 60.225 171.825 60.575 172.445 ;
        RECT 59.885 171.245 60.350 171.635 ;
        RECT 60.745 171.375 60.915 172.735 ;
        RECT 61.085 171.545 61.545 172.595 ;
        RECT 60.520 171.205 60.915 171.375 ;
        RECT 60.520 171.075 60.690 171.205 ;
        RECT 59.545 170.745 60.225 171.075 ;
        RECT 60.440 170.745 60.690 171.075 ;
        RECT 61.280 170.760 61.605 171.545 ;
        RECT 61.775 170.745 61.945 172.865 ;
        RECT 62.615 172.575 62.870 172.865 ;
        RECT 62.120 172.405 62.870 172.575 ;
        RECT 62.120 171.415 62.350 172.405 ;
        RECT 63.945 172.325 64.275 172.955 ;
        RECT 82.455 172.475 82.625 172.955 ;
        RECT 83.295 172.475 83.465 172.955 ;
        RECT 84.135 172.475 84.305 172.955 ;
        RECT 62.520 171.585 62.870 172.235 ;
        RECT 63.945 171.725 64.195 172.325 ;
        RECT 82.455 172.305 83.090 172.475 ;
        RECT 83.295 172.305 84.305 172.475 ;
        RECT 85.240 172.495 85.525 172.955 ;
        RECT 85.240 172.325 86.195 172.495 ;
        RECT 82.920 172.135 83.090 172.305 ;
        RECT 83.805 172.275 84.305 172.305 ;
        RECT 64.365 171.885 64.695 172.135 ;
        RECT 82.370 171.895 82.750 172.135 ;
        RECT 82.920 171.965 83.420 172.135 ;
        RECT 82.920 171.725 83.090 171.965 ;
        RECT 83.810 171.765 84.305 172.275 ;
        RECT 62.120 171.245 62.870 171.415 ;
        RECT 62.615 170.745 62.870 171.245 ;
        RECT 63.945 170.745 64.275 171.725 ;
        RECT 82.375 171.555 83.090 171.725 ;
        RECT 83.295 171.595 84.305 171.765 ;
        RECT 85.125 171.595 85.815 172.155 ;
        RECT 82.375 170.745 82.705 171.555 ;
        RECT 83.295 170.745 83.465 171.595 ;
        RECT 84.135 170.745 84.305 171.595 ;
        RECT 85.985 171.425 86.195 172.325 ;
        RECT 85.240 171.205 86.195 171.425 ;
        RECT 86.365 172.155 86.765 172.955 ;
        RECT 86.955 172.495 87.235 172.955 ;
        RECT 86.955 172.325 88.080 172.495 ;
        RECT 88.250 172.385 88.635 172.955 ;
        RECT 87.630 172.215 88.080 172.325 ;
        RECT 86.365 171.595 87.460 172.155 ;
        RECT 87.630 171.885 88.185 172.215 ;
        RECT 85.240 170.745 85.525 171.205 ;
        RECT 86.365 170.745 86.765 171.595 ;
        RECT 87.630 171.425 88.080 171.885 ;
        RECT 88.355 171.715 88.635 172.385 ;
        RECT 90.165 172.325 90.495 172.955 ;
        RECT 89.745 171.885 90.075 172.135 ;
        RECT 90.245 171.725 90.495 172.325 ;
        RECT 86.955 171.205 88.080 171.425 ;
        RECT 86.955 170.745 87.235 171.205 ;
        RECT 88.250 170.745 88.635 171.715 ;
        RECT 90.165 170.745 90.495 171.725 ;
        RECT 91.110 172.415 91.365 172.945 ;
        RECT 92.085 172.745 93.155 172.915 ;
        RECT 91.110 171.765 91.320 172.415 ;
        RECT 92.085 172.390 92.405 172.745 ;
        RECT 92.080 172.215 92.405 172.390 ;
        RECT 91.490 171.915 92.405 172.215 ;
        RECT 92.575 172.175 92.815 172.575 ;
        RECT 92.985 172.515 93.155 172.745 ;
        RECT 93.685 172.675 94.635 172.955 ;
        RECT 94.855 172.765 95.205 172.935 ;
        RECT 92.985 172.345 93.515 172.515 ;
        RECT 91.490 171.885 92.230 171.915 ;
        RECT 91.110 170.885 91.365 171.765 ;
        RECT 92.060 171.295 92.230 171.885 ;
        RECT 92.575 171.805 93.115 172.175 ;
        RECT 93.295 172.065 93.515 172.345 ;
        RECT 93.685 171.895 93.855 172.675 ;
        RECT 93.450 171.725 93.855 171.895 ;
        RECT 94.025 171.885 94.375 172.505 ;
        RECT 93.450 171.635 93.620 171.725 ;
        RECT 94.545 171.715 94.755 172.505 ;
        RECT 92.400 171.465 93.620 171.635 ;
        RECT 94.080 171.555 94.755 171.715 ;
        RECT 92.060 171.125 92.860 171.295 ;
        RECT 92.690 170.835 92.860 171.125 ;
        RECT 93.450 171.085 93.620 171.465 ;
        RECT 93.790 171.545 94.755 171.555 ;
        RECT 94.945 172.375 95.205 172.765 ;
        RECT 96.620 172.735 97.475 172.905 ;
        RECT 97.680 172.735 98.175 172.905 ;
        RECT 94.945 171.685 95.115 172.375 ;
        RECT 95.285 172.025 95.455 172.205 ;
        RECT 95.625 172.195 96.415 172.445 ;
        RECT 96.620 172.025 96.790 172.735 ;
        RECT 96.960 172.225 97.315 172.445 ;
        RECT 95.285 171.855 96.975 172.025 ;
        RECT 93.790 171.255 94.250 171.545 ;
        RECT 94.945 171.515 96.445 171.685 ;
        RECT 94.945 171.375 95.115 171.515 ;
        RECT 94.555 171.205 95.115 171.375 ;
        RECT 93.450 170.745 94.320 171.085 ;
        RECT 94.555 170.745 94.725 171.205 ;
        RECT 95.560 171.175 96.635 171.345 ;
        RECT 95.560 170.835 95.730 171.175 ;
        RECT 96.465 170.835 96.635 171.175 ;
        RECT 96.805 171.075 96.975 171.855 ;
        RECT 97.145 171.635 97.315 172.225 ;
        RECT 97.485 171.825 97.835 172.445 ;
        RECT 97.145 171.245 97.610 171.635 ;
        RECT 98.005 171.375 98.175 172.735 ;
        RECT 98.345 171.545 98.805 172.595 ;
        RECT 97.780 171.205 98.175 171.375 ;
        RECT 97.780 171.075 97.950 171.205 ;
        RECT 96.805 170.745 97.485 171.075 ;
        RECT 97.700 170.745 97.950 171.075 ;
        RECT 98.540 170.760 98.865 171.545 ;
        RECT 99.035 170.745 99.205 172.865 ;
        RECT 99.875 172.575 100.130 172.865 ;
        RECT 99.380 172.405 100.130 172.575 ;
        RECT 105.895 172.485 106.150 172.930 ;
        RECT 106.750 172.485 107.010 172.930 ;
        RECT 99.380 171.415 99.610 172.405 ;
        RECT 104.905 172.315 107.935 172.485 ;
        RECT 99.780 171.585 100.130 172.235 ;
        RECT 104.905 171.750 105.205 172.315 ;
        RECT 105.380 171.920 107.595 172.145 ;
        RECT 107.765 171.750 107.935 172.315 ;
        RECT 104.905 171.580 107.935 171.750 ;
        RECT 108.125 172.325 108.465 172.955 ;
        RECT 109.075 172.475 109.405 172.955 ;
        RECT 109.970 172.475 110.300 172.955 ;
        RECT 108.125 171.715 108.300 172.325 ;
        RECT 109.075 172.305 110.300 172.475 ;
        RECT 110.930 172.345 111.430 172.955 ;
        RECT 108.470 171.965 109.165 172.135 ;
        RECT 108.995 171.715 109.165 171.965 ;
        RECT 109.340 171.935 109.760 172.135 ;
        RECT 109.930 171.935 110.260 172.135 ;
        RECT 110.430 171.935 110.760 172.135 ;
        RECT 110.930 171.715 111.100 172.345 ;
        RECT 113.625 172.325 113.955 172.955 ;
        RECT 111.285 171.885 111.635 172.135 ;
        RECT 113.205 171.885 113.535 172.135 ;
        RECT 113.705 171.725 113.955 172.325 ;
        RECT 99.380 171.245 100.130 171.415 ;
        RECT 99.875 170.745 100.130 171.245 ;
        RECT 105.460 170.775 105.720 171.580 ;
        RECT 106.320 170.775 106.575 171.580 ;
        RECT 107.180 170.775 107.435 171.580 ;
        RECT 108.125 170.745 108.465 171.715 ;
        RECT 108.995 171.545 111.430 171.715 ;
        RECT 109.970 170.745 110.300 171.545 ;
        RECT 111.100 170.745 111.430 171.545 ;
        RECT 113.625 170.745 113.955 171.725 ;
        RECT 115.950 172.415 116.205 172.945 ;
        RECT 116.925 172.745 117.995 172.915 ;
        RECT 115.950 171.765 116.160 172.415 ;
        RECT 116.925 172.390 117.245 172.745 ;
        RECT 116.920 172.215 117.245 172.390 ;
        RECT 116.330 171.915 117.245 172.215 ;
        RECT 117.415 172.175 117.655 172.575 ;
        RECT 117.825 172.515 117.995 172.745 ;
        RECT 118.525 172.675 119.475 172.955 ;
        RECT 119.695 172.765 120.045 172.935 ;
        RECT 117.825 172.345 118.355 172.515 ;
        RECT 116.330 171.885 117.070 171.915 ;
        RECT 115.950 170.885 116.205 171.765 ;
        RECT 116.900 171.295 117.070 171.885 ;
        RECT 117.415 171.805 117.955 172.175 ;
        RECT 118.135 172.065 118.355 172.345 ;
        RECT 118.525 171.895 118.695 172.675 ;
        RECT 118.290 171.725 118.695 171.895 ;
        RECT 118.865 171.885 119.215 172.505 ;
        RECT 118.290 171.635 118.460 171.725 ;
        RECT 119.385 171.715 119.595 172.505 ;
        RECT 117.240 171.465 118.460 171.635 ;
        RECT 118.920 171.555 119.595 171.715 ;
        RECT 116.900 171.125 117.700 171.295 ;
        RECT 117.530 170.835 117.700 171.125 ;
        RECT 118.290 171.085 118.460 171.465 ;
        RECT 118.630 171.545 119.595 171.555 ;
        RECT 119.785 172.375 120.045 172.765 ;
        RECT 121.460 172.735 122.315 172.905 ;
        RECT 122.520 172.735 123.015 172.905 ;
        RECT 119.785 171.685 119.955 172.375 ;
        RECT 120.125 172.025 120.295 172.205 ;
        RECT 120.465 172.195 121.255 172.445 ;
        RECT 121.460 172.025 121.630 172.735 ;
        RECT 121.800 172.225 122.155 172.445 ;
        RECT 120.125 171.855 121.815 172.025 ;
        RECT 118.630 171.255 119.090 171.545 ;
        RECT 119.785 171.515 121.285 171.685 ;
        RECT 119.785 171.375 119.955 171.515 ;
        RECT 119.395 171.205 119.955 171.375 ;
        RECT 118.290 170.745 119.160 171.085 ;
        RECT 119.395 170.745 119.565 171.205 ;
        RECT 120.400 171.175 121.475 171.345 ;
        RECT 120.400 170.835 120.570 171.175 ;
        RECT 121.305 170.835 121.475 171.175 ;
        RECT 121.645 171.075 121.815 171.855 ;
        RECT 121.985 171.635 122.155 172.225 ;
        RECT 122.325 171.825 122.675 172.445 ;
        RECT 121.985 171.245 122.450 171.635 ;
        RECT 122.845 171.375 123.015 172.735 ;
        RECT 123.185 171.545 123.645 172.595 ;
        RECT 122.620 171.205 123.015 171.375 ;
        RECT 122.620 171.075 122.790 171.205 ;
        RECT 121.645 170.745 122.325 171.075 ;
        RECT 122.540 170.745 122.790 171.075 ;
        RECT 123.380 170.760 123.705 171.545 ;
        RECT 123.875 170.745 124.045 172.865 ;
        RECT 124.715 172.575 124.970 172.865 ;
        RECT 124.220 172.405 124.970 172.575 ;
        RECT 124.220 171.415 124.450 172.405 ;
        RECT 124.620 171.585 124.970 172.235 ;
        RECT 124.220 171.245 124.970 171.415 ;
        RECT 124.715 170.745 124.970 171.245 ;
        RECT 27.605 169.255 27.935 170.235 ;
        RECT 30.825 169.255 31.155 170.235 ;
        RECT 31.880 169.775 32.165 170.235 ;
        RECT 31.880 169.555 32.835 169.775 ;
        RECT 27.605 168.655 27.855 169.255 ;
        RECT 28.025 168.845 28.355 169.095 ;
        RECT 30.825 168.655 31.075 169.255 ;
        RECT 31.245 168.845 31.575 169.095 ;
        RECT 31.765 168.825 32.455 169.385 ;
        RECT 32.625 168.655 32.835 169.555 ;
        RECT 27.605 168.025 27.935 168.655 ;
        RECT 30.825 168.025 31.155 168.655 ;
        RECT 31.880 168.485 32.835 168.655 ;
        RECT 33.005 169.385 33.405 170.235 ;
        RECT 33.595 169.775 33.875 170.235 ;
        RECT 33.595 169.555 34.720 169.775 ;
        RECT 33.005 168.825 34.100 169.385 ;
        RECT 34.270 169.095 34.720 169.555 ;
        RECT 34.890 169.265 35.275 170.235 ;
        RECT 31.880 168.025 32.165 168.485 ;
        RECT 33.005 168.025 33.405 168.825 ;
        RECT 34.270 168.765 34.825 169.095 ;
        RECT 34.270 168.655 34.720 168.765 ;
        RECT 33.595 168.485 34.720 168.655 ;
        RECT 34.995 168.595 35.275 169.265 ;
        RECT 36.105 169.065 36.435 170.235 ;
        RECT 37.165 169.065 37.525 170.235 ;
        RECT 45.565 169.265 45.905 170.235 ;
        RECT 47.410 169.435 47.740 170.235 ;
        RECT 48.540 169.435 48.870 170.235 ;
        RECT 46.435 169.265 48.870 169.435 ;
        RECT 53.020 169.400 53.280 170.205 ;
        RECT 53.880 169.400 54.135 170.205 ;
        RECT 54.740 169.400 54.995 170.205 ;
        RECT 68.655 169.475 68.825 170.235 ;
        RECT 36.105 168.785 37.525 169.065 ;
        RECT 33.595 168.025 33.875 168.485 ;
        RECT 34.890 168.025 35.275 168.595 ;
        RECT 37.165 168.450 37.525 168.785 ;
        RECT 37.695 168.515 38.035 169.095 ;
        RECT 45.565 168.655 45.740 169.265 ;
        RECT 46.435 169.015 46.605 169.265 ;
        RECT 45.910 168.845 46.605 169.015 ;
        RECT 46.780 168.845 47.200 169.045 ;
        RECT 47.370 168.845 47.700 169.045 ;
        RECT 47.870 168.845 48.200 169.045 ;
        RECT 36.905 168.025 37.525 168.450 ;
        RECT 45.565 168.025 45.905 168.655 ;
        RECT 46.515 168.505 47.740 168.675 ;
        RECT 46.515 168.025 46.845 168.505 ;
        RECT 47.410 168.025 47.740 168.505 ;
        RECT 48.370 168.635 48.540 169.265 ;
        RECT 52.465 169.230 55.495 169.400 ;
        RECT 68.655 169.305 69.370 169.475 ;
        RECT 69.540 169.330 69.795 170.235 ;
        RECT 48.725 168.845 49.075 169.095 ;
        RECT 52.465 168.665 52.765 169.230 ;
        RECT 52.940 168.835 55.155 169.060 ;
        RECT 55.325 168.665 55.495 169.230 ;
        RECT 68.565 168.755 68.920 169.125 ;
        RECT 69.200 169.095 69.370 169.305 ;
        RECT 69.200 168.765 69.455 169.095 ;
        RECT 48.370 168.025 48.870 168.635 ;
        RECT 52.465 168.495 55.495 168.665 ;
        RECT 69.200 168.575 69.370 168.765 ;
        RECT 69.625 168.600 69.795 169.330 ;
        RECT 53.455 168.050 53.710 168.495 ;
        RECT 54.310 168.050 54.570 168.495 ;
        RECT 68.655 168.405 69.370 168.575 ;
        RECT 68.655 168.025 68.825 168.405 ;
        RECT 69.540 168.025 69.795 168.600 ;
        RECT 70.845 169.330 71.100 170.235 ;
        RECT 71.815 169.475 71.985 170.235 ;
        RECT 70.845 168.600 71.015 169.330 ;
        RECT 71.270 169.305 71.985 169.475 ;
        RECT 72.705 169.435 73.015 170.235 ;
        RECT 73.665 169.775 73.925 170.235 ;
        RECT 74.525 169.775 74.785 170.235 ;
        RECT 77.475 170.065 79.505 170.235 ;
        RECT 73.665 169.605 74.785 169.775 ;
        RECT 71.270 169.095 71.440 169.305 ;
        RECT 72.705 169.265 73.735 169.435 ;
        RECT 71.185 168.765 71.440 169.095 ;
        RECT 70.845 168.025 71.100 168.600 ;
        RECT 71.270 168.575 71.440 168.765 ;
        RECT 71.720 168.755 72.075 169.125 ;
        RECT 71.270 168.405 71.985 168.575 ;
        RECT 71.815 168.025 71.985 168.405 ;
        RECT 72.705 168.355 72.875 169.265 ;
        RECT 73.045 168.525 73.395 169.095 ;
        RECT 73.565 169.015 73.735 169.265 ;
        RECT 74.525 169.355 74.785 169.605 ;
        RECT 76.385 169.645 76.900 170.055 ;
        RECT 74.525 169.185 75.280 169.355 ;
        RECT 73.565 168.845 74.705 169.015 ;
        RECT 74.875 168.675 75.280 169.185 ;
        RECT 73.630 168.505 75.280 168.675 ;
        RECT 76.385 168.835 76.725 169.645 ;
        RECT 77.475 169.400 77.645 170.065 ;
        RECT 78.040 169.725 79.165 169.895 ;
        RECT 76.895 169.210 77.645 169.400 ;
        RECT 77.815 169.385 78.825 169.555 ;
        RECT 76.385 168.665 77.615 168.835 ;
        RECT 72.705 168.025 73.005 168.355 ;
        RECT 73.630 168.115 73.925 168.505 ;
        RECT 74.525 168.115 74.785 168.505 ;
        RECT 76.660 168.060 76.905 168.665 ;
        RECT 77.815 168.025 78.005 169.385 ;
        RECT 78.175 168.365 78.450 169.185 ;
        RECT 78.655 168.585 78.825 169.385 ;
        RECT 78.995 168.595 79.165 169.725 ;
        RECT 79.335 169.095 79.505 170.065 ;
        RECT 80.015 169.265 80.350 170.235 ;
        RECT 79.335 168.765 79.530 169.095 ;
        RECT 79.755 168.765 80.010 169.095 ;
        RECT 79.755 168.595 79.925 168.765 ;
        RECT 80.180 168.595 80.350 169.265 ;
        RECT 80.900 169.425 81.155 170.095 ;
        RECT 81.800 169.685 82.130 170.195 ;
        RECT 80.900 168.705 81.080 169.425 ;
        RECT 81.800 169.095 82.050 169.685 ;
        RECT 82.400 169.535 82.570 170.145 ;
        RECT 83.300 169.855 83.540 170.145 ;
        RECT 84.340 169.935 84.970 170.185 ;
        RECT 84.340 169.855 84.510 169.935 ;
        RECT 85.940 169.855 86.110 170.145 ;
        RECT 86.910 170.020 87.740 170.190 ;
        RECT 83.300 169.685 84.510 169.855 ;
        RECT 81.250 168.765 82.050 169.095 ;
        RECT 78.995 168.425 79.925 168.595 ;
        RECT 78.995 168.390 79.170 168.425 ;
        RECT 78.175 168.195 78.455 168.365 ;
        RECT 78.175 168.025 78.450 168.195 ;
        RECT 78.640 168.025 79.170 168.390 ;
        RECT 80.095 168.025 80.350 168.595 ;
        RECT 80.815 168.565 81.080 168.705 ;
        RECT 80.815 168.535 81.155 168.565 ;
        RECT 80.900 168.035 81.155 168.535 ;
        RECT 81.800 168.115 82.050 168.765 ;
        RECT 82.250 169.515 82.570 169.535 ;
        RECT 82.250 169.345 84.170 169.515 ;
        RECT 82.250 168.450 82.440 169.345 ;
        RECT 84.340 169.175 84.510 169.685 ;
        RECT 84.680 169.425 85.200 169.735 ;
        RECT 82.610 169.005 84.510 169.175 ;
        RECT 82.610 168.945 82.940 169.005 ;
        RECT 83.090 168.775 83.420 168.835 ;
        RECT 82.760 168.505 83.420 168.775 ;
        RECT 82.250 168.120 82.570 168.450 ;
        RECT 83.610 168.245 83.780 169.005 ;
        RECT 84.680 168.835 84.860 169.245 ;
        RECT 83.950 168.665 84.280 168.785 ;
        RECT 85.030 168.665 85.200 169.425 ;
        RECT 83.950 168.495 85.200 168.665 ;
        RECT 85.370 169.605 86.740 169.855 ;
        RECT 85.370 168.835 85.560 169.605 ;
        RECT 86.490 169.345 86.740 169.605 ;
        RECT 85.730 169.175 85.980 169.335 ;
        RECT 86.910 169.175 87.080 170.020 ;
        RECT 87.975 169.735 88.145 170.235 ;
        RECT 87.250 169.345 87.750 169.725 ;
        RECT 87.975 169.565 88.670 169.735 ;
        RECT 85.730 169.005 87.080 169.175 ;
        RECT 86.660 168.965 87.080 169.005 ;
        RECT 85.370 168.495 85.790 168.835 ;
        RECT 86.080 168.505 86.490 168.835 ;
        RECT 83.610 168.075 84.460 168.245 ;
        RECT 85.540 168.065 85.790 168.495 ;
        RECT 86.660 168.235 86.830 168.965 ;
        RECT 87.000 168.415 87.350 168.785 ;
        RECT 87.530 168.475 87.750 169.345 ;
        RECT 87.920 168.775 88.330 169.395 ;
        RECT 88.500 168.595 88.670 169.565 ;
        RECT 87.975 168.405 88.670 168.595 ;
        RECT 86.660 168.035 87.675 168.235 ;
        RECT 87.975 168.075 88.145 168.405 ;
        RECT 88.860 168.115 89.085 170.235 ;
        RECT 89.755 169.735 89.925 170.235 ;
        RECT 92.195 170.065 94.225 170.235 ;
        RECT 89.260 169.565 89.925 169.735 ;
        RECT 91.105 169.645 91.620 170.055 ;
        RECT 89.260 168.575 89.490 169.565 ;
        RECT 89.660 168.745 90.010 169.395 ;
        RECT 91.105 168.835 91.445 169.645 ;
        RECT 92.195 169.400 92.365 170.065 ;
        RECT 92.760 169.725 93.885 169.895 ;
        RECT 91.615 169.210 92.365 169.400 ;
        RECT 92.535 169.385 93.545 169.555 ;
        RECT 91.105 168.665 92.335 168.835 ;
        RECT 89.260 168.405 89.925 168.575 ;
        RECT 89.755 168.115 89.925 168.405 ;
        RECT 91.380 168.060 91.625 168.665 ;
        RECT 92.535 168.025 92.725 169.385 ;
        RECT 92.895 169.045 93.170 169.185 ;
        RECT 92.895 168.875 93.175 169.045 ;
        RECT 92.895 168.025 93.170 168.875 ;
        RECT 93.375 168.585 93.545 169.385 ;
        RECT 93.715 168.595 93.885 169.725 ;
        RECT 94.055 169.095 94.225 170.065 ;
        RECT 94.735 169.265 95.070 170.235 ;
        RECT 96.255 169.475 96.425 170.235 ;
        RECT 96.255 169.305 96.920 169.475 ;
        RECT 97.105 169.330 97.375 170.235 ;
        RECT 94.055 168.765 94.250 169.095 ;
        RECT 94.475 168.765 94.730 169.095 ;
        RECT 94.475 168.595 94.645 168.765 ;
        RECT 94.900 168.595 95.070 169.265 ;
        RECT 96.750 169.160 96.920 169.305 ;
        RECT 96.185 168.755 96.515 169.125 ;
        RECT 96.750 168.830 97.035 169.160 ;
        RECT 93.715 168.425 94.645 168.595 ;
        RECT 93.715 168.390 93.890 168.425 ;
        RECT 93.360 168.025 93.890 168.390 ;
        RECT 94.815 168.025 95.070 168.595 ;
        RECT 96.750 168.575 96.920 168.830 ;
        RECT 96.255 168.405 96.920 168.575 ;
        RECT 97.205 168.530 97.375 169.330 ;
        RECT 96.255 168.025 96.425 168.405 ;
        RECT 97.115 168.025 97.375 168.530 ;
        RECT 102.610 169.215 102.865 170.095 ;
        RECT 104.190 169.855 104.360 170.145 ;
        RECT 103.560 169.685 104.360 169.855 ;
        RECT 104.950 169.895 105.820 170.235 ;
        RECT 102.610 168.565 102.820 169.215 ;
        RECT 103.560 169.095 103.730 169.685 ;
        RECT 104.950 169.515 105.120 169.895 ;
        RECT 106.055 169.775 106.225 170.235 ;
        RECT 107.060 169.805 107.230 170.145 ;
        RECT 107.965 169.805 108.135 170.145 ;
        RECT 103.900 169.345 105.120 169.515 ;
        RECT 105.290 169.435 105.750 169.725 ;
        RECT 106.055 169.605 106.615 169.775 ;
        RECT 107.060 169.635 108.135 169.805 ;
        RECT 108.305 169.905 108.985 170.235 ;
        RECT 109.200 169.905 109.450 170.235 ;
        RECT 106.445 169.465 106.615 169.605 ;
        RECT 105.290 169.425 106.255 169.435 ;
        RECT 104.950 169.255 105.120 169.345 ;
        RECT 105.580 169.265 106.255 169.425 ;
        RECT 102.990 169.065 103.730 169.095 ;
        RECT 102.990 168.765 103.905 169.065 ;
        RECT 103.580 168.590 103.905 168.765 ;
        RECT 102.610 168.035 102.865 168.565 ;
        RECT 103.585 168.235 103.905 168.590 ;
        RECT 104.075 168.805 104.615 169.175 ;
        RECT 104.950 169.085 105.355 169.255 ;
        RECT 104.075 168.405 104.315 168.805 ;
        RECT 104.795 168.635 105.015 168.915 ;
        RECT 104.485 168.465 105.015 168.635 ;
        RECT 104.485 168.235 104.655 168.465 ;
        RECT 103.585 168.065 104.655 168.235 ;
        RECT 105.185 168.305 105.355 169.085 ;
        RECT 105.525 168.475 105.875 169.095 ;
        RECT 106.045 168.475 106.255 169.265 ;
        RECT 106.445 169.295 107.945 169.465 ;
        RECT 106.445 168.605 106.615 169.295 ;
        RECT 108.305 169.125 108.475 169.905 ;
        RECT 109.280 169.775 109.450 169.905 ;
        RECT 106.785 168.955 108.475 169.125 ;
        RECT 108.645 169.345 109.110 169.735 ;
        RECT 109.280 169.605 109.675 169.775 ;
        RECT 106.785 168.775 106.955 168.955 ;
        RECT 105.185 168.025 106.135 168.305 ;
        RECT 106.445 168.215 106.705 168.605 ;
        RECT 107.125 168.535 107.915 168.785 ;
        RECT 106.355 168.045 106.705 168.215 ;
        RECT 108.120 168.245 108.290 168.955 ;
        RECT 108.645 168.755 108.815 169.345 ;
        RECT 108.460 168.535 108.815 168.755 ;
        RECT 108.985 168.535 109.335 169.155 ;
        RECT 109.505 168.245 109.675 169.605 ;
        RECT 110.040 169.435 110.365 170.220 ;
        RECT 109.845 168.385 110.305 169.435 ;
        RECT 108.120 168.075 108.975 168.245 ;
        RECT 109.180 168.075 109.675 168.245 ;
        RECT 110.535 168.115 110.705 170.235 ;
        RECT 111.375 169.735 111.630 170.235 ;
        RECT 110.880 169.565 111.630 169.735 ;
        RECT 110.880 168.575 111.110 169.565 ;
        RECT 111.280 168.745 111.630 169.395 ;
        RECT 112.730 169.265 113.065 170.235 ;
        RECT 113.575 170.065 115.605 170.235 ;
        RECT 112.730 168.595 112.900 169.265 ;
        RECT 113.575 169.095 113.745 170.065 ;
        RECT 113.070 168.765 113.325 169.095 ;
        RECT 113.550 168.765 113.745 169.095 ;
        RECT 113.915 169.725 115.040 169.895 ;
        RECT 113.155 168.595 113.325 168.765 ;
        RECT 113.915 168.595 114.085 169.725 ;
        RECT 110.880 168.405 111.630 168.575 ;
        RECT 111.375 168.115 111.630 168.405 ;
        RECT 112.730 168.025 112.985 168.595 ;
        RECT 113.155 168.425 114.085 168.595 ;
        RECT 114.255 169.385 115.265 169.555 ;
        RECT 114.255 168.585 114.425 169.385 ;
        RECT 114.630 169.045 114.905 169.185 ;
        RECT 114.625 168.875 114.905 169.045 ;
        RECT 113.910 168.390 114.085 168.425 ;
        RECT 113.910 168.025 114.440 168.390 ;
        RECT 114.630 168.025 114.905 168.875 ;
        RECT 115.075 168.025 115.265 169.385 ;
        RECT 115.435 169.400 115.605 170.065 ;
        RECT 116.180 169.645 116.695 170.055 ;
        RECT 115.435 169.210 116.185 169.400 ;
        RECT 116.355 168.835 116.695 169.645 ;
        RECT 115.465 168.665 116.695 168.835 ;
        RECT 116.865 169.265 117.250 170.235 ;
        RECT 118.265 169.775 118.545 170.235 ;
        RECT 117.420 169.555 118.545 169.775 ;
        RECT 116.175 168.060 116.420 168.665 ;
        RECT 116.865 168.595 117.145 169.265 ;
        RECT 117.420 169.095 117.870 169.555 ;
        RECT 118.735 169.385 119.135 170.235 ;
        RECT 119.975 169.775 120.260 170.235 ;
        RECT 117.315 168.765 117.870 169.095 ;
        RECT 118.040 168.825 119.135 169.385 ;
        RECT 117.420 168.655 117.870 168.765 ;
        RECT 116.865 168.025 117.250 168.595 ;
        RECT 117.420 168.485 118.545 168.655 ;
        RECT 118.265 168.025 118.545 168.485 ;
        RECT 118.735 168.025 119.135 168.825 ;
        RECT 119.305 169.555 120.260 169.775 ;
        RECT 119.305 168.655 119.515 169.555 ;
        RECT 119.685 168.825 120.375 169.385 ;
        RECT 120.985 169.255 121.315 170.235 ;
        RECT 122.435 169.800 122.620 170.205 ;
        RECT 120.565 168.845 120.895 169.095 ;
        RECT 121.065 168.655 121.315 169.255 ;
        RECT 119.305 168.485 120.260 168.655 ;
        RECT 119.975 168.025 120.260 168.485 ;
        RECT 120.985 168.025 121.315 168.655 ;
        RECT 121.955 169.625 122.620 169.800 ;
        RECT 121.955 168.595 122.295 169.625 ;
        RECT 123.325 169.435 123.595 170.205 ;
        RECT 122.465 169.265 123.595 169.435 ;
        RECT 122.465 168.765 122.715 169.265 ;
        RECT 121.955 168.425 122.640 168.595 ;
        RECT 122.435 168.025 122.640 168.425 ;
        RECT 123.425 168.355 123.595 169.265 ;
        RECT 123.335 168.025 123.595 168.355 ;
        RECT 123.765 169.330 124.035 170.235 ;
        RECT 124.715 169.475 124.885 170.235 ;
        RECT 123.765 168.530 123.935 169.330 ;
        RECT 124.220 169.305 124.885 169.475 ;
        RECT 124.220 169.160 124.390 169.305 ;
        RECT 124.105 168.830 124.390 169.160 ;
        RECT 124.220 168.575 124.390 168.830 ;
        RECT 124.625 168.755 124.955 169.125 ;
        RECT 123.765 168.025 124.025 168.530 ;
        RECT 124.220 168.405 124.885 168.575 ;
        RECT 124.715 168.025 124.885 168.405 ;
        RECT 18.430 166.975 18.685 167.505 ;
        RECT 19.405 167.305 20.475 167.475 ;
        RECT 18.430 166.325 18.640 166.975 ;
        RECT 19.405 166.950 19.725 167.305 ;
        RECT 19.400 166.775 19.725 166.950 ;
        RECT 18.810 166.475 19.725 166.775 ;
        RECT 19.895 166.735 20.135 167.135 ;
        RECT 20.305 167.075 20.475 167.305 ;
        RECT 21.005 167.235 21.955 167.515 ;
        RECT 22.175 167.325 22.525 167.495 ;
        RECT 20.305 166.905 20.835 167.075 ;
        RECT 18.810 166.445 19.550 166.475 ;
        RECT 18.430 165.445 18.685 166.325 ;
        RECT 19.380 165.855 19.550 166.445 ;
        RECT 19.895 166.365 20.435 166.735 ;
        RECT 20.615 166.625 20.835 166.905 ;
        RECT 21.005 166.455 21.175 167.235 ;
        RECT 20.770 166.285 21.175 166.455 ;
        RECT 21.345 166.445 21.695 167.065 ;
        RECT 20.770 166.195 20.940 166.285 ;
        RECT 21.865 166.275 22.075 167.065 ;
        RECT 19.720 166.025 20.940 166.195 ;
        RECT 21.400 166.115 22.075 166.275 ;
        RECT 19.380 165.685 20.180 165.855 ;
        RECT 20.010 165.395 20.180 165.685 ;
        RECT 20.770 165.645 20.940 166.025 ;
        RECT 21.110 166.105 22.075 166.115 ;
        RECT 22.265 166.935 22.525 167.325 ;
        RECT 23.940 167.295 24.795 167.465 ;
        RECT 25.000 167.295 25.495 167.465 ;
        RECT 22.265 166.245 22.435 166.935 ;
        RECT 22.605 166.585 22.775 166.765 ;
        RECT 22.945 166.755 23.735 167.005 ;
        RECT 23.940 166.585 24.110 167.295 ;
        RECT 24.280 166.785 24.635 167.005 ;
        RECT 22.605 166.415 24.295 166.585 ;
        RECT 21.110 165.815 21.570 166.105 ;
        RECT 22.265 166.075 23.765 166.245 ;
        RECT 22.265 165.935 22.435 166.075 ;
        RECT 21.875 165.765 22.435 165.935 ;
        RECT 20.770 165.305 21.640 165.645 ;
        RECT 21.875 165.305 22.045 165.765 ;
        RECT 22.880 165.735 23.955 165.905 ;
        RECT 22.880 165.395 23.050 165.735 ;
        RECT 23.785 165.395 23.955 165.735 ;
        RECT 24.125 165.635 24.295 166.415 ;
        RECT 24.465 166.195 24.635 166.785 ;
        RECT 24.805 166.385 25.155 167.005 ;
        RECT 24.465 165.805 24.930 166.195 ;
        RECT 25.325 165.935 25.495 167.295 ;
        RECT 25.665 166.105 26.125 167.155 ;
        RECT 25.100 165.765 25.495 165.935 ;
        RECT 25.100 165.635 25.270 165.765 ;
        RECT 24.125 165.305 24.805 165.635 ;
        RECT 25.020 165.305 25.270 165.635 ;
        RECT 25.860 165.320 26.185 166.105 ;
        RECT 26.355 165.305 26.525 167.425 ;
        RECT 27.195 167.135 27.450 167.425 ;
        RECT 26.700 166.965 27.450 167.135 ;
        RECT 28.185 167.035 28.445 167.490 ;
        RECT 29.055 167.035 29.315 167.490 ;
        RECT 29.915 167.035 30.175 167.490 ;
        RECT 30.775 167.035 31.035 167.490 ;
        RECT 31.620 167.035 31.895 167.490 ;
        RECT 32.480 167.035 32.740 167.490 ;
        RECT 33.340 167.035 33.600 167.490 ;
        RECT 34.200 167.035 34.460 167.490 ;
        RECT 26.700 165.975 26.930 166.965 ;
        RECT 27.715 166.865 34.460 167.035 ;
        RECT 27.100 166.145 27.450 166.795 ;
        RECT 27.715 166.275 28.880 166.865 ;
        RECT 35.060 166.695 35.310 167.505 ;
        RECT 35.920 166.695 36.170 167.505 ;
        RECT 37.745 167.010 38.005 167.515 ;
        RECT 38.695 167.135 38.865 167.515 ;
        RECT 29.050 166.445 36.170 166.695 ;
        RECT 36.340 166.445 36.655 167.005 ;
        RECT 27.715 166.050 34.460 166.275 ;
        RECT 26.700 165.805 27.450 165.975 ;
        RECT 27.195 165.305 27.450 165.805 ;
        RECT 28.155 165.310 28.445 166.050 ;
        RECT 29.055 166.035 34.460 166.050 ;
        RECT 29.055 165.310 29.315 166.035 ;
        RECT 29.915 165.310 30.175 166.035 ;
        RECT 30.775 165.310 31.035 166.035 ;
        RECT 31.620 165.310 31.880 166.035 ;
        RECT 32.480 165.310 32.740 166.035 ;
        RECT 33.340 165.310 33.600 166.035 ;
        RECT 34.200 165.310 34.460 166.035 ;
        RECT 35.060 165.310 35.310 166.445 ;
        RECT 35.925 165.305 36.170 166.445 ;
        RECT 37.745 166.210 37.915 167.010 ;
        RECT 38.200 166.965 38.865 167.135 ;
        RECT 38.200 166.710 38.370 166.965 ;
        RECT 39.565 166.885 39.895 167.515 ;
        RECT 41.055 167.135 41.225 167.515 ;
        RECT 41.055 166.965 41.720 167.135 ;
        RECT 41.915 167.010 42.175 167.515 ;
        RECT 38.085 166.380 38.370 166.710 ;
        RECT 38.605 166.415 38.935 166.785 ;
        RECT 38.200 166.235 38.370 166.380 ;
        RECT 39.565 166.285 39.815 166.885 ;
        RECT 39.985 166.445 40.315 166.695 ;
        RECT 40.985 166.415 41.315 166.785 ;
        RECT 41.550 166.710 41.720 166.965 ;
        RECT 41.550 166.380 41.835 166.710 ;
        RECT 37.745 165.305 38.015 166.210 ;
        RECT 38.200 166.065 38.865 166.235 ;
        RECT 38.695 165.305 38.865 166.065 ;
        RECT 39.565 165.305 39.895 166.285 ;
        RECT 41.550 166.235 41.720 166.380 ;
        RECT 41.055 166.065 41.720 166.235 ;
        RECT 42.005 166.210 42.175 167.010 ;
        RECT 42.785 166.885 43.115 167.515 ;
        RECT 43.840 167.055 44.125 167.515 ;
        RECT 43.840 166.885 44.795 167.055 ;
        RECT 42.365 166.445 42.695 166.695 ;
        RECT 42.865 166.285 43.115 166.885 ;
        RECT 41.055 165.305 41.225 166.065 ;
        RECT 41.905 165.305 42.175 166.210 ;
        RECT 42.785 165.305 43.115 166.285 ;
        RECT 43.725 166.155 44.415 166.715 ;
        RECT 44.585 165.985 44.795 166.885 ;
        RECT 43.840 165.765 44.795 165.985 ;
        RECT 44.965 166.715 45.365 167.515 ;
        RECT 45.555 167.055 45.835 167.515 ;
        RECT 45.555 166.885 46.680 167.055 ;
        RECT 46.850 166.945 47.235 167.515 ;
        RECT 46.230 166.775 46.680 166.885 ;
        RECT 44.965 166.155 46.060 166.715 ;
        RECT 46.230 166.445 46.785 166.775 ;
        RECT 43.840 165.305 44.125 165.765 ;
        RECT 44.965 165.305 45.365 166.155 ;
        RECT 46.230 165.985 46.680 166.445 ;
        RECT 46.955 166.275 47.235 166.945 ;
        RECT 45.555 165.765 46.680 165.985 ;
        RECT 45.555 165.305 45.835 165.765 ;
        RECT 46.850 165.305 47.235 166.275 ;
        RECT 47.410 166.975 47.665 167.505 ;
        RECT 48.385 167.305 49.455 167.475 ;
        RECT 47.410 166.325 47.620 166.975 ;
        RECT 48.385 166.950 48.705 167.305 ;
        RECT 48.380 166.775 48.705 166.950 ;
        RECT 47.790 166.475 48.705 166.775 ;
        RECT 48.875 166.735 49.115 167.135 ;
        RECT 49.285 167.075 49.455 167.305 ;
        RECT 49.985 167.235 50.935 167.515 ;
        RECT 51.155 167.325 51.505 167.495 ;
        RECT 49.285 166.905 49.815 167.075 ;
        RECT 47.790 166.445 48.530 166.475 ;
        RECT 47.410 165.445 47.665 166.325 ;
        RECT 48.360 165.855 48.530 166.445 ;
        RECT 48.875 166.365 49.415 166.735 ;
        RECT 49.595 166.625 49.815 166.905 ;
        RECT 49.985 166.455 50.155 167.235 ;
        RECT 49.750 166.285 50.155 166.455 ;
        RECT 50.325 166.445 50.675 167.065 ;
        RECT 49.750 166.195 49.920 166.285 ;
        RECT 50.845 166.275 51.055 167.065 ;
        RECT 48.700 166.025 49.920 166.195 ;
        RECT 50.380 166.115 51.055 166.275 ;
        RECT 48.360 165.685 49.160 165.855 ;
        RECT 48.990 165.395 49.160 165.685 ;
        RECT 49.750 165.645 49.920 166.025 ;
        RECT 50.090 166.105 51.055 166.115 ;
        RECT 51.245 166.935 51.505 167.325 ;
        RECT 52.920 167.295 53.775 167.465 ;
        RECT 53.980 167.295 54.475 167.465 ;
        RECT 51.245 166.245 51.415 166.935 ;
        RECT 51.585 166.585 51.755 166.765 ;
        RECT 51.925 166.755 52.715 167.005 ;
        RECT 52.920 166.585 53.090 167.295 ;
        RECT 53.260 166.785 53.615 167.005 ;
        RECT 51.585 166.415 53.275 166.585 ;
        RECT 50.090 165.815 50.550 166.105 ;
        RECT 51.245 166.075 52.745 166.245 ;
        RECT 51.245 165.935 51.415 166.075 ;
        RECT 50.855 165.765 51.415 165.935 ;
        RECT 49.750 165.305 50.620 165.645 ;
        RECT 50.855 165.305 51.025 165.765 ;
        RECT 51.860 165.735 52.935 165.905 ;
        RECT 51.860 165.395 52.030 165.735 ;
        RECT 52.765 165.395 52.935 165.735 ;
        RECT 53.105 165.635 53.275 166.415 ;
        RECT 53.445 166.195 53.615 166.785 ;
        RECT 53.785 166.385 54.135 167.005 ;
        RECT 53.445 165.805 53.910 166.195 ;
        RECT 54.305 165.935 54.475 167.295 ;
        RECT 54.645 166.105 55.105 167.155 ;
        RECT 54.080 165.765 54.475 165.935 ;
        RECT 54.080 165.635 54.250 165.765 ;
        RECT 53.105 165.305 53.785 165.635 ;
        RECT 54.000 165.305 54.250 165.635 ;
        RECT 54.840 165.320 55.165 166.105 ;
        RECT 55.335 165.305 55.505 167.425 ;
        RECT 56.175 167.135 56.430 167.425 ;
        RECT 55.680 166.965 56.430 167.135 ;
        RECT 55.680 165.975 55.910 166.965 ;
        RECT 57.965 166.885 58.295 167.515 ;
        RECT 60.475 167.035 60.645 167.515 ;
        RECT 61.315 167.035 61.485 167.515 ;
        RECT 62.155 167.035 62.325 167.515 ;
        RECT 56.080 166.145 56.430 166.795 ;
        RECT 57.965 166.285 58.215 166.885 ;
        RECT 60.475 166.865 61.485 167.035 ;
        RECT 61.690 166.865 62.325 167.035 ;
        RECT 65.075 167.035 65.245 167.515 ;
        RECT 65.915 167.035 66.085 167.515 ;
        RECT 66.755 167.035 66.925 167.515 ;
        RECT 67.695 167.035 67.955 167.425 ;
        RECT 68.555 167.035 68.850 167.425 ;
        RECT 69.475 167.185 69.775 167.515 ;
        RECT 65.075 166.865 66.085 167.035 ;
        RECT 66.290 166.865 66.925 167.035 ;
        RECT 67.200 166.865 68.850 167.035 ;
        RECT 58.385 166.445 58.715 166.695 ;
        RECT 60.475 166.665 60.970 166.865 ;
        RECT 61.690 166.695 61.860 166.865 ;
        RECT 65.075 166.835 65.575 166.865 ;
        RECT 60.475 166.495 60.975 166.665 ;
        RECT 61.360 166.525 61.860 166.695 ;
        RECT 60.475 166.325 60.970 166.495 ;
        RECT 55.680 165.805 56.430 165.975 ;
        RECT 56.175 165.305 56.430 165.805 ;
        RECT 57.965 165.305 58.295 166.285 ;
        RECT 60.475 166.155 61.485 166.325 ;
        RECT 60.475 165.305 60.645 166.155 ;
        RECT 61.315 165.305 61.485 166.155 ;
        RECT 61.690 166.285 61.860 166.525 ;
        RECT 62.030 166.455 62.410 166.695 ;
        RECT 65.075 166.325 65.570 166.835 ;
        RECT 66.290 166.695 66.460 166.865 ;
        RECT 65.960 166.525 66.460 166.695 ;
        RECT 61.690 166.115 62.405 166.285 ;
        RECT 62.075 165.305 62.405 166.115 ;
        RECT 65.075 166.155 66.085 166.325 ;
        RECT 65.075 165.305 65.245 166.155 ;
        RECT 65.915 165.305 66.085 166.155 ;
        RECT 66.290 166.285 66.460 166.525 ;
        RECT 66.630 166.455 67.010 166.695 ;
        RECT 67.200 166.355 67.605 166.865 ;
        RECT 67.775 166.525 68.915 166.695 ;
        RECT 66.290 166.115 67.005 166.285 ;
        RECT 67.200 166.185 67.955 166.355 ;
        RECT 66.675 165.305 67.005 166.115 ;
        RECT 67.695 165.935 67.955 166.185 ;
        RECT 68.745 166.275 68.915 166.525 ;
        RECT 69.085 166.445 69.435 167.015 ;
        RECT 69.605 166.275 69.775 167.185 ;
        RECT 71.335 167.155 71.665 167.515 ;
        RECT 72.365 167.155 72.695 167.515 ;
        RECT 71.335 166.945 72.695 167.155 ;
        RECT 73.205 166.925 73.915 167.515 ;
        RECT 71.325 166.445 71.635 166.775 ;
        RECT 71.845 166.445 72.220 166.775 ;
        RECT 72.540 166.445 73.035 166.775 ;
        RECT 68.745 166.105 69.775 166.275 ;
        RECT 67.695 165.765 68.815 165.935 ;
        RECT 67.695 165.305 67.955 165.765 ;
        RECT 68.555 165.305 68.815 165.765 ;
        RECT 69.465 165.305 69.775 166.105 ;
        RECT 71.845 165.520 72.015 166.445 ;
        RECT 72.185 165.955 72.515 166.175 ;
        RECT 72.710 166.155 73.035 166.445 ;
        RECT 73.210 166.155 73.540 166.695 ;
        RECT 73.710 165.955 73.915 166.925 ;
        RECT 72.185 165.725 73.915 165.955 ;
        RECT 72.185 165.325 72.515 165.725 ;
        RECT 73.215 165.305 73.915 165.725 ;
        RECT 75.840 166.975 76.095 167.505 ;
        RECT 75.840 166.115 76.020 166.975 ;
        RECT 76.740 166.775 76.990 167.425 ;
        RECT 76.190 166.445 76.990 166.775 ;
        RECT 75.840 165.645 76.095 166.115 ;
        RECT 75.755 165.475 76.095 165.645 ;
        RECT 75.840 165.445 76.095 165.475 ;
        RECT 76.740 165.855 76.990 166.445 ;
        RECT 77.190 167.090 77.510 167.420 ;
        RECT 78.550 167.295 79.400 167.465 ;
        RECT 77.190 166.195 77.380 167.090 ;
        RECT 77.700 166.765 78.360 167.035 ;
        RECT 78.030 166.705 78.360 166.765 ;
        RECT 77.550 166.535 77.880 166.595 ;
        RECT 78.550 166.535 78.720 167.295 ;
        RECT 80.480 167.045 80.730 167.475 ;
        RECT 78.890 166.875 80.140 167.045 ;
        RECT 78.890 166.755 79.220 166.875 ;
        RECT 77.550 166.365 79.450 166.535 ;
        RECT 77.190 166.025 79.110 166.195 ;
        RECT 77.190 166.005 77.510 166.025 ;
        RECT 76.740 165.345 77.070 165.855 ;
        RECT 77.340 165.395 77.510 166.005 ;
        RECT 79.280 165.855 79.450 166.365 ;
        RECT 79.620 166.295 79.800 166.705 ;
        RECT 79.970 166.115 80.140 166.875 ;
        RECT 78.240 165.685 79.450 165.855 ;
        RECT 79.620 165.805 80.140 166.115 ;
        RECT 80.310 166.705 80.730 167.045 ;
        RECT 81.600 167.305 82.615 167.505 ;
        RECT 81.020 166.705 81.430 167.035 ;
        RECT 80.310 165.935 80.500 166.705 ;
        RECT 81.600 166.575 81.770 167.305 ;
        RECT 82.915 167.135 83.085 167.465 ;
        RECT 81.940 166.755 82.290 167.125 ;
        RECT 81.600 166.535 82.020 166.575 ;
        RECT 80.670 166.365 82.020 166.535 ;
        RECT 80.670 166.205 80.920 166.365 ;
        RECT 81.430 165.935 81.680 166.195 ;
        RECT 80.310 165.685 81.680 165.935 ;
        RECT 78.240 165.395 78.480 165.685 ;
        RECT 79.280 165.605 79.450 165.685 ;
        RECT 79.280 165.355 79.910 165.605 ;
        RECT 80.880 165.395 81.050 165.685 ;
        RECT 81.850 165.520 82.020 166.365 ;
        RECT 82.470 166.195 82.690 167.065 ;
        RECT 82.915 166.945 83.610 167.135 ;
        RECT 82.190 165.815 82.690 166.195 ;
        RECT 82.860 166.145 83.270 166.765 ;
        RECT 83.440 165.975 83.610 166.945 ;
        RECT 82.915 165.805 83.610 165.975 ;
        RECT 81.850 165.350 82.680 165.520 ;
        RECT 82.915 165.305 83.085 165.805 ;
        RECT 83.800 165.305 84.025 167.425 ;
        RECT 84.695 167.135 84.865 167.425 ;
        RECT 84.200 166.965 84.865 167.135 ;
        RECT 84.200 165.975 84.430 166.965 ;
        RECT 85.565 166.885 85.895 167.515 ;
        RECT 86.945 166.885 87.275 167.515 ;
        RECT 97.460 166.975 97.715 167.505 ;
        RECT 84.600 166.145 84.950 166.795 ;
        RECT 85.565 166.285 85.815 166.885 ;
        RECT 85.985 166.445 86.315 166.695 ;
        RECT 86.945 166.285 87.195 166.885 ;
        RECT 87.365 166.445 87.695 166.695 ;
        RECT 84.200 165.805 84.865 165.975 ;
        RECT 84.695 165.305 84.865 165.805 ;
        RECT 85.565 165.305 85.895 166.285 ;
        RECT 86.945 165.305 87.275 166.285 ;
        RECT 97.460 166.115 97.640 166.975 ;
        RECT 98.360 166.775 98.610 167.425 ;
        RECT 97.810 166.445 98.610 166.775 ;
        RECT 97.460 165.645 97.715 166.115 ;
        RECT 97.375 165.475 97.715 165.645 ;
        RECT 97.460 165.445 97.715 165.475 ;
        RECT 98.360 165.855 98.610 166.445 ;
        RECT 98.810 167.090 99.130 167.420 ;
        RECT 100.170 167.295 101.020 167.465 ;
        RECT 98.810 166.195 99.000 167.090 ;
        RECT 99.320 166.765 99.980 167.035 ;
        RECT 99.650 166.705 99.980 166.765 ;
        RECT 99.170 166.535 99.500 166.595 ;
        RECT 100.170 166.535 100.340 167.295 ;
        RECT 102.100 167.045 102.350 167.475 ;
        RECT 100.510 166.875 101.760 167.045 ;
        RECT 100.510 166.755 100.840 166.875 ;
        RECT 99.170 166.365 101.070 166.535 ;
        RECT 98.810 166.025 100.730 166.195 ;
        RECT 98.810 166.005 99.130 166.025 ;
        RECT 98.360 165.345 98.690 165.855 ;
        RECT 98.960 165.395 99.130 166.005 ;
        RECT 100.900 165.855 101.070 166.365 ;
        RECT 101.240 166.295 101.420 166.705 ;
        RECT 101.590 166.115 101.760 166.875 ;
        RECT 99.860 165.685 101.070 165.855 ;
        RECT 101.240 165.805 101.760 166.115 ;
        RECT 101.930 166.705 102.350 167.045 ;
        RECT 103.220 167.305 104.235 167.505 ;
        RECT 102.640 166.705 103.050 167.035 ;
        RECT 101.930 165.935 102.120 166.705 ;
        RECT 103.220 166.575 103.390 167.305 ;
        RECT 104.535 167.135 104.705 167.465 ;
        RECT 103.560 166.755 103.910 167.125 ;
        RECT 103.220 166.535 103.640 166.575 ;
        RECT 102.290 166.365 103.640 166.535 ;
        RECT 102.290 166.205 102.540 166.365 ;
        RECT 103.050 165.935 103.300 166.195 ;
        RECT 101.930 165.685 103.300 165.935 ;
        RECT 99.860 165.395 100.100 165.685 ;
        RECT 100.900 165.605 101.070 165.685 ;
        RECT 100.900 165.355 101.530 165.605 ;
        RECT 102.500 165.395 102.670 165.685 ;
        RECT 103.470 165.520 103.640 166.365 ;
        RECT 104.090 166.195 104.310 167.065 ;
        RECT 104.535 166.945 105.230 167.135 ;
        RECT 103.810 165.815 104.310 166.195 ;
        RECT 104.480 166.145 104.890 166.765 ;
        RECT 105.060 165.975 105.230 166.945 ;
        RECT 104.535 165.805 105.230 165.975 ;
        RECT 103.470 165.350 104.300 165.520 ;
        RECT 104.535 165.305 104.705 165.805 ;
        RECT 105.420 165.305 105.645 167.425 ;
        RECT 106.315 167.135 106.485 167.425 ;
        RECT 105.820 166.965 106.485 167.135 ;
        RECT 107.320 167.055 107.605 167.515 ;
        RECT 105.820 165.975 106.050 166.965 ;
        RECT 107.320 166.885 108.275 167.055 ;
        RECT 106.220 166.145 106.570 166.795 ;
        RECT 107.205 166.155 107.895 166.715 ;
        RECT 108.065 165.985 108.275 166.885 ;
        RECT 105.820 165.805 106.485 165.975 ;
        RECT 106.315 165.305 106.485 165.805 ;
        RECT 107.320 165.765 108.275 165.985 ;
        RECT 108.445 166.715 108.845 167.515 ;
        RECT 109.035 167.055 109.315 167.515 ;
        RECT 109.035 166.885 110.160 167.055 ;
        RECT 110.330 166.945 110.715 167.515 ;
        RECT 109.710 166.775 110.160 166.885 ;
        RECT 108.445 166.155 109.540 166.715 ;
        RECT 109.710 166.445 110.265 166.775 ;
        RECT 107.320 165.305 107.605 165.765 ;
        RECT 108.445 165.305 108.845 166.155 ;
        RECT 109.710 165.985 110.160 166.445 ;
        RECT 110.435 166.275 110.715 166.945 ;
        RECT 109.035 165.765 110.160 165.985 ;
        RECT 109.035 165.305 109.315 165.765 ;
        RECT 110.330 165.305 110.715 166.275 ;
        RECT 110.885 166.945 111.270 167.515 ;
        RECT 112.285 167.055 112.565 167.515 ;
        RECT 110.885 166.275 111.165 166.945 ;
        RECT 111.440 166.885 112.565 167.055 ;
        RECT 111.440 166.775 111.890 166.885 ;
        RECT 111.335 166.445 111.890 166.775 ;
        RECT 112.755 166.715 113.155 167.515 ;
        RECT 113.995 167.055 114.280 167.515 ;
        RECT 110.885 165.305 111.270 166.275 ;
        RECT 111.440 165.985 111.890 166.445 ;
        RECT 112.060 166.155 113.155 166.715 ;
        RECT 111.440 165.765 112.565 165.985 ;
        RECT 112.285 165.305 112.565 165.765 ;
        RECT 112.755 165.305 113.155 166.155 ;
        RECT 113.325 166.885 114.280 167.055 ;
        RECT 115.950 166.975 116.205 167.505 ;
        RECT 116.925 167.305 117.995 167.475 ;
        RECT 113.325 165.985 113.535 166.885 ;
        RECT 113.705 166.155 114.395 166.715 ;
        RECT 115.950 166.325 116.160 166.975 ;
        RECT 116.925 166.950 117.245 167.305 ;
        RECT 116.920 166.775 117.245 166.950 ;
        RECT 116.330 166.475 117.245 166.775 ;
        RECT 117.415 166.735 117.655 167.135 ;
        RECT 117.825 167.075 117.995 167.305 ;
        RECT 118.525 167.235 119.475 167.515 ;
        RECT 119.695 167.325 120.045 167.495 ;
        RECT 117.825 166.905 118.355 167.075 ;
        RECT 116.330 166.445 117.070 166.475 ;
        RECT 113.325 165.765 114.280 165.985 ;
        RECT 113.995 165.305 114.280 165.765 ;
        RECT 115.950 165.445 116.205 166.325 ;
        RECT 116.900 165.855 117.070 166.445 ;
        RECT 117.415 166.365 117.955 166.735 ;
        RECT 118.135 166.625 118.355 166.905 ;
        RECT 118.525 166.455 118.695 167.235 ;
        RECT 118.290 166.285 118.695 166.455 ;
        RECT 118.865 166.445 119.215 167.065 ;
        RECT 118.290 166.195 118.460 166.285 ;
        RECT 119.385 166.275 119.595 167.065 ;
        RECT 117.240 166.025 118.460 166.195 ;
        RECT 118.920 166.115 119.595 166.275 ;
        RECT 116.900 165.685 117.700 165.855 ;
        RECT 117.530 165.395 117.700 165.685 ;
        RECT 118.290 165.645 118.460 166.025 ;
        RECT 118.630 166.105 119.595 166.115 ;
        RECT 119.785 166.935 120.045 167.325 ;
        RECT 121.460 167.295 122.315 167.465 ;
        RECT 122.520 167.295 123.015 167.465 ;
        RECT 119.785 166.245 119.955 166.935 ;
        RECT 120.125 166.585 120.295 166.765 ;
        RECT 120.465 166.755 121.255 167.005 ;
        RECT 121.460 166.585 121.630 167.295 ;
        RECT 121.800 166.785 122.155 167.005 ;
        RECT 120.125 166.415 121.815 166.585 ;
        RECT 118.630 165.815 119.090 166.105 ;
        RECT 119.785 166.075 121.285 166.245 ;
        RECT 119.785 165.935 119.955 166.075 ;
        RECT 119.395 165.765 119.955 165.935 ;
        RECT 118.290 165.305 119.160 165.645 ;
        RECT 119.395 165.305 119.565 165.765 ;
        RECT 120.400 165.735 121.475 165.905 ;
        RECT 120.400 165.395 120.570 165.735 ;
        RECT 121.305 165.395 121.475 165.735 ;
        RECT 121.645 165.635 121.815 166.415 ;
        RECT 121.985 166.195 122.155 166.785 ;
        RECT 122.325 166.385 122.675 167.005 ;
        RECT 121.985 165.805 122.450 166.195 ;
        RECT 122.845 165.935 123.015 167.295 ;
        RECT 123.185 166.105 123.645 167.155 ;
        RECT 122.620 165.765 123.015 165.935 ;
        RECT 122.620 165.635 122.790 165.765 ;
        RECT 121.645 165.305 122.325 165.635 ;
        RECT 122.540 165.305 122.790 165.635 ;
        RECT 123.380 165.320 123.705 166.105 ;
        RECT 123.875 165.305 124.045 167.425 ;
        RECT 124.715 167.135 124.970 167.425 ;
        RECT 124.220 166.965 124.970 167.135 ;
        RECT 124.220 165.975 124.450 166.965 ;
        RECT 124.620 166.145 124.970 166.795 ;
        RECT 124.220 165.805 124.970 165.975 ;
        RECT 124.715 165.305 124.970 165.805 ;
        RECT 25.785 163.890 26.055 164.795 ;
        RECT 26.735 164.035 26.905 164.795 ;
        RECT 25.785 163.090 25.955 163.890 ;
        RECT 26.240 163.865 26.905 164.035 ;
        RECT 26.240 163.720 26.410 163.865 ;
        RECT 26.125 163.390 26.410 163.720 ;
        RECT 27.170 163.775 27.425 164.655 ;
        RECT 28.750 164.415 28.920 164.705 ;
        RECT 28.120 164.245 28.920 164.415 ;
        RECT 29.510 164.455 30.380 164.795 ;
        RECT 26.240 163.135 26.410 163.390 ;
        RECT 26.645 163.315 26.975 163.685 ;
        RECT 25.785 162.585 26.045 163.090 ;
        RECT 26.240 162.965 26.905 163.135 ;
        RECT 26.735 162.585 26.905 162.965 ;
        RECT 27.170 163.125 27.380 163.775 ;
        RECT 28.120 163.655 28.290 164.245 ;
        RECT 29.510 164.075 29.680 164.455 ;
        RECT 30.615 164.335 30.785 164.795 ;
        RECT 31.620 164.365 31.790 164.705 ;
        RECT 32.525 164.365 32.695 164.705 ;
        RECT 28.460 163.905 29.680 164.075 ;
        RECT 29.850 163.995 30.310 164.285 ;
        RECT 30.615 164.165 31.175 164.335 ;
        RECT 31.620 164.195 32.695 164.365 ;
        RECT 32.865 164.465 33.545 164.795 ;
        RECT 33.760 164.465 34.010 164.795 ;
        RECT 31.005 164.025 31.175 164.165 ;
        RECT 29.850 163.985 30.815 163.995 ;
        RECT 29.510 163.815 29.680 163.905 ;
        RECT 30.140 163.825 30.815 163.985 ;
        RECT 27.550 163.625 28.290 163.655 ;
        RECT 27.550 163.325 28.465 163.625 ;
        RECT 28.140 163.150 28.465 163.325 ;
        RECT 27.170 162.595 27.425 163.125 ;
        RECT 28.145 162.795 28.465 163.150 ;
        RECT 28.635 163.365 29.175 163.735 ;
        RECT 29.510 163.645 29.915 163.815 ;
        RECT 28.635 162.965 28.875 163.365 ;
        RECT 29.355 163.195 29.575 163.475 ;
        RECT 29.045 163.025 29.575 163.195 ;
        RECT 29.045 162.795 29.215 163.025 ;
        RECT 28.145 162.625 29.215 162.795 ;
        RECT 29.745 162.865 29.915 163.645 ;
        RECT 30.085 163.035 30.435 163.655 ;
        RECT 30.605 163.035 30.815 163.825 ;
        RECT 31.005 163.855 32.505 164.025 ;
        RECT 31.005 163.165 31.175 163.855 ;
        RECT 32.865 163.685 33.035 164.465 ;
        RECT 33.840 164.335 34.010 164.465 ;
        RECT 31.345 163.515 33.035 163.685 ;
        RECT 33.205 163.905 33.670 164.295 ;
        RECT 33.840 164.165 34.235 164.335 ;
        RECT 31.345 163.335 31.515 163.515 ;
        RECT 29.745 162.585 30.695 162.865 ;
        RECT 31.005 162.775 31.265 163.165 ;
        RECT 31.685 163.095 32.475 163.345 ;
        RECT 30.915 162.605 31.265 162.775 ;
        RECT 32.680 162.805 32.850 163.515 ;
        RECT 33.205 163.315 33.375 163.905 ;
        RECT 33.020 163.095 33.375 163.315 ;
        RECT 33.545 163.095 33.895 163.715 ;
        RECT 34.065 162.805 34.235 164.165 ;
        RECT 34.600 163.995 34.925 164.780 ;
        RECT 34.405 162.945 34.865 163.995 ;
        RECT 32.680 162.635 33.535 162.805 ;
        RECT 33.740 162.635 34.235 162.805 ;
        RECT 35.095 162.675 35.265 164.795 ;
        RECT 35.935 164.295 36.190 164.795 ;
        RECT 35.440 164.125 36.190 164.295 ;
        RECT 35.440 163.135 35.670 164.125 ;
        RECT 35.840 163.305 36.190 163.955 ;
        RECT 36.370 163.775 36.625 164.655 ;
        RECT 37.950 164.415 38.120 164.705 ;
        RECT 37.320 164.245 38.120 164.415 ;
        RECT 38.710 164.455 39.580 164.795 ;
        RECT 35.440 162.965 36.190 163.135 ;
        RECT 35.935 162.675 36.190 162.965 ;
        RECT 36.370 163.125 36.580 163.775 ;
        RECT 37.320 163.655 37.490 164.245 ;
        RECT 38.710 164.075 38.880 164.455 ;
        RECT 39.815 164.335 39.985 164.795 ;
        RECT 40.820 164.365 40.990 164.705 ;
        RECT 41.725 164.365 41.895 164.705 ;
        RECT 37.660 163.905 38.880 164.075 ;
        RECT 39.050 163.995 39.510 164.285 ;
        RECT 39.815 164.165 40.375 164.335 ;
        RECT 40.820 164.195 41.895 164.365 ;
        RECT 42.065 164.465 42.745 164.795 ;
        RECT 42.960 164.465 43.210 164.795 ;
        RECT 40.205 164.025 40.375 164.165 ;
        RECT 39.050 163.985 40.015 163.995 ;
        RECT 38.710 163.815 38.880 163.905 ;
        RECT 39.340 163.825 40.015 163.985 ;
        RECT 36.750 163.625 37.490 163.655 ;
        RECT 36.750 163.325 37.665 163.625 ;
        RECT 37.340 163.150 37.665 163.325 ;
        RECT 36.370 162.595 36.625 163.125 ;
        RECT 37.345 162.795 37.665 163.150 ;
        RECT 37.835 163.365 38.375 163.735 ;
        RECT 38.710 163.645 39.115 163.815 ;
        RECT 37.835 162.965 38.075 163.365 ;
        RECT 38.555 163.195 38.775 163.475 ;
        RECT 38.245 163.025 38.775 163.195 ;
        RECT 38.245 162.795 38.415 163.025 ;
        RECT 37.345 162.625 38.415 162.795 ;
        RECT 38.945 162.865 39.115 163.645 ;
        RECT 39.285 163.035 39.635 163.655 ;
        RECT 39.805 163.035 40.015 163.825 ;
        RECT 40.205 163.855 41.705 164.025 ;
        RECT 40.205 163.165 40.375 163.855 ;
        RECT 42.065 163.685 42.235 164.465 ;
        RECT 43.040 164.335 43.210 164.465 ;
        RECT 40.545 163.515 42.235 163.685 ;
        RECT 42.405 163.905 42.870 164.295 ;
        RECT 43.040 164.165 43.435 164.335 ;
        RECT 40.545 163.335 40.715 163.515 ;
        RECT 38.945 162.585 39.895 162.865 ;
        RECT 40.205 162.775 40.465 163.165 ;
        RECT 40.885 163.095 41.675 163.345 ;
        RECT 40.115 162.605 40.465 162.775 ;
        RECT 41.880 162.805 42.050 163.515 ;
        RECT 42.405 163.315 42.575 163.905 ;
        RECT 42.220 163.095 42.575 163.315 ;
        RECT 42.745 163.095 43.095 163.715 ;
        RECT 43.265 162.805 43.435 164.165 ;
        RECT 43.800 163.995 44.125 164.780 ;
        RECT 43.605 162.945 44.065 163.995 ;
        RECT 41.880 162.635 42.735 162.805 ;
        RECT 42.940 162.635 43.435 162.805 ;
        RECT 44.295 162.675 44.465 164.795 ;
        RECT 45.135 164.295 45.390 164.795 ;
        RECT 44.640 164.125 45.390 164.295 ;
        RECT 44.640 163.135 44.870 164.125 ;
        RECT 45.040 163.305 45.390 163.955 ;
        RECT 45.570 163.825 45.905 164.795 ;
        RECT 46.415 164.625 48.445 164.795 ;
        RECT 45.570 163.155 45.740 163.825 ;
        RECT 46.415 163.655 46.585 164.625 ;
        RECT 45.910 163.325 46.165 163.655 ;
        RECT 46.390 163.325 46.585 163.655 ;
        RECT 46.755 164.285 47.880 164.455 ;
        RECT 45.995 163.155 46.165 163.325 ;
        RECT 46.755 163.155 46.925 164.285 ;
        RECT 44.640 162.965 45.390 163.135 ;
        RECT 45.135 162.675 45.390 162.965 ;
        RECT 45.570 162.585 45.825 163.155 ;
        RECT 45.995 162.985 46.925 163.155 ;
        RECT 47.095 163.945 48.105 164.115 ;
        RECT 47.095 163.145 47.265 163.945 ;
        RECT 47.470 163.605 47.745 163.745 ;
        RECT 47.465 163.435 47.745 163.605 ;
        RECT 46.750 162.950 46.925 162.985 ;
        RECT 46.750 162.585 47.280 162.950 ;
        RECT 47.470 162.585 47.745 163.435 ;
        RECT 47.915 162.585 48.105 163.945 ;
        RECT 48.275 163.960 48.445 164.625 ;
        RECT 51.715 164.625 53.745 164.795 ;
        RECT 49.020 164.205 49.535 164.615 ;
        RECT 48.275 163.770 49.025 163.960 ;
        RECT 49.195 163.395 49.535 164.205 ;
        RECT 48.305 163.225 49.535 163.395 ;
        RECT 50.625 164.205 51.140 164.615 ;
        RECT 50.625 163.395 50.965 164.205 ;
        RECT 51.715 163.960 51.885 164.625 ;
        RECT 52.280 164.285 53.405 164.455 ;
        RECT 51.135 163.770 51.885 163.960 ;
        RECT 52.055 163.945 53.065 164.115 ;
        RECT 50.625 163.225 51.855 163.395 ;
        RECT 49.015 162.620 49.260 163.225 ;
        RECT 50.900 162.620 51.145 163.225 ;
        RECT 52.055 162.585 52.245 163.945 ;
        RECT 52.415 163.605 52.690 163.745 ;
        RECT 52.415 163.435 52.695 163.605 ;
        RECT 52.415 162.585 52.690 163.435 ;
        RECT 52.895 163.145 53.065 163.945 ;
        RECT 53.235 163.155 53.405 164.285 ;
        RECT 53.575 163.655 53.745 164.625 ;
        RECT 54.255 163.825 54.590 164.795 ;
        RECT 53.575 163.325 53.770 163.655 ;
        RECT 53.995 163.325 54.250 163.655 ;
        RECT 53.995 163.155 54.165 163.325 ;
        RECT 54.420 163.155 54.590 163.825 ;
        RECT 53.235 162.985 54.165 163.155 ;
        RECT 53.235 162.950 53.410 162.985 ;
        RECT 52.880 162.585 53.410 162.950 ;
        RECT 54.335 162.585 54.590 163.155 ;
        RECT 54.770 163.775 55.025 164.655 ;
        RECT 56.350 164.415 56.520 164.705 ;
        RECT 55.720 164.245 56.520 164.415 ;
        RECT 57.110 164.455 57.980 164.795 ;
        RECT 54.770 163.125 54.980 163.775 ;
        RECT 55.720 163.655 55.890 164.245 ;
        RECT 57.110 164.075 57.280 164.455 ;
        RECT 58.215 164.335 58.385 164.795 ;
        RECT 59.220 164.365 59.390 164.705 ;
        RECT 60.125 164.365 60.295 164.705 ;
        RECT 56.060 163.905 57.280 164.075 ;
        RECT 57.450 163.995 57.910 164.285 ;
        RECT 58.215 164.165 58.775 164.335 ;
        RECT 59.220 164.195 60.295 164.365 ;
        RECT 60.465 164.465 61.145 164.795 ;
        RECT 61.360 164.465 61.610 164.795 ;
        RECT 58.605 164.025 58.775 164.165 ;
        RECT 57.450 163.985 58.415 163.995 ;
        RECT 57.110 163.815 57.280 163.905 ;
        RECT 57.740 163.825 58.415 163.985 ;
        RECT 55.150 163.625 55.890 163.655 ;
        RECT 55.150 163.325 56.065 163.625 ;
        RECT 55.740 163.150 56.065 163.325 ;
        RECT 54.770 162.595 55.025 163.125 ;
        RECT 55.745 162.795 56.065 163.150 ;
        RECT 56.235 163.365 56.775 163.735 ;
        RECT 57.110 163.645 57.515 163.815 ;
        RECT 56.235 162.965 56.475 163.365 ;
        RECT 56.955 163.195 57.175 163.475 ;
        RECT 56.645 163.025 57.175 163.195 ;
        RECT 56.645 162.795 56.815 163.025 ;
        RECT 55.745 162.625 56.815 162.795 ;
        RECT 57.345 162.865 57.515 163.645 ;
        RECT 57.685 163.035 58.035 163.655 ;
        RECT 58.205 163.035 58.415 163.825 ;
        RECT 58.605 163.855 60.105 164.025 ;
        RECT 58.605 163.165 58.775 163.855 ;
        RECT 60.465 163.685 60.635 164.465 ;
        RECT 61.440 164.335 61.610 164.465 ;
        RECT 58.945 163.515 60.635 163.685 ;
        RECT 60.805 163.905 61.270 164.295 ;
        RECT 61.440 164.165 61.835 164.335 ;
        RECT 58.945 163.335 59.115 163.515 ;
        RECT 57.345 162.585 58.295 162.865 ;
        RECT 58.605 162.775 58.865 163.165 ;
        RECT 59.285 163.095 60.075 163.345 ;
        RECT 58.515 162.605 58.865 162.775 ;
        RECT 60.280 162.805 60.450 163.515 ;
        RECT 60.805 163.315 60.975 163.905 ;
        RECT 60.620 163.095 60.975 163.315 ;
        RECT 61.145 163.095 61.495 163.715 ;
        RECT 61.665 162.805 61.835 164.165 ;
        RECT 62.200 163.995 62.525 164.780 ;
        RECT 62.005 162.945 62.465 163.995 ;
        RECT 60.280 162.635 61.135 162.805 ;
        RECT 61.340 162.635 61.835 162.805 ;
        RECT 62.695 162.675 62.865 164.795 ;
        RECT 63.535 164.295 63.790 164.795 ;
        RECT 63.040 164.125 63.790 164.295 ;
        RECT 67.695 164.335 67.955 164.795 ;
        RECT 68.555 164.335 68.815 164.795 ;
        RECT 67.695 164.165 68.815 164.335 ;
        RECT 63.040 163.135 63.270 164.125 ;
        RECT 63.440 163.305 63.790 163.955 ;
        RECT 67.695 163.915 67.955 164.165 ;
        RECT 69.465 163.995 69.775 164.795 ;
        RECT 79.315 164.625 81.345 164.795 ;
        RECT 67.200 163.745 67.955 163.915 ;
        RECT 68.745 163.825 69.775 163.995 ;
        RECT 67.200 163.235 67.605 163.745 ;
        RECT 68.745 163.575 68.915 163.825 ;
        RECT 67.775 163.405 68.915 163.575 ;
        RECT 63.040 162.965 63.790 163.135 ;
        RECT 67.200 163.065 68.850 163.235 ;
        RECT 69.085 163.085 69.435 163.655 ;
        RECT 63.535 162.675 63.790 162.965 ;
        RECT 67.695 162.675 67.955 163.065 ;
        RECT 68.555 162.675 68.850 163.065 ;
        RECT 69.605 162.915 69.775 163.825 ;
        RECT 78.225 164.205 78.740 164.615 ;
        RECT 78.225 163.395 78.565 164.205 ;
        RECT 79.315 163.960 79.485 164.625 ;
        RECT 79.880 164.285 81.005 164.455 ;
        RECT 78.735 163.770 79.485 163.960 ;
        RECT 79.655 163.945 80.665 164.115 ;
        RECT 78.225 163.225 79.455 163.395 ;
        RECT 69.475 162.585 69.775 162.915 ;
        RECT 78.500 162.620 78.745 163.225 ;
        RECT 79.655 162.585 79.845 163.945 ;
        RECT 80.015 162.925 80.290 163.745 ;
        RECT 80.495 163.145 80.665 163.945 ;
        RECT 80.835 163.155 81.005 164.285 ;
        RECT 81.175 163.655 81.345 164.625 ;
        RECT 81.855 163.825 82.190 164.795 ;
        RECT 82.455 164.035 82.625 164.795 ;
        RECT 82.455 163.865 83.120 164.035 ;
        RECT 83.305 163.890 83.575 164.795 ;
        RECT 81.175 163.325 81.370 163.655 ;
        RECT 81.595 163.325 81.850 163.655 ;
        RECT 81.595 163.155 81.765 163.325 ;
        RECT 82.020 163.155 82.190 163.825 ;
        RECT 82.950 163.720 83.120 163.865 ;
        RECT 82.385 163.315 82.715 163.685 ;
        RECT 82.950 163.390 83.235 163.720 ;
        RECT 80.835 162.985 81.765 163.155 ;
        RECT 80.835 162.950 81.010 162.985 ;
        RECT 80.015 162.755 80.295 162.925 ;
        RECT 80.015 162.585 80.290 162.755 ;
        RECT 80.480 162.585 81.010 162.950 ;
        RECT 81.935 162.585 82.190 163.155 ;
        RECT 82.950 163.135 83.120 163.390 ;
        RECT 82.455 162.965 83.120 163.135 ;
        RECT 83.405 163.090 83.575 163.890 ;
        RECT 85.675 164.035 85.845 164.795 ;
        RECT 85.675 163.865 86.340 164.035 ;
        RECT 86.525 163.890 86.795 164.795 ;
        RECT 94.495 164.625 96.525 164.795 ;
        RECT 86.170 163.720 86.340 163.865 ;
        RECT 85.605 163.315 85.935 163.685 ;
        RECT 86.170 163.390 86.455 163.720 ;
        RECT 86.170 163.135 86.340 163.390 ;
        RECT 82.455 162.585 82.625 162.965 ;
        RECT 83.315 162.585 83.575 163.090 ;
        RECT 85.675 162.965 86.340 163.135 ;
        RECT 86.625 163.090 86.795 163.890 ;
        RECT 93.405 164.205 93.920 164.615 ;
        RECT 93.405 163.395 93.745 164.205 ;
        RECT 94.495 163.960 94.665 164.625 ;
        RECT 95.060 164.285 96.185 164.455 ;
        RECT 93.915 163.770 94.665 163.960 ;
        RECT 94.835 163.945 95.845 164.115 ;
        RECT 93.405 163.225 94.635 163.395 ;
        RECT 85.675 162.585 85.845 162.965 ;
        RECT 86.535 162.585 86.795 163.090 ;
        RECT 93.680 162.620 93.925 163.225 ;
        RECT 94.835 162.585 95.025 163.945 ;
        RECT 95.195 163.265 95.470 163.745 ;
        RECT 95.195 163.095 95.475 163.265 ;
        RECT 95.675 163.145 95.845 163.945 ;
        RECT 96.015 163.155 96.185 164.285 ;
        RECT 96.355 163.655 96.525 164.625 ;
        RECT 97.035 163.825 97.370 164.795 ;
        RECT 98.635 164.625 100.665 164.795 ;
        RECT 96.355 163.325 96.550 163.655 ;
        RECT 96.775 163.325 97.030 163.655 ;
        RECT 96.775 163.155 96.945 163.325 ;
        RECT 97.200 163.155 97.370 163.825 ;
        RECT 97.545 164.205 98.060 164.615 ;
        RECT 97.545 163.395 97.885 164.205 ;
        RECT 98.635 163.960 98.805 164.625 ;
        RECT 99.200 164.285 100.325 164.455 ;
        RECT 98.055 163.770 98.805 163.960 ;
        RECT 98.975 163.945 99.985 164.115 ;
        RECT 97.545 163.225 98.775 163.395 ;
        RECT 95.195 162.585 95.470 163.095 ;
        RECT 96.015 162.985 96.945 163.155 ;
        RECT 96.015 162.950 96.190 162.985 ;
        RECT 95.660 162.585 96.190 162.950 ;
        RECT 97.115 162.585 97.370 163.155 ;
        RECT 97.820 162.620 98.065 163.225 ;
        RECT 98.975 162.585 99.165 163.945 ;
        RECT 99.335 163.605 99.610 163.745 ;
        RECT 99.335 163.435 99.615 163.605 ;
        RECT 99.335 162.585 99.610 163.435 ;
        RECT 99.815 163.145 99.985 163.945 ;
        RECT 100.155 163.155 100.325 164.285 ;
        RECT 100.495 163.655 100.665 164.625 ;
        RECT 101.175 163.825 101.510 164.795 ;
        RECT 100.495 163.325 100.690 163.655 ;
        RECT 100.915 163.325 101.170 163.655 ;
        RECT 100.915 163.155 101.085 163.325 ;
        RECT 101.340 163.155 101.510 163.825 ;
        RECT 100.155 162.985 101.085 163.155 ;
        RECT 100.155 162.950 100.330 162.985 ;
        RECT 99.800 162.585 100.330 162.950 ;
        RECT 101.255 162.585 101.510 163.155 ;
        RECT 102.145 163.825 102.530 164.795 ;
        RECT 103.545 164.335 103.825 164.795 ;
        RECT 102.700 164.115 103.825 164.335 ;
        RECT 102.145 163.155 102.425 163.825 ;
        RECT 102.700 163.655 103.150 164.115 ;
        RECT 104.015 163.945 104.415 164.795 ;
        RECT 105.255 164.335 105.540 164.795 ;
        RECT 102.595 163.325 103.150 163.655 ;
        RECT 103.320 163.385 104.415 163.945 ;
        RECT 102.700 163.215 103.150 163.325 ;
        RECT 102.145 162.585 102.530 163.155 ;
        RECT 102.700 163.045 103.825 163.215 ;
        RECT 103.545 162.585 103.825 163.045 ;
        RECT 104.015 162.585 104.415 163.385 ;
        RECT 104.585 164.115 105.540 164.335 ;
        RECT 104.585 163.215 104.795 164.115 ;
        RECT 104.965 163.385 105.655 163.945 ;
        RECT 106.750 163.825 107.085 164.795 ;
        RECT 107.595 164.625 109.625 164.795 ;
        RECT 104.585 163.045 105.540 163.215 ;
        RECT 105.255 162.585 105.540 163.045 ;
        RECT 106.750 163.155 106.920 163.825 ;
        RECT 107.595 163.655 107.765 164.625 ;
        RECT 107.090 163.325 107.345 163.655 ;
        RECT 107.570 163.325 107.765 163.655 ;
        RECT 107.935 164.285 109.060 164.455 ;
        RECT 107.175 163.155 107.345 163.325 ;
        RECT 107.935 163.155 108.105 164.285 ;
        RECT 106.750 162.585 107.005 163.155 ;
        RECT 107.175 162.985 108.105 163.155 ;
        RECT 108.275 163.945 109.285 164.115 ;
        RECT 108.275 163.145 108.445 163.945 ;
        RECT 107.930 162.950 108.105 162.985 ;
        RECT 107.930 162.585 108.460 162.950 ;
        RECT 108.650 162.925 108.925 163.745 ;
        RECT 108.645 162.755 108.925 162.925 ;
        RECT 108.650 162.585 108.925 162.755 ;
        RECT 109.095 162.585 109.285 163.945 ;
        RECT 109.455 163.960 109.625 164.625 ;
        RECT 110.200 164.205 110.715 164.615 ;
        RECT 109.455 163.770 110.205 163.960 ;
        RECT 110.375 163.395 110.715 164.205 ;
        RECT 109.485 163.225 110.715 163.395 ;
        RECT 111.325 163.815 111.655 164.795 ;
        RECT 110.195 162.620 110.440 163.225 ;
        RECT 111.325 163.215 111.575 163.815 ;
        RECT 113.190 163.775 113.445 164.655 ;
        RECT 114.770 164.415 114.940 164.705 ;
        RECT 114.140 164.245 114.940 164.415 ;
        RECT 115.530 164.455 116.400 164.795 ;
        RECT 111.745 163.405 112.075 163.655 ;
        RECT 111.325 162.585 111.655 163.215 ;
        RECT 113.190 163.125 113.400 163.775 ;
        RECT 114.140 163.655 114.310 164.245 ;
        RECT 115.530 164.075 115.700 164.455 ;
        RECT 116.635 164.335 116.805 164.795 ;
        RECT 117.640 164.365 117.810 164.705 ;
        RECT 118.545 164.365 118.715 164.705 ;
        RECT 114.480 163.905 115.700 164.075 ;
        RECT 115.870 163.995 116.330 164.285 ;
        RECT 116.635 164.165 117.195 164.335 ;
        RECT 117.640 164.195 118.715 164.365 ;
        RECT 118.885 164.465 119.565 164.795 ;
        RECT 119.780 164.465 120.030 164.795 ;
        RECT 117.025 164.025 117.195 164.165 ;
        RECT 115.870 163.985 116.835 163.995 ;
        RECT 115.530 163.815 115.700 163.905 ;
        RECT 116.160 163.825 116.835 163.985 ;
        RECT 113.570 163.625 114.310 163.655 ;
        RECT 113.570 163.325 114.485 163.625 ;
        RECT 114.160 163.150 114.485 163.325 ;
        RECT 113.190 162.595 113.445 163.125 ;
        RECT 114.165 162.795 114.485 163.150 ;
        RECT 114.655 163.365 115.195 163.735 ;
        RECT 115.530 163.645 115.935 163.815 ;
        RECT 114.655 162.965 114.895 163.365 ;
        RECT 115.375 163.195 115.595 163.475 ;
        RECT 115.065 163.025 115.595 163.195 ;
        RECT 115.065 162.795 115.235 163.025 ;
        RECT 114.165 162.625 115.235 162.795 ;
        RECT 115.765 162.865 115.935 163.645 ;
        RECT 116.105 163.035 116.455 163.655 ;
        RECT 116.625 163.035 116.835 163.825 ;
        RECT 117.025 163.855 118.525 164.025 ;
        RECT 117.025 163.165 117.195 163.855 ;
        RECT 118.885 163.685 119.055 164.465 ;
        RECT 119.860 164.335 120.030 164.465 ;
        RECT 117.365 163.515 119.055 163.685 ;
        RECT 119.225 163.905 119.690 164.295 ;
        RECT 119.860 164.165 120.255 164.335 ;
        RECT 117.365 163.335 117.535 163.515 ;
        RECT 115.765 162.585 116.715 162.865 ;
        RECT 117.025 162.775 117.285 163.165 ;
        RECT 117.705 163.095 118.495 163.345 ;
        RECT 116.935 162.605 117.285 162.775 ;
        RECT 118.700 162.805 118.870 163.515 ;
        RECT 119.225 163.315 119.395 163.905 ;
        RECT 119.040 163.095 119.395 163.315 ;
        RECT 119.565 163.095 119.915 163.715 ;
        RECT 120.085 162.805 120.255 164.165 ;
        RECT 120.620 163.995 120.945 164.780 ;
        RECT 120.425 162.945 120.885 163.995 ;
        RECT 118.700 162.635 119.555 162.805 ;
        RECT 119.760 162.635 120.255 162.805 ;
        RECT 121.115 162.675 121.285 164.795 ;
        RECT 121.955 164.295 122.210 164.795 ;
        RECT 121.460 164.125 122.210 164.295 ;
        RECT 121.460 163.135 121.690 164.125 ;
        RECT 121.860 163.305 122.210 163.955 ;
        RECT 122.385 163.890 122.655 164.795 ;
        RECT 123.335 164.035 123.505 164.795 ;
        RECT 121.460 162.965 122.210 163.135 ;
        RECT 121.955 162.675 122.210 162.965 ;
        RECT 122.385 163.090 122.555 163.890 ;
        RECT 122.840 163.865 123.505 164.035 ;
        RECT 122.840 163.720 123.010 163.865 ;
        RECT 122.725 163.390 123.010 163.720 ;
        RECT 122.840 163.135 123.010 163.390 ;
        RECT 123.245 163.315 123.575 163.685 ;
        RECT 122.385 162.585 122.645 163.090 ;
        RECT 122.840 162.965 123.505 163.135 ;
        RECT 123.335 162.585 123.505 162.965 ;
        RECT 18.340 161.535 18.595 162.065 ;
        RECT 18.340 160.675 18.520 161.535 ;
        RECT 19.240 161.335 19.490 161.985 ;
        RECT 18.690 161.005 19.490 161.335 ;
        RECT 18.340 160.205 18.595 160.675 ;
        RECT 18.255 160.035 18.595 160.205 ;
        RECT 18.340 160.005 18.595 160.035 ;
        RECT 19.240 160.415 19.490 161.005 ;
        RECT 19.690 161.650 20.010 161.980 ;
        RECT 21.050 161.855 21.900 162.025 ;
        RECT 19.690 160.755 19.880 161.650 ;
        RECT 20.200 161.325 20.860 161.595 ;
        RECT 20.530 161.265 20.860 161.325 ;
        RECT 20.050 161.095 20.380 161.155 ;
        RECT 21.050 161.095 21.220 161.855 ;
        RECT 22.980 161.605 23.230 162.035 ;
        RECT 21.390 161.435 22.640 161.605 ;
        RECT 21.390 161.315 21.720 161.435 ;
        RECT 20.050 160.925 21.950 161.095 ;
        RECT 19.690 160.585 21.610 160.755 ;
        RECT 19.690 160.565 20.010 160.585 ;
        RECT 19.240 159.905 19.570 160.415 ;
        RECT 19.840 159.955 20.010 160.565 ;
        RECT 21.780 160.415 21.950 160.925 ;
        RECT 22.120 160.855 22.300 161.265 ;
        RECT 22.470 160.675 22.640 161.435 ;
        RECT 20.740 160.245 21.950 160.415 ;
        RECT 22.120 160.365 22.640 160.675 ;
        RECT 22.810 161.265 23.230 161.605 ;
        RECT 24.100 161.865 25.115 162.065 ;
        RECT 23.520 161.265 23.930 161.595 ;
        RECT 22.810 160.495 23.000 161.265 ;
        RECT 24.100 161.135 24.270 161.865 ;
        RECT 25.415 161.695 25.585 162.025 ;
        RECT 24.440 161.315 24.790 161.685 ;
        RECT 24.100 161.095 24.520 161.135 ;
        RECT 23.170 160.925 24.520 161.095 ;
        RECT 23.170 160.765 23.420 160.925 ;
        RECT 23.930 160.495 24.180 160.755 ;
        RECT 22.810 160.245 24.180 160.495 ;
        RECT 20.740 159.955 20.980 160.245 ;
        RECT 21.780 160.165 21.950 160.245 ;
        RECT 21.780 159.915 22.410 160.165 ;
        RECT 23.380 159.955 23.550 160.245 ;
        RECT 24.350 160.080 24.520 160.925 ;
        RECT 24.970 160.755 25.190 161.625 ;
        RECT 25.415 161.505 26.110 161.695 ;
        RECT 24.690 160.375 25.190 160.755 ;
        RECT 25.360 160.705 25.770 161.325 ;
        RECT 25.940 160.535 26.110 161.505 ;
        RECT 25.415 160.365 26.110 160.535 ;
        RECT 24.350 159.910 25.180 160.080 ;
        RECT 25.415 159.865 25.585 160.365 ;
        RECT 26.300 159.865 26.525 161.985 ;
        RECT 27.195 161.695 27.365 161.985 ;
        RECT 26.700 161.525 27.365 161.695 ;
        RECT 26.700 160.535 26.930 161.525 ;
        RECT 27.630 161.505 27.885 162.075 ;
        RECT 28.810 161.710 29.340 162.075 ;
        RECT 28.810 161.675 28.985 161.710 ;
        RECT 28.055 161.505 28.985 161.675 ;
        RECT 27.100 160.705 27.450 161.355 ;
        RECT 27.630 160.835 27.800 161.505 ;
        RECT 28.055 161.335 28.225 161.505 ;
        RECT 27.970 161.005 28.225 161.335 ;
        RECT 28.450 161.005 28.645 161.335 ;
        RECT 26.700 160.365 27.365 160.535 ;
        RECT 27.195 159.865 27.365 160.365 ;
        RECT 27.630 159.865 27.965 160.835 ;
        RECT 28.475 160.035 28.645 161.005 ;
        RECT 28.815 160.375 28.985 161.505 ;
        RECT 29.155 160.715 29.325 161.515 ;
        RECT 29.530 161.225 29.805 162.075 ;
        RECT 29.525 161.055 29.805 161.225 ;
        RECT 29.530 160.915 29.805 161.055 ;
        RECT 29.975 160.715 30.165 162.075 ;
        RECT 31.075 161.435 31.320 162.040 ;
        RECT 33.420 161.435 33.665 162.040 ;
        RECT 30.365 161.265 31.595 161.435 ;
        RECT 29.155 160.545 30.165 160.715 ;
        RECT 30.335 160.700 31.085 160.890 ;
        RECT 28.815 160.205 29.940 160.375 ;
        RECT 30.335 160.035 30.505 160.700 ;
        RECT 31.255 160.455 31.595 161.265 ;
        RECT 31.080 160.045 31.595 160.455 ;
        RECT 33.145 161.265 34.375 161.435 ;
        RECT 33.145 160.455 33.485 161.265 ;
        RECT 33.655 160.700 34.405 160.890 ;
        RECT 33.145 160.045 33.660 160.455 ;
        RECT 28.475 159.865 30.505 160.035 ;
        RECT 34.235 160.035 34.405 160.700 ;
        RECT 34.575 160.715 34.765 162.075 ;
        RECT 34.935 161.225 35.210 162.075 ;
        RECT 35.400 161.710 35.930 162.075 ;
        RECT 35.755 161.675 35.930 161.710 ;
        RECT 34.935 161.055 35.215 161.225 ;
        RECT 34.935 160.915 35.210 161.055 ;
        RECT 35.415 160.715 35.585 161.515 ;
        RECT 34.575 160.545 35.585 160.715 ;
        RECT 35.755 161.505 36.685 161.675 ;
        RECT 36.855 161.505 37.110 162.075 ;
        RECT 35.755 160.375 35.925 161.505 ;
        RECT 36.515 161.335 36.685 161.505 ;
        RECT 34.800 160.205 35.925 160.375 ;
        RECT 36.095 161.005 36.290 161.335 ;
        RECT 36.515 161.005 36.770 161.335 ;
        RECT 36.095 160.035 36.265 161.005 ;
        RECT 36.940 160.835 37.110 161.505 ;
        RECT 34.235 159.865 36.265 160.035 ;
        RECT 36.775 159.865 37.110 160.835 ;
        RECT 41.885 161.505 42.270 162.075 ;
        RECT 43.285 161.615 43.565 162.075 ;
        RECT 41.885 160.835 42.165 161.505 ;
        RECT 42.440 161.445 43.565 161.615 ;
        RECT 42.440 161.335 42.890 161.445 ;
        RECT 42.335 161.005 42.890 161.335 ;
        RECT 43.755 161.275 44.155 162.075 ;
        RECT 44.995 161.615 45.280 162.075 ;
        RECT 41.885 159.865 42.270 160.835 ;
        RECT 42.440 160.545 42.890 161.005 ;
        RECT 43.060 160.715 44.155 161.275 ;
        RECT 42.440 160.325 43.565 160.545 ;
        RECT 43.285 159.865 43.565 160.325 ;
        RECT 43.755 159.865 44.155 160.715 ;
        RECT 44.325 161.445 45.280 161.615 ;
        RECT 47.060 161.615 47.345 162.075 ;
        RECT 47.060 161.445 48.015 161.615 ;
        RECT 44.325 160.545 44.535 161.445 ;
        RECT 44.705 160.715 45.395 161.275 ;
        RECT 46.945 160.715 47.635 161.275 ;
        RECT 47.805 160.545 48.015 161.445 ;
        RECT 44.325 160.325 45.280 160.545 ;
        RECT 44.995 159.865 45.280 160.325 ;
        RECT 47.060 160.325 48.015 160.545 ;
        RECT 48.185 161.275 48.585 162.075 ;
        RECT 48.775 161.615 49.055 162.075 ;
        RECT 48.775 161.445 49.900 161.615 ;
        RECT 50.070 161.505 50.455 162.075 ;
        RECT 49.450 161.335 49.900 161.445 ;
        RECT 48.185 160.715 49.280 161.275 ;
        RECT 49.450 161.005 50.005 161.335 ;
        RECT 47.060 159.865 47.345 160.325 ;
        RECT 48.185 159.865 48.585 160.715 ;
        RECT 49.450 160.545 49.900 161.005 ;
        RECT 50.175 160.835 50.455 161.505 ;
        RECT 50.900 161.435 51.145 162.040 ;
        RECT 48.775 160.325 49.900 160.545 ;
        RECT 48.775 159.865 49.055 160.325 ;
        RECT 50.070 159.865 50.455 160.835 ;
        RECT 50.625 161.265 51.855 161.435 ;
        RECT 50.625 160.455 50.965 161.265 ;
        RECT 51.135 160.700 51.885 160.890 ;
        RECT 50.625 160.045 51.140 160.455 ;
        RECT 51.715 160.035 51.885 160.700 ;
        RECT 52.055 160.715 52.245 162.075 ;
        RECT 52.415 161.565 52.690 162.075 ;
        RECT 52.880 161.710 53.410 162.075 ;
        RECT 53.235 161.675 53.410 161.710 ;
        RECT 52.415 161.395 52.695 161.565 ;
        RECT 52.415 160.915 52.690 161.395 ;
        RECT 52.895 160.715 53.065 161.515 ;
        RECT 52.055 160.545 53.065 160.715 ;
        RECT 53.235 161.505 54.165 161.675 ;
        RECT 54.335 161.505 54.590 162.075 ;
        RECT 53.235 160.375 53.405 161.505 ;
        RECT 53.995 161.335 54.165 161.505 ;
        RECT 52.280 160.205 53.405 160.375 ;
        RECT 53.575 161.005 53.770 161.335 ;
        RECT 53.995 161.005 54.250 161.335 ;
        RECT 53.575 160.035 53.745 161.005 ;
        RECT 54.420 160.835 54.590 161.505 ;
        RECT 54.880 161.615 55.165 162.075 ;
        RECT 54.880 161.445 55.835 161.615 ;
        RECT 51.715 159.865 53.745 160.035 ;
        RECT 54.255 159.865 54.590 160.835 ;
        RECT 54.765 160.715 55.455 161.275 ;
        RECT 55.625 160.545 55.835 161.445 ;
        RECT 54.880 160.325 55.835 160.545 ;
        RECT 56.005 161.275 56.405 162.075 ;
        RECT 56.595 161.615 56.875 162.075 ;
        RECT 56.595 161.445 57.720 161.615 ;
        RECT 57.890 161.505 58.275 162.075 ;
        RECT 58.995 161.695 59.165 162.075 ;
        RECT 58.995 161.525 59.660 161.695 ;
        RECT 59.855 161.570 60.115 162.075 ;
        RECT 57.270 161.335 57.720 161.445 ;
        RECT 56.005 160.715 57.100 161.275 ;
        RECT 57.270 161.005 57.825 161.335 ;
        RECT 54.880 159.865 55.165 160.325 ;
        RECT 56.005 159.865 56.405 160.715 ;
        RECT 57.270 160.545 57.720 161.005 ;
        RECT 57.995 160.835 58.275 161.505 ;
        RECT 58.925 160.975 59.255 161.345 ;
        RECT 59.490 161.270 59.660 161.525 ;
        RECT 56.595 160.325 57.720 160.545 ;
        RECT 56.595 159.865 56.875 160.325 ;
        RECT 57.890 159.865 58.275 160.835 ;
        RECT 59.490 160.940 59.775 161.270 ;
        RECT 59.490 160.795 59.660 160.940 ;
        RECT 58.995 160.625 59.660 160.795 ;
        RECT 59.945 160.770 60.115 161.570 ;
        RECT 58.995 159.865 59.165 160.625 ;
        RECT 59.845 159.865 60.115 160.770 ;
        RECT 65.325 161.500 65.580 162.075 ;
        RECT 66.295 161.695 66.465 162.075 ;
        RECT 65.750 161.525 66.465 161.695 ;
        RECT 65.325 160.770 65.495 161.500 ;
        RECT 65.750 161.335 65.920 161.525 ;
        RECT 67.165 161.500 67.420 162.075 ;
        RECT 68.135 161.695 68.305 162.075 ;
        RECT 67.590 161.525 68.305 161.695 ;
        RECT 68.655 161.695 68.825 162.075 ;
        RECT 68.655 161.525 69.370 161.695 ;
        RECT 65.665 161.005 65.920 161.335 ;
        RECT 65.750 160.795 65.920 161.005 ;
        RECT 66.200 160.975 66.555 161.345 ;
        RECT 65.325 159.865 65.580 160.770 ;
        RECT 65.750 160.625 66.465 160.795 ;
        RECT 66.295 159.865 66.465 160.625 ;
        RECT 67.165 160.770 67.335 161.500 ;
        RECT 67.590 161.335 67.760 161.525 ;
        RECT 67.505 161.005 67.760 161.335 ;
        RECT 67.590 160.795 67.760 161.005 ;
        RECT 68.040 160.975 68.395 161.345 ;
        RECT 68.565 160.975 68.920 161.345 ;
        RECT 69.200 161.335 69.370 161.525 ;
        RECT 69.540 161.500 69.795 162.075 ;
        RECT 70.495 161.695 70.665 162.075 ;
        RECT 70.495 161.525 71.210 161.695 ;
        RECT 69.200 161.005 69.455 161.335 ;
        RECT 69.200 160.795 69.370 161.005 ;
        RECT 67.165 159.865 67.420 160.770 ;
        RECT 67.590 160.625 68.305 160.795 ;
        RECT 68.135 159.865 68.305 160.625 ;
        RECT 68.655 160.625 69.370 160.795 ;
        RECT 69.625 160.770 69.795 161.500 ;
        RECT 70.405 160.975 70.760 161.345 ;
        RECT 71.040 161.335 71.210 161.525 ;
        RECT 71.380 161.500 71.635 162.075 ;
        RECT 71.040 161.005 71.295 161.335 ;
        RECT 71.040 160.795 71.210 161.005 ;
        RECT 68.655 159.865 68.825 160.625 ;
        RECT 69.540 159.865 69.795 160.770 ;
        RECT 70.495 160.625 71.210 160.795 ;
        RECT 71.465 160.770 71.635 161.500 ;
        RECT 70.495 159.865 70.665 160.625 ;
        RECT 71.380 159.865 71.635 160.770 ;
        RECT 80.965 161.445 81.295 162.075 ;
        RECT 80.965 160.845 81.215 161.445 ;
        RECT 82.180 161.435 82.425 162.040 ;
        RECT 81.905 161.265 83.135 161.435 ;
        RECT 81.385 161.005 81.715 161.255 ;
        RECT 80.965 159.865 81.295 160.845 ;
        RECT 81.905 160.455 82.245 161.265 ;
        RECT 82.415 160.700 83.165 160.890 ;
        RECT 81.905 160.045 82.420 160.455 ;
        RECT 82.995 160.035 83.165 160.700 ;
        RECT 83.335 160.715 83.525 162.075 ;
        RECT 83.695 161.225 83.970 162.075 ;
        RECT 84.160 161.710 84.690 162.075 ;
        RECT 84.515 161.675 84.690 161.710 ;
        RECT 83.695 161.055 83.975 161.225 ;
        RECT 83.695 160.915 83.970 161.055 ;
        RECT 84.175 160.715 84.345 161.515 ;
        RECT 83.335 160.545 84.345 160.715 ;
        RECT 84.515 161.505 85.445 161.675 ;
        RECT 85.615 161.505 85.870 162.075 ;
        RECT 86.595 161.695 86.765 162.075 ;
        RECT 86.595 161.525 87.260 161.695 ;
        RECT 87.455 161.570 87.715 162.075 ;
        RECT 89.640 161.905 89.895 162.065 ;
        RECT 89.555 161.735 89.895 161.905 ;
        RECT 84.515 160.375 84.685 161.505 ;
        RECT 85.275 161.335 85.445 161.505 ;
        RECT 83.560 160.205 84.685 160.375 ;
        RECT 84.855 161.005 85.050 161.335 ;
        RECT 85.275 161.005 85.530 161.335 ;
        RECT 84.855 160.035 85.025 161.005 ;
        RECT 85.700 160.835 85.870 161.505 ;
        RECT 86.525 160.975 86.855 161.345 ;
        RECT 87.090 161.270 87.260 161.525 ;
        RECT 82.995 159.865 85.025 160.035 ;
        RECT 85.535 159.865 85.870 160.835 ;
        RECT 87.090 160.940 87.375 161.270 ;
        RECT 87.090 160.795 87.260 160.940 ;
        RECT 86.595 160.625 87.260 160.795 ;
        RECT 87.545 160.770 87.715 161.570 ;
        RECT 86.595 159.865 86.765 160.625 ;
        RECT 87.445 159.865 87.715 160.770 ;
        RECT 89.640 161.535 89.895 161.735 ;
        RECT 89.640 160.675 89.820 161.535 ;
        RECT 90.540 161.335 90.790 161.985 ;
        RECT 89.990 161.005 90.790 161.335 ;
        RECT 89.640 160.005 89.895 160.675 ;
        RECT 90.540 160.415 90.790 161.005 ;
        RECT 90.990 161.650 91.310 161.980 ;
        RECT 92.350 161.855 93.200 162.025 ;
        RECT 90.990 160.755 91.180 161.650 ;
        RECT 91.500 161.325 92.160 161.595 ;
        RECT 91.830 161.265 92.160 161.325 ;
        RECT 91.350 161.095 91.680 161.155 ;
        RECT 92.350 161.095 92.520 161.855 ;
        RECT 94.280 161.605 94.530 162.035 ;
        RECT 92.690 161.435 93.940 161.605 ;
        RECT 92.690 161.315 93.020 161.435 ;
        RECT 91.350 160.925 93.250 161.095 ;
        RECT 90.990 160.585 92.910 160.755 ;
        RECT 90.990 160.565 91.310 160.585 ;
        RECT 90.540 159.905 90.870 160.415 ;
        RECT 91.140 159.955 91.310 160.565 ;
        RECT 93.080 160.415 93.250 160.925 ;
        RECT 93.420 160.855 93.600 161.265 ;
        RECT 93.770 160.675 93.940 161.435 ;
        RECT 92.040 160.245 93.250 160.415 ;
        RECT 93.420 160.365 93.940 160.675 ;
        RECT 94.110 161.265 94.530 161.605 ;
        RECT 95.400 161.865 96.415 162.065 ;
        RECT 94.820 161.265 95.230 161.595 ;
        RECT 94.110 160.495 94.300 161.265 ;
        RECT 95.400 161.135 95.570 161.865 ;
        RECT 96.715 161.695 96.885 162.025 ;
        RECT 95.740 161.315 96.090 161.685 ;
        RECT 95.400 161.095 95.820 161.135 ;
        RECT 94.470 160.925 95.820 161.095 ;
        RECT 94.470 160.765 94.720 160.925 ;
        RECT 95.230 160.495 95.480 160.755 ;
        RECT 94.110 160.245 95.480 160.495 ;
        RECT 92.040 159.955 92.280 160.245 ;
        RECT 93.080 160.165 93.250 160.245 ;
        RECT 93.080 159.915 93.710 160.165 ;
        RECT 94.680 159.955 94.850 160.245 ;
        RECT 95.650 160.080 95.820 160.925 ;
        RECT 96.270 160.755 96.490 161.625 ;
        RECT 96.715 161.505 97.410 161.695 ;
        RECT 95.990 160.375 96.490 160.755 ;
        RECT 96.660 160.705 97.070 161.325 ;
        RECT 97.240 160.535 97.410 161.505 ;
        RECT 96.715 160.365 97.410 160.535 ;
        RECT 95.650 159.910 96.480 160.080 ;
        RECT 96.715 159.865 96.885 160.365 ;
        RECT 97.600 159.865 97.825 161.985 ;
        RECT 98.495 161.695 98.665 161.985 ;
        RECT 98.000 161.525 98.665 161.695 ;
        RECT 99.935 161.695 100.105 162.075 ;
        RECT 99.935 161.525 100.600 161.695 ;
        RECT 100.795 161.570 101.055 162.075 ;
        RECT 98.000 160.535 98.230 161.525 ;
        RECT 98.400 160.705 98.750 161.355 ;
        RECT 99.865 160.975 100.195 161.345 ;
        RECT 100.430 161.270 100.600 161.525 ;
        RECT 100.430 160.940 100.715 161.270 ;
        RECT 100.430 160.795 100.600 160.940 ;
        RECT 99.935 160.625 100.600 160.795 ;
        RECT 100.885 160.770 101.055 161.570 ;
        RECT 98.000 160.365 98.665 160.535 ;
        RECT 98.495 159.865 98.665 160.365 ;
        RECT 99.935 159.865 100.105 160.625 ;
        RECT 100.785 159.865 101.055 160.770 ;
        RECT 101.665 161.445 101.995 162.075 ;
        RECT 102.605 161.505 102.990 162.075 ;
        RECT 104.005 161.615 104.285 162.075 ;
        RECT 101.665 160.845 101.915 161.445 ;
        RECT 102.085 161.005 102.415 161.255 ;
        RECT 101.665 159.865 101.995 160.845 ;
        RECT 102.605 160.835 102.885 161.505 ;
        RECT 103.160 161.445 104.285 161.615 ;
        RECT 103.160 161.335 103.610 161.445 ;
        RECT 103.055 161.005 103.610 161.335 ;
        RECT 104.475 161.275 104.875 162.075 ;
        RECT 105.715 161.615 106.000 162.075 ;
        RECT 102.605 159.865 102.990 160.835 ;
        RECT 103.160 160.545 103.610 161.005 ;
        RECT 103.780 160.715 104.875 161.275 ;
        RECT 103.160 160.325 104.285 160.545 ;
        RECT 104.005 159.865 104.285 160.325 ;
        RECT 104.475 159.865 104.875 160.715 ;
        RECT 105.045 161.445 106.000 161.615 ;
        RECT 106.860 161.615 107.145 162.075 ;
        RECT 106.860 161.445 107.815 161.615 ;
        RECT 105.045 160.545 105.255 161.445 ;
        RECT 105.425 160.715 106.115 161.275 ;
        RECT 106.745 160.715 107.435 161.275 ;
        RECT 107.605 160.545 107.815 161.445 ;
        RECT 105.045 160.325 106.000 160.545 ;
        RECT 105.715 159.865 106.000 160.325 ;
        RECT 106.860 160.325 107.815 160.545 ;
        RECT 107.985 161.275 108.385 162.075 ;
        RECT 108.575 161.615 108.855 162.075 ;
        RECT 108.575 161.445 109.700 161.615 ;
        RECT 109.870 161.505 110.255 162.075 ;
        RECT 109.250 161.335 109.700 161.445 ;
        RECT 107.985 160.715 109.080 161.275 ;
        RECT 109.250 161.005 109.805 161.335 ;
        RECT 106.860 159.865 107.145 160.325 ;
        RECT 107.985 159.865 108.385 160.715 ;
        RECT 109.250 160.545 109.700 161.005 ;
        RECT 109.975 160.835 110.255 161.505 ;
        RECT 110.700 161.435 110.945 162.040 ;
        RECT 108.575 160.325 109.700 160.545 ;
        RECT 108.575 159.865 108.855 160.325 ;
        RECT 109.870 159.865 110.255 160.835 ;
        RECT 110.425 161.265 111.655 161.435 ;
        RECT 110.425 160.455 110.765 161.265 ;
        RECT 110.935 160.700 111.685 160.890 ;
        RECT 110.425 160.045 110.940 160.455 ;
        RECT 111.515 160.035 111.685 160.700 ;
        RECT 111.855 160.715 112.045 162.075 ;
        RECT 112.215 161.225 112.490 162.075 ;
        RECT 112.680 161.710 113.210 162.075 ;
        RECT 113.035 161.675 113.210 161.710 ;
        RECT 112.215 161.055 112.495 161.225 ;
        RECT 112.215 160.915 112.490 161.055 ;
        RECT 112.695 160.715 112.865 161.515 ;
        RECT 111.855 160.545 112.865 160.715 ;
        RECT 113.035 161.505 113.965 161.675 ;
        RECT 114.135 161.505 114.390 162.075 ;
        RECT 113.035 160.375 113.205 161.505 ;
        RECT 113.795 161.335 113.965 161.505 ;
        RECT 112.080 160.205 113.205 160.375 ;
        RECT 113.375 161.005 113.570 161.335 ;
        RECT 113.795 161.005 114.050 161.335 ;
        RECT 113.375 160.035 113.545 161.005 ;
        RECT 114.220 160.835 114.390 161.505 ;
        RECT 115.300 161.435 115.545 162.040 ;
        RECT 111.515 159.865 113.545 160.035 ;
        RECT 114.055 159.865 114.390 160.835 ;
        RECT 115.025 161.265 116.255 161.435 ;
        RECT 115.025 160.455 115.365 161.265 ;
        RECT 115.535 160.700 116.285 160.890 ;
        RECT 115.025 160.045 115.540 160.455 ;
        RECT 116.115 160.035 116.285 160.700 ;
        RECT 116.455 160.715 116.645 162.075 ;
        RECT 116.815 161.905 117.090 162.075 ;
        RECT 116.815 161.735 117.095 161.905 ;
        RECT 116.815 160.915 117.090 161.735 ;
        RECT 117.280 161.710 117.810 162.075 ;
        RECT 117.635 161.675 117.810 161.710 ;
        RECT 117.295 160.715 117.465 161.515 ;
        RECT 116.455 160.545 117.465 160.715 ;
        RECT 117.635 161.505 118.565 161.675 ;
        RECT 118.735 161.505 118.990 162.075 ;
        RECT 117.635 160.375 117.805 161.505 ;
        RECT 118.395 161.335 118.565 161.505 ;
        RECT 116.680 160.205 117.805 160.375 ;
        RECT 117.975 161.005 118.170 161.335 ;
        RECT 118.395 161.005 118.650 161.335 ;
        RECT 117.975 160.035 118.145 161.005 ;
        RECT 118.820 160.835 118.990 161.505 ;
        RECT 119.280 161.615 119.565 162.075 ;
        RECT 119.280 161.445 120.235 161.615 ;
        RECT 116.115 159.865 118.145 160.035 ;
        RECT 118.655 159.865 118.990 160.835 ;
        RECT 119.165 160.715 119.855 161.275 ;
        RECT 120.025 160.545 120.235 161.445 ;
        RECT 119.280 160.325 120.235 160.545 ;
        RECT 120.405 161.275 120.805 162.075 ;
        RECT 120.995 161.615 121.275 162.075 ;
        RECT 120.995 161.445 122.120 161.615 ;
        RECT 122.290 161.505 122.675 162.075 ;
        RECT 122.935 161.695 123.105 162.075 ;
        RECT 122.935 161.525 123.600 161.695 ;
        RECT 123.795 161.570 124.055 162.075 ;
        RECT 121.670 161.335 122.120 161.445 ;
        RECT 120.405 160.715 121.500 161.275 ;
        RECT 121.670 161.005 122.225 161.335 ;
        RECT 119.280 159.865 119.565 160.325 ;
        RECT 120.405 159.865 120.805 160.715 ;
        RECT 121.670 160.545 122.120 161.005 ;
        RECT 122.395 160.835 122.675 161.505 ;
        RECT 122.865 160.975 123.195 161.345 ;
        RECT 123.430 161.270 123.600 161.525 ;
        RECT 120.995 160.325 122.120 160.545 ;
        RECT 120.995 159.865 121.275 160.325 ;
        RECT 122.290 159.865 122.675 160.835 ;
        RECT 123.430 160.940 123.715 161.270 ;
        RECT 123.430 160.795 123.600 160.940 ;
        RECT 122.935 160.625 123.600 160.795 ;
        RECT 123.885 160.770 124.055 161.570 ;
        RECT 122.935 159.865 123.105 160.625 ;
        RECT 123.785 159.865 124.055 160.770 ;
        RECT 17.945 158.375 18.275 159.355 ;
        RECT 19.325 158.375 19.655 159.355 ;
        RECT 21.355 159.185 23.385 159.355 ;
        RECT 17.945 157.775 18.195 158.375 ;
        RECT 18.365 157.965 18.695 158.215 ;
        RECT 18.905 157.965 19.235 158.215 ;
        RECT 19.405 157.775 19.655 158.375 ;
        RECT 20.265 158.765 20.780 159.175 ;
        RECT 20.265 157.955 20.605 158.765 ;
        RECT 21.355 158.520 21.525 159.185 ;
        RECT 21.920 158.845 23.045 159.015 ;
        RECT 20.775 158.330 21.525 158.520 ;
        RECT 21.695 158.505 22.705 158.675 ;
        RECT 20.265 157.785 21.495 157.955 ;
        RECT 17.945 157.145 18.275 157.775 ;
        RECT 19.325 157.145 19.655 157.775 ;
        RECT 20.540 157.180 20.785 157.785 ;
        RECT 21.695 157.145 21.885 158.505 ;
        RECT 22.055 157.485 22.330 158.305 ;
        RECT 22.535 157.705 22.705 158.505 ;
        RECT 22.875 157.715 23.045 158.845 ;
        RECT 23.215 158.215 23.385 159.185 ;
        RECT 23.895 158.385 24.230 159.355 ;
        RECT 24.955 158.595 25.125 159.355 ;
        RECT 24.955 158.425 25.620 158.595 ;
        RECT 25.805 158.450 26.075 159.355 ;
        RECT 23.215 157.885 23.410 158.215 ;
        RECT 23.635 157.885 23.890 158.215 ;
        RECT 23.635 157.715 23.805 157.885 ;
        RECT 24.060 157.715 24.230 158.385 ;
        RECT 25.450 158.280 25.620 158.425 ;
        RECT 24.885 157.875 25.215 158.245 ;
        RECT 25.450 157.950 25.735 158.280 ;
        RECT 22.875 157.545 23.805 157.715 ;
        RECT 22.875 157.510 23.050 157.545 ;
        RECT 22.055 157.315 22.335 157.485 ;
        RECT 22.055 157.145 22.330 157.315 ;
        RECT 22.520 157.145 23.050 157.510 ;
        RECT 23.975 157.145 24.230 157.715 ;
        RECT 25.450 157.695 25.620 157.950 ;
        RECT 24.955 157.525 25.620 157.695 ;
        RECT 25.905 157.650 26.075 158.450 ;
        RECT 24.955 157.145 25.125 157.525 ;
        RECT 25.815 157.145 26.075 157.650 ;
        RECT 32.225 158.385 32.610 159.355 ;
        RECT 33.625 158.895 33.905 159.355 ;
        RECT 32.780 158.675 33.905 158.895 ;
        RECT 32.225 157.715 32.505 158.385 ;
        RECT 32.780 158.215 33.230 158.675 ;
        RECT 34.095 158.505 34.495 159.355 ;
        RECT 35.335 158.895 35.620 159.355 ;
        RECT 32.675 157.885 33.230 158.215 ;
        RECT 33.400 157.945 34.495 158.505 ;
        RECT 32.780 157.775 33.230 157.885 ;
        RECT 32.225 157.145 32.610 157.715 ;
        RECT 32.780 157.605 33.905 157.775 ;
        RECT 33.625 157.145 33.905 157.605 ;
        RECT 34.095 157.145 34.495 157.945 ;
        RECT 34.665 158.675 35.620 158.895 ;
        RECT 34.665 157.775 34.875 158.675 ;
        RECT 43.010 158.555 43.340 159.355 ;
        RECT 44.140 158.555 44.470 159.355 ;
        RECT 35.045 157.945 35.735 158.505 ;
        RECT 43.010 158.385 45.445 158.555 ;
        RECT 45.975 158.385 46.315 159.355 ;
        RECT 42.805 157.965 43.155 158.215 ;
        RECT 34.665 157.605 35.620 157.775 ;
        RECT 43.340 157.755 43.510 158.385 ;
        RECT 43.680 157.965 44.010 158.165 ;
        RECT 44.180 157.965 44.510 158.165 ;
        RECT 44.680 157.965 45.100 158.165 ;
        RECT 45.275 158.135 45.445 158.385 ;
        RECT 45.275 157.965 45.970 158.135 ;
        RECT 35.335 157.145 35.620 157.605 ;
        RECT 43.010 157.145 43.510 157.755 ;
        RECT 44.140 157.625 45.365 157.795 ;
        RECT 46.140 157.775 46.315 158.385 ;
        RECT 44.140 157.145 44.470 157.625 ;
        RECT 45.035 157.145 45.365 157.625 ;
        RECT 45.975 157.145 46.315 157.775 ;
        RECT 46.485 158.385 46.825 159.355 ;
        RECT 48.330 158.555 48.660 159.355 ;
        RECT 49.460 158.555 49.790 159.355 ;
        RECT 47.355 158.385 49.790 158.555 ;
        RECT 50.625 158.385 50.965 159.355 ;
        RECT 52.470 158.555 52.800 159.355 ;
        RECT 53.600 158.555 53.930 159.355 ;
        RECT 51.495 158.385 53.930 158.555 ;
        RECT 54.765 158.450 55.035 159.355 ;
        RECT 55.715 158.595 55.885 159.355 ;
        RECT 46.485 157.775 46.660 158.385 ;
        RECT 47.355 158.135 47.525 158.385 ;
        RECT 46.830 157.965 47.525 158.135 ;
        RECT 47.700 157.965 48.120 158.165 ;
        RECT 48.290 157.965 48.620 158.165 ;
        RECT 48.790 157.965 49.120 158.165 ;
        RECT 46.485 157.145 46.825 157.775 ;
        RECT 47.435 157.625 48.660 157.795 ;
        RECT 47.435 157.145 47.765 157.625 ;
        RECT 48.330 157.145 48.660 157.625 ;
        RECT 49.290 157.755 49.460 158.385 ;
        RECT 49.645 157.965 49.995 158.215 ;
        RECT 50.625 157.775 50.800 158.385 ;
        RECT 51.495 158.135 51.665 158.385 ;
        RECT 50.970 157.965 51.665 158.135 ;
        RECT 51.840 157.965 52.260 158.165 ;
        RECT 52.430 157.965 52.760 158.165 ;
        RECT 52.930 157.965 53.260 158.165 ;
        RECT 49.290 157.145 49.790 157.755 ;
        RECT 50.625 157.145 50.965 157.775 ;
        RECT 51.575 157.625 52.800 157.795 ;
        RECT 51.575 157.145 51.905 157.625 ;
        RECT 52.470 157.145 52.800 157.625 ;
        RECT 53.430 157.755 53.600 158.385 ;
        RECT 53.785 157.965 54.135 158.215 ;
        RECT 53.430 157.145 53.930 157.755 ;
        RECT 54.765 157.650 54.935 158.450 ;
        RECT 55.220 158.425 55.885 158.595 ;
        RECT 62.315 158.505 62.485 159.355 ;
        RECT 63.155 158.505 63.325 159.355 ;
        RECT 63.915 158.545 64.245 159.355 ;
        RECT 55.220 158.280 55.390 158.425 ;
        RECT 55.105 157.950 55.390 158.280 ;
        RECT 62.315 158.335 63.325 158.505 ;
        RECT 63.530 158.375 64.245 158.545 ;
        RECT 68.655 158.595 68.825 159.355 ;
        RECT 68.655 158.425 69.370 158.595 ;
        RECT 69.540 158.450 69.795 159.355 ;
        RECT 55.220 157.695 55.390 157.950 ;
        RECT 55.625 157.875 55.955 158.245 ;
        RECT 62.315 158.165 62.810 158.335 ;
        RECT 62.315 157.995 62.815 158.165 ;
        RECT 63.530 158.135 63.700 158.375 ;
        RECT 62.315 157.795 62.810 157.995 ;
        RECT 63.200 157.965 63.700 158.135 ;
        RECT 63.870 157.965 64.250 158.205 ;
        RECT 63.530 157.795 63.700 157.965 ;
        RECT 68.565 157.875 68.920 158.245 ;
        RECT 69.200 158.215 69.370 158.425 ;
        RECT 69.200 157.885 69.455 158.215 ;
        RECT 54.765 157.145 55.025 157.650 ;
        RECT 55.220 157.525 55.885 157.695 ;
        RECT 55.715 157.145 55.885 157.525 ;
        RECT 62.315 157.625 63.325 157.795 ;
        RECT 63.530 157.625 64.165 157.795 ;
        RECT 69.200 157.695 69.370 157.885 ;
        RECT 69.625 157.720 69.795 158.450 ;
        RECT 70.495 158.595 70.665 159.355 ;
        RECT 70.495 158.425 71.210 158.595 ;
        RECT 71.380 158.450 71.635 159.355 ;
        RECT 70.405 157.875 70.760 158.245 ;
        RECT 71.040 158.215 71.210 158.425 ;
        RECT 71.040 157.885 71.295 158.215 ;
        RECT 62.315 157.145 62.485 157.625 ;
        RECT 63.155 157.145 63.325 157.625 ;
        RECT 63.995 157.145 64.165 157.625 ;
        RECT 68.655 157.525 69.370 157.695 ;
        RECT 68.655 157.145 68.825 157.525 ;
        RECT 69.540 157.145 69.795 157.720 ;
        RECT 71.040 157.695 71.210 157.885 ;
        RECT 71.465 157.720 71.635 158.450 ;
        RECT 72.450 158.555 72.780 159.355 ;
        RECT 73.580 158.555 73.910 159.355 ;
        RECT 72.450 158.385 74.885 158.555 ;
        RECT 75.415 158.385 75.755 159.355 ;
        RECT 72.245 157.965 72.595 158.215 ;
        RECT 72.780 157.755 72.950 158.385 ;
        RECT 73.120 157.965 73.450 158.165 ;
        RECT 73.620 157.965 73.950 158.165 ;
        RECT 74.120 157.965 74.540 158.165 ;
        RECT 74.715 158.135 74.885 158.385 ;
        RECT 74.715 157.965 75.410 158.135 ;
        RECT 70.495 157.525 71.210 157.695 ;
        RECT 70.495 157.145 70.665 157.525 ;
        RECT 71.380 157.145 71.635 157.720 ;
        RECT 72.450 157.145 72.950 157.755 ;
        RECT 73.580 157.625 74.805 157.795 ;
        RECT 75.580 157.775 75.755 158.385 ;
        RECT 73.580 157.145 73.910 157.625 ;
        RECT 74.475 157.145 74.805 157.625 ;
        RECT 75.415 157.145 75.755 157.775 ;
        RECT 76.845 158.385 77.185 159.355 ;
        RECT 78.690 158.555 79.020 159.355 ;
        RECT 79.820 158.555 80.150 159.355 ;
        RECT 77.715 158.385 80.150 158.555 ;
        RECT 80.900 158.545 81.155 159.215 ;
        RECT 81.800 158.805 82.130 159.315 ;
        RECT 80.900 158.505 81.080 158.545 ;
        RECT 76.845 157.775 77.020 158.385 ;
        RECT 77.715 158.135 77.885 158.385 ;
        RECT 77.190 157.965 77.885 158.135 ;
        RECT 78.060 157.965 78.480 158.165 ;
        RECT 78.650 157.965 78.980 158.165 ;
        RECT 79.150 157.965 79.480 158.165 ;
        RECT 76.845 157.145 77.185 157.775 ;
        RECT 77.795 157.625 79.020 157.795 ;
        RECT 77.795 157.145 78.125 157.625 ;
        RECT 78.690 157.145 79.020 157.625 ;
        RECT 79.650 157.755 79.820 158.385 ;
        RECT 80.815 158.335 81.080 158.505 ;
        RECT 80.005 157.965 80.355 158.215 ;
        RECT 79.650 157.145 80.150 157.755 ;
        RECT 80.900 157.685 81.080 158.335 ;
        RECT 81.800 158.215 82.050 158.805 ;
        RECT 82.400 158.655 82.570 159.265 ;
        RECT 83.300 158.975 83.540 159.265 ;
        RECT 84.340 159.055 84.970 159.305 ;
        RECT 84.340 158.975 84.510 159.055 ;
        RECT 85.940 158.975 86.110 159.265 ;
        RECT 86.910 159.140 87.740 159.310 ;
        RECT 83.300 158.805 84.510 158.975 ;
        RECT 81.250 157.885 82.050 158.215 ;
        RECT 80.900 157.155 81.155 157.685 ;
        RECT 81.800 157.235 82.050 157.885 ;
        RECT 82.250 158.635 82.570 158.655 ;
        RECT 82.250 158.465 84.170 158.635 ;
        RECT 82.250 157.570 82.440 158.465 ;
        RECT 84.340 158.295 84.510 158.805 ;
        RECT 84.680 158.545 85.200 158.855 ;
        RECT 82.610 158.125 84.510 158.295 ;
        RECT 82.610 158.065 82.940 158.125 ;
        RECT 83.090 157.895 83.420 157.955 ;
        RECT 82.760 157.625 83.420 157.895 ;
        RECT 82.250 157.240 82.570 157.570 ;
        RECT 83.610 157.365 83.780 158.125 ;
        RECT 84.680 157.955 84.860 158.365 ;
        RECT 83.950 157.785 84.280 157.905 ;
        RECT 85.030 157.785 85.200 158.545 ;
        RECT 83.950 157.615 85.200 157.785 ;
        RECT 85.370 158.725 86.740 158.975 ;
        RECT 85.370 157.955 85.560 158.725 ;
        RECT 86.490 158.465 86.740 158.725 ;
        RECT 85.730 158.295 85.980 158.455 ;
        RECT 86.910 158.295 87.080 159.140 ;
        RECT 87.975 158.855 88.145 159.355 ;
        RECT 87.250 158.465 87.750 158.845 ;
        RECT 87.975 158.685 88.670 158.855 ;
        RECT 85.730 158.125 87.080 158.295 ;
        RECT 86.660 158.085 87.080 158.125 ;
        RECT 85.370 157.615 85.790 157.955 ;
        RECT 86.080 157.625 86.490 157.955 ;
        RECT 83.610 157.195 84.460 157.365 ;
        RECT 85.540 157.185 85.790 157.615 ;
        RECT 86.660 157.355 86.830 158.085 ;
        RECT 87.000 157.535 87.350 157.905 ;
        RECT 87.530 157.595 87.750 158.465 ;
        RECT 87.920 157.895 88.330 158.515 ;
        RECT 88.500 157.715 88.670 158.685 ;
        RECT 87.975 157.525 88.670 157.715 ;
        RECT 86.660 157.155 87.675 157.355 ;
        RECT 87.975 157.195 88.145 157.525 ;
        RECT 88.860 157.235 89.085 159.355 ;
        RECT 89.755 158.855 89.925 159.355 ;
        RECT 89.260 158.685 89.925 158.855 ;
        RECT 89.260 157.695 89.490 158.685 ;
        RECT 89.660 157.865 90.010 158.515 ;
        RECT 93.385 158.375 93.715 159.355 ;
        RECT 96.165 158.450 96.435 159.355 ;
        RECT 97.115 158.595 97.285 159.355 ;
        RECT 93.385 157.775 93.635 158.375 ;
        RECT 93.805 157.965 94.135 158.215 ;
        RECT 89.260 157.525 89.925 157.695 ;
        RECT 89.755 157.235 89.925 157.525 ;
        RECT 93.385 157.145 93.715 157.775 ;
        RECT 96.165 157.650 96.335 158.450 ;
        RECT 96.620 158.425 97.285 158.595 ;
        RECT 105.455 158.595 105.625 159.355 ;
        RECT 105.455 158.425 106.120 158.595 ;
        RECT 106.305 158.450 106.575 159.355 ;
        RECT 96.620 158.280 96.790 158.425 ;
        RECT 96.505 157.950 96.790 158.280 ;
        RECT 105.950 158.280 106.120 158.425 ;
        RECT 96.620 157.695 96.790 157.950 ;
        RECT 97.025 157.875 97.355 158.245 ;
        RECT 105.385 157.875 105.715 158.245 ;
        RECT 105.950 157.950 106.235 158.280 ;
        RECT 105.950 157.695 106.120 157.950 ;
        RECT 96.165 157.145 96.425 157.650 ;
        RECT 96.620 157.525 97.285 157.695 ;
        RECT 97.115 157.145 97.285 157.525 ;
        RECT 105.455 157.525 106.120 157.695 ;
        RECT 106.405 157.650 106.575 158.450 ;
        RECT 105.455 157.145 105.625 157.525 ;
        RECT 106.315 157.145 106.575 157.650 ;
        RECT 119.815 158.505 119.985 159.355 ;
        RECT 120.655 158.505 120.825 159.355 ;
        RECT 121.415 158.545 121.745 159.355 ;
        RECT 119.815 158.335 120.825 158.505 ;
        RECT 121.030 158.375 121.745 158.545 ;
        RECT 119.815 157.825 120.310 158.335 ;
        RECT 121.030 158.135 121.200 158.375 ;
        RECT 120.700 157.965 121.200 158.135 ;
        RECT 121.370 157.965 121.750 158.205 ;
        RECT 119.815 157.795 120.315 157.825 ;
        RECT 121.030 157.795 121.200 157.965 ;
        RECT 119.815 157.625 120.825 157.795 ;
        RECT 121.030 157.625 121.665 157.795 ;
        RECT 119.815 157.145 119.985 157.625 ;
        RECT 120.655 157.145 120.825 157.625 ;
        RECT 121.495 157.145 121.665 157.625 ;
        RECT 16.960 156.465 17.215 156.625 ;
        RECT 16.875 156.295 17.215 156.465 ;
        RECT 16.960 156.095 17.215 156.295 ;
        RECT 16.960 155.235 17.140 156.095 ;
        RECT 17.860 155.895 18.110 156.545 ;
        RECT 17.310 155.565 18.110 155.895 ;
        RECT 16.960 154.565 17.215 155.235 ;
        RECT 17.860 154.975 18.110 155.565 ;
        RECT 18.310 156.210 18.630 156.540 ;
        RECT 19.670 156.415 20.520 156.585 ;
        RECT 18.310 155.315 18.500 156.210 ;
        RECT 18.820 155.885 19.480 156.155 ;
        RECT 19.150 155.825 19.480 155.885 ;
        RECT 18.670 155.655 19.000 155.715 ;
        RECT 19.670 155.655 19.840 156.415 ;
        RECT 21.600 156.165 21.850 156.595 ;
        RECT 20.010 155.995 21.260 156.165 ;
        RECT 20.010 155.875 20.340 155.995 ;
        RECT 18.670 155.485 20.570 155.655 ;
        RECT 18.310 155.145 20.230 155.315 ;
        RECT 18.310 155.125 18.630 155.145 ;
        RECT 17.860 154.465 18.190 154.975 ;
        RECT 18.460 154.515 18.630 155.125 ;
        RECT 20.400 154.975 20.570 155.485 ;
        RECT 20.740 155.415 20.920 155.825 ;
        RECT 21.090 155.235 21.260 155.995 ;
        RECT 19.360 154.805 20.570 154.975 ;
        RECT 20.740 154.925 21.260 155.235 ;
        RECT 21.430 155.825 21.850 156.165 ;
        RECT 22.720 156.425 23.735 156.625 ;
        RECT 22.140 155.825 22.550 156.155 ;
        RECT 21.430 155.055 21.620 155.825 ;
        RECT 22.720 155.695 22.890 156.425 ;
        RECT 24.035 156.255 24.205 156.585 ;
        RECT 23.060 155.875 23.410 156.245 ;
        RECT 22.720 155.655 23.140 155.695 ;
        RECT 21.790 155.485 23.140 155.655 ;
        RECT 21.790 155.325 22.040 155.485 ;
        RECT 22.550 155.055 22.800 155.315 ;
        RECT 21.430 154.805 22.800 155.055 ;
        RECT 19.360 154.515 19.600 154.805 ;
        RECT 20.400 154.725 20.570 154.805 ;
        RECT 20.400 154.475 21.030 154.725 ;
        RECT 22.000 154.515 22.170 154.805 ;
        RECT 22.970 154.640 23.140 155.485 ;
        RECT 23.590 155.315 23.810 156.185 ;
        RECT 24.035 156.065 24.730 156.255 ;
        RECT 23.310 154.935 23.810 155.315 ;
        RECT 23.980 155.265 24.390 155.885 ;
        RECT 24.560 155.095 24.730 156.065 ;
        RECT 24.035 154.925 24.730 155.095 ;
        RECT 22.970 154.470 23.800 154.640 ;
        RECT 24.035 154.425 24.205 154.925 ;
        RECT 24.920 154.425 25.145 156.545 ;
        RECT 25.815 156.255 25.985 156.545 ;
        RECT 25.320 156.085 25.985 156.255 ;
        RECT 26.245 156.130 26.505 156.635 ;
        RECT 27.195 156.255 27.365 156.635 ;
        RECT 25.320 155.095 25.550 156.085 ;
        RECT 25.720 155.265 26.070 155.915 ;
        RECT 26.245 155.330 26.415 156.130 ;
        RECT 26.700 156.085 27.365 156.255 ;
        RECT 32.340 156.175 32.625 156.635 ;
        RECT 26.700 155.830 26.870 156.085 ;
        RECT 32.340 156.005 33.295 156.175 ;
        RECT 26.585 155.500 26.870 155.830 ;
        RECT 27.105 155.535 27.435 155.905 ;
        RECT 26.700 155.355 26.870 155.500 ;
        RECT 25.320 154.925 25.985 155.095 ;
        RECT 25.815 154.425 25.985 154.925 ;
        RECT 26.245 154.425 26.515 155.330 ;
        RECT 26.700 155.185 27.365 155.355 ;
        RECT 32.225 155.275 32.915 155.835 ;
        RECT 27.195 154.425 27.365 155.185 ;
        RECT 33.085 155.105 33.295 156.005 ;
        RECT 32.340 154.885 33.295 155.105 ;
        RECT 33.465 155.835 33.865 156.635 ;
        RECT 34.055 156.175 34.335 156.635 ;
        RECT 34.055 156.005 35.180 156.175 ;
        RECT 35.350 156.065 35.735 156.635 ;
        RECT 34.730 155.895 35.180 156.005 ;
        RECT 33.465 155.275 34.560 155.835 ;
        RECT 34.730 155.565 35.285 155.895 ;
        RECT 32.340 154.425 32.625 154.885 ;
        RECT 33.465 154.425 33.865 155.275 ;
        RECT 34.730 155.105 35.180 155.565 ;
        RECT 35.455 155.395 35.735 156.065 ;
        RECT 34.055 154.885 35.180 155.105 ;
        RECT 34.055 154.425 34.335 154.885 ;
        RECT 35.350 154.425 35.735 155.395 ;
        RECT 40.045 156.005 40.385 156.635 ;
        RECT 40.995 156.155 41.325 156.635 ;
        RECT 41.890 156.155 42.220 156.635 ;
        RECT 40.045 155.395 40.220 156.005 ;
        RECT 40.995 155.985 42.220 156.155 ;
        RECT 42.850 156.025 43.350 156.635 ;
        RECT 40.390 155.645 41.085 155.815 ;
        RECT 40.915 155.395 41.085 155.645 ;
        RECT 41.260 155.615 41.680 155.815 ;
        RECT 41.850 155.615 42.180 155.815 ;
        RECT 42.350 155.615 42.680 155.815 ;
        RECT 42.850 155.395 43.020 156.025 ;
        RECT 43.725 156.005 44.065 156.635 ;
        RECT 44.675 156.155 45.005 156.635 ;
        RECT 45.570 156.155 45.900 156.635 ;
        RECT 43.205 155.565 43.555 155.815 ;
        RECT 43.725 155.395 43.900 156.005 ;
        RECT 44.675 155.985 45.900 156.155 ;
        RECT 46.530 156.025 47.030 156.635 ;
        RECT 47.610 156.025 48.110 156.635 ;
        RECT 44.070 155.645 44.765 155.815 ;
        RECT 44.940 155.785 45.360 155.815 ;
        RECT 44.595 155.395 44.765 155.645 ;
        RECT 44.935 155.615 45.360 155.785 ;
        RECT 45.530 155.615 45.860 155.815 ;
        RECT 46.030 155.615 46.360 155.815 ;
        RECT 46.530 155.395 46.700 156.025 ;
        RECT 46.885 155.565 47.235 155.815 ;
        RECT 47.405 155.565 47.755 155.815 ;
        RECT 47.940 155.395 48.110 156.025 ;
        RECT 48.740 156.155 49.070 156.635 ;
        RECT 49.635 156.155 49.965 156.635 ;
        RECT 48.740 155.985 49.965 156.155 ;
        RECT 50.575 156.005 50.915 156.635 ;
        RECT 48.280 155.615 48.610 155.815 ;
        RECT 48.780 155.615 49.110 155.815 ;
        RECT 49.280 155.615 49.700 155.815 ;
        RECT 49.875 155.645 50.570 155.815 ;
        RECT 49.875 155.395 50.045 155.645 ;
        RECT 50.740 155.395 50.915 156.005 ;
        RECT 40.045 154.425 40.385 155.395 ;
        RECT 40.915 155.225 43.350 155.395 ;
        RECT 41.890 154.425 42.220 155.225 ;
        RECT 43.020 154.425 43.350 155.225 ;
        RECT 43.725 154.425 44.065 155.395 ;
        RECT 44.595 155.225 47.030 155.395 ;
        RECT 45.570 154.425 45.900 155.225 ;
        RECT 46.700 154.425 47.030 155.225 ;
        RECT 47.610 155.225 50.045 155.395 ;
        RECT 47.610 154.425 47.940 155.225 ;
        RECT 48.740 154.425 49.070 155.225 ;
        RECT 50.575 154.425 50.915 155.395 ;
        RECT 53.760 156.095 54.015 156.625 ;
        RECT 53.760 155.235 53.940 156.095 ;
        RECT 54.660 155.895 54.910 156.545 ;
        RECT 54.110 155.565 54.910 155.895 ;
        RECT 53.760 154.765 54.015 155.235 ;
        RECT 53.675 154.595 54.015 154.765 ;
        RECT 53.760 154.565 54.015 154.595 ;
        RECT 54.660 154.975 54.910 155.565 ;
        RECT 55.110 156.210 55.430 156.540 ;
        RECT 56.470 156.415 57.320 156.585 ;
        RECT 55.110 155.315 55.300 156.210 ;
        RECT 55.620 155.885 56.280 156.155 ;
        RECT 55.950 155.825 56.280 155.885 ;
        RECT 55.470 155.655 55.800 155.715 ;
        RECT 56.470 155.655 56.640 156.415 ;
        RECT 58.400 156.165 58.650 156.595 ;
        RECT 56.810 155.995 58.060 156.165 ;
        RECT 56.810 155.875 57.140 155.995 ;
        RECT 55.470 155.485 57.370 155.655 ;
        RECT 55.110 155.145 57.030 155.315 ;
        RECT 55.110 155.125 55.430 155.145 ;
        RECT 54.660 154.465 54.990 154.975 ;
        RECT 55.260 154.515 55.430 155.125 ;
        RECT 57.200 154.975 57.370 155.485 ;
        RECT 57.540 155.415 57.720 155.825 ;
        RECT 57.890 155.235 58.060 155.995 ;
        RECT 56.160 154.805 57.370 154.975 ;
        RECT 57.540 154.925 58.060 155.235 ;
        RECT 58.230 155.825 58.650 156.165 ;
        RECT 59.520 156.425 60.535 156.625 ;
        RECT 58.940 155.825 59.350 156.155 ;
        RECT 58.230 155.055 58.420 155.825 ;
        RECT 59.520 155.695 59.690 156.425 ;
        RECT 60.835 156.255 61.005 156.585 ;
        RECT 59.860 155.875 60.210 156.245 ;
        RECT 59.520 155.655 59.940 155.695 ;
        RECT 58.590 155.485 59.940 155.655 ;
        RECT 58.590 155.325 58.840 155.485 ;
        RECT 59.350 155.055 59.600 155.315 ;
        RECT 58.230 154.805 59.600 155.055 ;
        RECT 56.160 154.515 56.400 154.805 ;
        RECT 57.200 154.725 57.370 154.805 ;
        RECT 57.200 154.475 57.830 154.725 ;
        RECT 58.800 154.515 58.970 154.805 ;
        RECT 59.770 154.640 59.940 155.485 ;
        RECT 60.390 155.315 60.610 156.185 ;
        RECT 60.835 156.065 61.530 156.255 ;
        RECT 60.110 154.935 60.610 155.315 ;
        RECT 60.780 155.265 61.190 155.885 ;
        RECT 61.360 155.095 61.530 156.065 ;
        RECT 60.835 154.925 61.530 155.095 ;
        RECT 59.770 154.470 60.600 154.640 ;
        RECT 60.835 154.425 61.005 154.925 ;
        RECT 61.720 154.425 61.945 156.545 ;
        RECT 62.615 156.255 62.785 156.545 ;
        RECT 62.120 156.085 62.785 156.255 ;
        RECT 62.120 155.095 62.350 156.085 ;
        RECT 63.945 156.005 64.275 156.635 ;
        RECT 67.285 156.155 67.545 156.610 ;
        RECT 68.155 156.155 68.415 156.610 ;
        RECT 69.015 156.155 69.275 156.610 ;
        RECT 69.875 156.155 70.135 156.610 ;
        RECT 70.720 156.155 70.995 156.610 ;
        RECT 71.580 156.155 71.840 156.610 ;
        RECT 72.440 156.155 72.700 156.610 ;
        RECT 73.300 156.155 73.560 156.610 ;
        RECT 62.520 155.265 62.870 155.915 ;
        RECT 63.525 155.565 63.855 155.815 ;
        RECT 64.025 155.405 64.275 156.005 ;
        RECT 66.815 155.985 73.560 156.155 ;
        RECT 66.815 155.445 67.980 155.985 ;
        RECT 74.160 155.815 74.410 156.625 ;
        RECT 75.020 155.815 75.270 156.625 ;
        RECT 76.130 156.025 76.630 156.635 ;
        RECT 68.150 155.565 75.270 155.815 ;
        RECT 75.925 155.565 76.275 155.815 ;
        RECT 62.120 154.925 62.785 155.095 ;
        RECT 62.615 154.425 62.785 154.925 ;
        RECT 63.945 154.425 64.275 155.405 ;
        RECT 66.785 155.395 67.980 155.445 ;
        RECT 66.785 155.275 73.560 155.395 ;
        RECT 66.815 155.170 73.560 155.275 ;
        RECT 67.255 154.430 67.545 155.170 ;
        RECT 68.155 155.155 73.560 155.170 ;
        RECT 68.155 154.430 68.415 155.155 ;
        RECT 69.015 154.430 69.275 155.155 ;
        RECT 69.875 154.430 70.135 155.155 ;
        RECT 70.720 154.430 70.980 155.155 ;
        RECT 71.580 154.430 71.840 155.155 ;
        RECT 72.440 154.430 72.700 155.155 ;
        RECT 73.300 154.430 73.560 155.155 ;
        RECT 74.160 154.430 74.410 155.565 ;
        RECT 75.025 154.425 75.270 155.565 ;
        RECT 76.460 155.395 76.630 156.025 ;
        RECT 77.260 156.155 77.590 156.635 ;
        RECT 78.155 156.155 78.485 156.635 ;
        RECT 77.260 155.985 78.485 156.155 ;
        RECT 79.095 156.005 79.435 156.635 ;
        RECT 76.800 155.615 77.130 155.815 ;
        RECT 77.300 155.615 77.630 155.815 ;
        RECT 77.800 155.615 78.220 155.815 ;
        RECT 78.395 155.645 79.090 155.815 ;
        RECT 78.395 155.395 78.565 155.645 ;
        RECT 79.260 155.395 79.435 156.005 ;
        RECT 76.130 155.225 78.565 155.395 ;
        RECT 76.130 154.425 76.460 155.225 ;
        RECT 77.260 154.425 77.590 155.225 ;
        RECT 79.095 154.425 79.435 155.395 ;
        RECT 80.525 156.005 80.865 156.635 ;
        RECT 81.475 156.155 81.805 156.635 ;
        RECT 82.370 156.155 82.700 156.635 ;
        RECT 80.525 155.395 80.700 156.005 ;
        RECT 81.475 155.985 82.700 156.155 ;
        RECT 83.330 156.025 83.830 156.635 ;
        RECT 80.870 155.645 81.565 155.815 ;
        RECT 81.395 155.395 81.565 155.645 ;
        RECT 81.740 155.615 82.160 155.815 ;
        RECT 82.330 155.615 82.660 155.815 ;
        RECT 82.830 155.615 83.160 155.815 ;
        RECT 83.330 155.395 83.500 156.025 ;
        RECT 97.545 156.005 97.885 156.635 ;
        RECT 98.495 156.155 98.825 156.635 ;
        RECT 99.390 156.155 99.720 156.635 ;
        RECT 83.685 155.565 84.035 155.815 ;
        RECT 97.545 155.395 97.720 156.005 ;
        RECT 98.495 155.985 99.720 156.155 ;
        RECT 100.350 156.025 100.850 156.635 ;
        RECT 103.730 156.025 104.230 156.635 ;
        RECT 97.890 155.645 98.585 155.815 ;
        RECT 98.415 155.395 98.585 155.645 ;
        RECT 98.760 155.615 99.180 155.815 ;
        RECT 99.350 155.615 99.680 155.815 ;
        RECT 99.850 155.615 100.180 155.815 ;
        RECT 100.350 155.395 100.520 156.025 ;
        RECT 100.705 155.565 101.055 155.815 ;
        RECT 103.525 155.565 103.875 155.815 ;
        RECT 104.060 155.395 104.230 156.025 ;
        RECT 104.860 156.155 105.190 156.635 ;
        RECT 105.755 156.155 106.085 156.635 ;
        RECT 104.860 155.985 106.085 156.155 ;
        RECT 106.695 156.005 107.035 156.635 ;
        RECT 107.410 156.025 107.910 156.635 ;
        RECT 104.400 155.615 104.730 155.815 ;
        RECT 104.900 155.615 105.230 155.815 ;
        RECT 105.400 155.615 105.820 155.815 ;
        RECT 105.995 155.645 106.690 155.815 ;
        RECT 105.995 155.395 106.165 155.645 ;
        RECT 106.860 155.395 107.035 156.005 ;
        RECT 107.205 155.565 107.555 155.815 ;
        RECT 107.740 155.395 107.910 156.025 ;
        RECT 108.540 156.155 108.870 156.635 ;
        RECT 109.435 156.155 109.765 156.635 ;
        RECT 108.540 155.985 109.765 156.155 ;
        RECT 110.375 156.005 110.715 156.635 ;
        RECT 108.080 155.615 108.410 155.815 ;
        RECT 108.580 155.615 108.910 155.815 ;
        RECT 109.080 155.615 109.500 155.815 ;
        RECT 109.675 155.645 110.370 155.815 ;
        RECT 109.675 155.395 109.845 155.645 ;
        RECT 110.540 155.395 110.715 156.005 ;
        RECT 80.525 154.425 80.865 155.395 ;
        RECT 81.395 155.225 83.830 155.395 ;
        RECT 82.370 154.425 82.700 155.225 ;
        RECT 83.500 154.425 83.830 155.225 ;
        RECT 97.545 154.425 97.885 155.395 ;
        RECT 98.415 155.225 100.850 155.395 ;
        RECT 99.390 154.425 99.720 155.225 ;
        RECT 100.520 154.425 100.850 155.225 ;
        RECT 103.730 155.225 106.165 155.395 ;
        RECT 103.730 154.425 104.060 155.225 ;
        RECT 104.860 154.425 105.190 155.225 ;
        RECT 106.695 154.425 107.035 155.395 ;
        RECT 107.410 155.225 109.845 155.395 ;
        RECT 107.410 154.425 107.740 155.225 ;
        RECT 108.540 154.425 108.870 155.225 ;
        RECT 110.375 154.425 110.715 155.395 ;
        RECT 110.885 156.005 111.225 156.635 ;
        RECT 111.835 156.155 112.165 156.635 ;
        RECT 112.730 156.155 113.060 156.635 ;
        RECT 110.885 155.395 111.060 156.005 ;
        RECT 111.835 155.985 113.060 156.155 ;
        RECT 113.690 156.025 114.190 156.635 ;
        RECT 116.495 156.155 116.665 156.635 ;
        RECT 117.335 156.155 117.505 156.635 ;
        RECT 118.175 156.155 118.345 156.635 ;
        RECT 111.230 155.645 111.925 155.815 ;
        RECT 111.755 155.395 111.925 155.645 ;
        RECT 112.100 155.615 112.520 155.815 ;
        RECT 112.690 155.615 113.020 155.815 ;
        RECT 113.190 155.615 113.520 155.815 ;
        RECT 113.690 155.395 113.860 156.025 ;
        RECT 116.495 155.985 117.130 156.155 ;
        RECT 117.335 155.985 118.345 156.155 ;
        RECT 116.960 155.815 117.130 155.985 ;
        RECT 114.045 155.565 114.395 155.815 ;
        RECT 116.410 155.575 116.790 155.815 ;
        RECT 116.960 155.645 117.460 155.815 ;
        RECT 116.960 155.405 117.130 155.645 ;
        RECT 117.850 155.445 118.345 155.985 ;
        RECT 110.885 154.425 111.225 155.395 ;
        RECT 111.755 155.225 114.190 155.395 ;
        RECT 112.730 154.425 113.060 155.225 ;
        RECT 113.860 154.425 114.190 155.225 ;
        RECT 116.415 155.235 117.130 155.405 ;
        RECT 117.335 155.275 118.345 155.445 ;
        RECT 116.415 154.425 116.745 155.235 ;
        RECT 117.335 154.425 117.505 155.275 ;
        RECT 118.175 154.425 118.345 155.275 ;
        RECT 21.355 153.745 23.385 153.915 ;
        RECT 20.265 153.325 20.780 153.735 ;
        RECT 20.265 152.515 20.605 153.325 ;
        RECT 21.355 153.080 21.525 153.745 ;
        RECT 21.920 153.405 23.045 153.575 ;
        RECT 20.775 152.890 21.525 153.080 ;
        RECT 21.695 153.065 22.705 153.235 ;
        RECT 20.265 152.345 21.495 152.515 ;
        RECT 20.540 151.740 20.785 152.345 ;
        RECT 21.695 151.705 21.885 153.065 ;
        RECT 22.055 152.045 22.330 152.865 ;
        RECT 22.535 152.265 22.705 153.065 ;
        RECT 22.875 152.275 23.045 153.405 ;
        RECT 23.215 152.775 23.385 153.745 ;
        RECT 23.895 152.945 24.230 153.915 ;
        RECT 23.215 152.445 23.410 152.775 ;
        RECT 23.635 152.445 23.890 152.775 ;
        RECT 23.635 152.275 23.805 152.445 ;
        RECT 24.060 152.275 24.230 152.945 ;
        RECT 31.285 152.935 31.615 153.915 ;
        RECT 32.315 153.155 32.485 153.915 ;
        RECT 32.315 152.985 32.980 153.155 ;
        RECT 33.165 153.010 33.435 153.915 ;
        RECT 30.865 152.525 31.195 152.775 ;
        RECT 31.365 152.335 31.615 152.935 ;
        RECT 32.810 152.840 32.980 152.985 ;
        RECT 32.245 152.435 32.575 152.805 ;
        RECT 32.810 152.510 33.095 152.840 ;
        RECT 22.875 152.105 23.805 152.275 ;
        RECT 22.875 152.070 23.050 152.105 ;
        RECT 22.055 151.875 22.335 152.045 ;
        RECT 22.055 151.705 22.330 151.875 ;
        RECT 22.520 151.705 23.050 152.070 ;
        RECT 23.975 151.705 24.230 152.275 ;
        RECT 31.285 151.705 31.615 152.335 ;
        RECT 32.810 152.255 32.980 152.510 ;
        RECT 32.315 152.085 32.980 152.255 ;
        RECT 33.265 152.210 33.435 153.010 ;
        RECT 32.315 151.705 32.485 152.085 ;
        RECT 33.175 151.705 33.435 152.210 ;
        RECT 33.610 152.945 33.945 153.915 ;
        RECT 34.455 153.745 36.485 153.915 ;
        RECT 33.610 152.275 33.780 152.945 ;
        RECT 34.455 152.775 34.625 153.745 ;
        RECT 33.950 152.445 34.205 152.775 ;
        RECT 34.430 152.445 34.625 152.775 ;
        RECT 34.795 153.405 35.920 153.575 ;
        RECT 34.035 152.275 34.205 152.445 ;
        RECT 34.795 152.275 34.965 153.405 ;
        RECT 33.610 151.705 33.865 152.275 ;
        RECT 34.035 152.105 34.965 152.275 ;
        RECT 35.135 153.065 36.145 153.235 ;
        RECT 35.135 152.265 35.305 153.065 ;
        RECT 35.510 152.725 35.785 152.865 ;
        RECT 35.505 152.555 35.785 152.725 ;
        RECT 34.790 152.070 34.965 152.105 ;
        RECT 34.790 151.705 35.320 152.070 ;
        RECT 35.510 151.705 35.785 152.555 ;
        RECT 35.955 151.705 36.145 153.065 ;
        RECT 36.315 153.080 36.485 153.745 ;
        RECT 37.060 153.325 37.575 153.735 ;
        RECT 36.315 152.890 37.065 153.080 ;
        RECT 37.235 152.515 37.575 153.325 ;
        RECT 36.345 152.345 37.575 152.515 ;
        RECT 37.745 152.945 38.085 153.915 ;
        RECT 39.590 153.115 39.920 153.915 ;
        RECT 40.720 153.115 41.050 153.915 ;
        RECT 38.615 152.945 41.050 153.115 ;
        RECT 37.055 151.740 37.300 152.345 ;
        RECT 37.745 152.335 37.920 152.945 ;
        RECT 38.615 152.695 38.785 152.945 ;
        RECT 38.090 152.525 38.785 152.695 ;
        RECT 38.960 152.525 39.380 152.725 ;
        RECT 39.550 152.525 39.880 152.725 ;
        RECT 40.050 152.525 40.380 152.725 ;
        RECT 37.745 151.705 38.085 152.335 ;
        RECT 38.695 152.185 39.920 152.355 ;
        RECT 38.695 151.705 39.025 152.185 ;
        RECT 39.590 151.705 39.920 152.185 ;
        RECT 40.550 152.315 40.720 152.945 ;
        RECT 57.505 152.935 57.835 153.915 ;
        RECT 40.905 152.525 41.255 152.775 ;
        RECT 57.085 152.525 57.415 152.775 ;
        RECT 57.585 152.335 57.835 152.935 ;
        RECT 40.550 151.705 41.050 152.315 ;
        RECT 57.505 151.705 57.835 152.335 ;
        RECT 58.820 153.105 59.075 153.775 ;
        RECT 59.720 153.365 60.050 153.875 ;
        RECT 58.820 152.245 59.000 153.105 ;
        RECT 59.720 152.775 59.970 153.365 ;
        RECT 60.320 153.215 60.490 153.825 ;
        RECT 61.220 153.535 61.460 153.825 ;
        RECT 62.260 153.615 62.890 153.865 ;
        RECT 62.260 153.535 62.430 153.615 ;
        RECT 63.860 153.535 64.030 153.825 ;
        RECT 64.830 153.700 65.660 153.870 ;
        RECT 61.220 153.365 62.430 153.535 ;
        RECT 59.170 152.445 59.970 152.775 ;
        RECT 58.820 152.045 59.075 152.245 ;
        RECT 58.735 151.875 59.075 152.045 ;
        RECT 58.820 151.715 59.075 151.875 ;
        RECT 59.720 151.795 59.970 152.445 ;
        RECT 60.170 153.195 60.490 153.215 ;
        RECT 60.170 153.025 62.090 153.195 ;
        RECT 60.170 152.130 60.360 153.025 ;
        RECT 62.260 152.855 62.430 153.365 ;
        RECT 62.600 153.105 63.120 153.415 ;
        RECT 60.530 152.685 62.430 152.855 ;
        RECT 60.530 152.625 60.860 152.685 ;
        RECT 61.010 152.455 61.340 152.515 ;
        RECT 60.680 152.185 61.340 152.455 ;
        RECT 60.170 151.800 60.490 152.130 ;
        RECT 61.530 151.925 61.700 152.685 ;
        RECT 62.600 152.515 62.780 152.925 ;
        RECT 61.870 152.345 62.200 152.465 ;
        RECT 62.950 152.345 63.120 153.105 ;
        RECT 61.870 152.175 63.120 152.345 ;
        RECT 63.290 153.285 64.660 153.535 ;
        RECT 63.290 152.515 63.480 153.285 ;
        RECT 64.410 153.025 64.660 153.285 ;
        RECT 63.650 152.855 63.900 153.015 ;
        RECT 64.830 152.855 65.000 153.700 ;
        RECT 65.895 153.415 66.065 153.915 ;
        RECT 65.170 153.025 65.670 153.405 ;
        RECT 65.895 153.245 66.590 153.415 ;
        RECT 63.650 152.685 65.000 152.855 ;
        RECT 64.580 152.645 65.000 152.685 ;
        RECT 63.290 152.175 63.710 152.515 ;
        RECT 64.000 152.185 64.410 152.515 ;
        RECT 61.530 151.755 62.380 151.925 ;
        RECT 63.460 151.745 63.710 152.175 ;
        RECT 64.580 151.915 64.750 152.645 ;
        RECT 64.920 152.095 65.270 152.465 ;
        RECT 65.450 152.155 65.670 153.025 ;
        RECT 65.840 152.455 66.250 153.075 ;
        RECT 66.420 152.275 66.590 153.245 ;
        RECT 65.895 152.085 66.590 152.275 ;
        RECT 64.580 151.715 65.595 151.915 ;
        RECT 65.895 151.755 66.065 152.085 ;
        RECT 66.780 151.795 67.005 153.915 ;
        RECT 67.675 153.415 67.845 153.915 ;
        RECT 67.180 153.245 67.845 153.415 ;
        RECT 67.180 152.255 67.410 153.245 ;
        RECT 71.415 153.155 71.585 153.915 ;
        RECT 67.580 152.425 67.930 153.075 ;
        RECT 71.415 152.985 72.130 153.155 ;
        RECT 72.300 153.010 72.555 153.915 ;
        RECT 71.325 152.435 71.680 152.805 ;
        RECT 71.960 152.775 72.130 152.985 ;
        RECT 71.960 152.445 72.215 152.775 ;
        RECT 71.960 152.255 72.130 152.445 ;
        RECT 72.385 152.280 72.555 153.010 ;
        RECT 73.685 152.775 73.855 153.700 ;
        RECT 74.025 153.495 74.355 153.895 ;
        RECT 75.055 153.495 75.755 153.915 ;
        RECT 74.025 153.265 75.755 153.495 ;
        RECT 74.025 153.045 74.355 153.265 ;
        RECT 74.550 152.775 74.875 153.065 ;
        RECT 73.165 152.445 73.475 152.775 ;
        RECT 73.685 152.445 74.060 152.775 ;
        RECT 74.380 152.445 74.875 152.775 ;
        RECT 75.050 152.525 75.380 153.065 ;
        RECT 75.550 152.295 75.755 153.265 ;
        RECT 91.085 152.935 91.415 153.915 ;
        RECT 90.665 152.525 90.995 152.775 ;
        RECT 91.165 152.335 91.415 152.935 ;
        RECT 67.180 152.085 67.845 152.255 ;
        RECT 67.675 151.795 67.845 152.085 ;
        RECT 71.415 152.085 72.130 152.255 ;
        RECT 71.415 151.705 71.585 152.085 ;
        RECT 72.300 151.705 72.555 152.280 ;
        RECT 73.175 152.065 74.535 152.275 ;
        RECT 73.175 151.705 73.505 152.065 ;
        RECT 74.205 151.705 74.535 152.065 ;
        RECT 75.045 151.705 75.755 152.295 ;
        RECT 91.085 151.705 91.415 152.335 ;
        RECT 105.365 152.945 105.705 153.915 ;
        RECT 107.210 153.115 107.540 153.915 ;
        RECT 108.340 153.115 108.670 153.915 ;
        RECT 106.235 152.945 108.670 153.115 ;
        RECT 109.045 152.945 109.385 153.915 ;
        RECT 110.890 153.115 111.220 153.915 ;
        RECT 112.020 153.115 112.350 153.915 ;
        RECT 109.915 152.945 112.350 153.115 ;
        RECT 105.365 152.335 105.540 152.945 ;
        RECT 106.235 152.695 106.405 152.945 ;
        RECT 105.710 152.525 106.405 152.695 ;
        RECT 106.580 152.525 107.000 152.725 ;
        RECT 107.170 152.525 107.500 152.725 ;
        RECT 107.670 152.525 108.000 152.725 ;
        RECT 105.365 151.705 105.705 152.335 ;
        RECT 106.315 152.185 107.540 152.355 ;
        RECT 106.315 151.705 106.645 152.185 ;
        RECT 107.210 151.705 107.540 152.185 ;
        RECT 108.170 152.315 108.340 152.945 ;
        RECT 108.525 152.525 108.875 152.775 ;
        RECT 109.045 152.335 109.220 152.945 ;
        RECT 109.915 152.695 110.085 152.945 ;
        RECT 109.390 152.525 110.085 152.695 ;
        RECT 110.260 152.525 110.680 152.725 ;
        RECT 110.850 152.525 111.180 152.725 ;
        RECT 111.350 152.525 111.680 152.725 ;
        RECT 108.170 151.705 108.670 152.315 ;
        RECT 109.045 151.705 109.385 152.335 ;
        RECT 109.995 152.185 111.220 152.355 ;
        RECT 109.995 151.705 110.325 152.185 ;
        RECT 110.890 151.705 111.220 152.185 ;
        RECT 111.850 152.315 112.020 152.945 ;
        RECT 119.145 152.935 119.475 153.915 ;
        RECT 120.635 153.155 120.805 153.915 ;
        RECT 120.635 152.985 121.300 153.155 ;
        RECT 121.485 153.010 121.755 153.915 ;
        RECT 112.205 152.525 112.555 152.775 ;
        RECT 119.145 152.335 119.395 152.935 ;
        RECT 121.130 152.840 121.300 152.985 ;
        RECT 119.565 152.525 119.895 152.775 ;
        RECT 120.565 152.435 120.895 152.805 ;
        RECT 121.130 152.510 121.415 152.840 ;
        RECT 111.850 151.705 112.350 152.315 ;
        RECT 119.145 151.705 119.475 152.335 ;
        RECT 121.130 152.255 121.300 152.510 ;
        RECT 120.635 152.085 121.300 152.255 ;
        RECT 121.585 152.210 121.755 153.010 ;
        RECT 120.635 151.705 120.805 152.085 ;
        RECT 121.495 151.705 121.755 152.210 ;
        RECT 16.500 150.655 16.755 151.185 ;
        RECT 16.500 149.795 16.680 150.655 ;
        RECT 17.400 150.455 17.650 151.105 ;
        RECT 16.850 150.125 17.650 150.455 ;
        RECT 16.500 149.325 16.755 149.795 ;
        RECT 16.415 149.155 16.755 149.325 ;
        RECT 16.500 149.125 16.755 149.155 ;
        RECT 17.400 149.535 17.650 150.125 ;
        RECT 17.850 150.770 18.170 151.100 ;
        RECT 19.210 150.975 20.060 151.145 ;
        RECT 17.850 149.875 18.040 150.770 ;
        RECT 18.360 150.445 19.020 150.715 ;
        RECT 18.690 150.385 19.020 150.445 ;
        RECT 18.210 150.215 18.540 150.275 ;
        RECT 19.210 150.215 19.380 150.975 ;
        RECT 21.140 150.725 21.390 151.155 ;
        RECT 19.550 150.555 20.800 150.725 ;
        RECT 19.550 150.435 19.880 150.555 ;
        RECT 18.210 150.045 20.110 150.215 ;
        RECT 17.850 149.705 19.770 149.875 ;
        RECT 17.850 149.685 18.170 149.705 ;
        RECT 17.400 149.025 17.730 149.535 ;
        RECT 18.000 149.075 18.170 149.685 ;
        RECT 19.940 149.535 20.110 150.045 ;
        RECT 20.280 149.975 20.460 150.385 ;
        RECT 20.630 149.795 20.800 150.555 ;
        RECT 18.900 149.365 20.110 149.535 ;
        RECT 20.280 149.485 20.800 149.795 ;
        RECT 20.970 150.385 21.390 150.725 ;
        RECT 22.260 150.985 23.275 151.185 ;
        RECT 21.680 150.385 22.090 150.715 ;
        RECT 20.970 149.615 21.160 150.385 ;
        RECT 22.260 150.255 22.430 150.985 ;
        RECT 23.575 150.815 23.745 151.145 ;
        RECT 22.600 150.435 22.950 150.805 ;
        RECT 22.260 150.215 22.680 150.255 ;
        RECT 21.330 150.045 22.680 150.215 ;
        RECT 21.330 149.885 21.580 150.045 ;
        RECT 22.090 149.615 22.340 149.875 ;
        RECT 20.970 149.365 22.340 149.615 ;
        RECT 18.900 149.075 19.140 149.365 ;
        RECT 19.940 149.285 20.110 149.365 ;
        RECT 19.940 149.035 20.570 149.285 ;
        RECT 21.540 149.075 21.710 149.365 ;
        RECT 22.510 149.200 22.680 150.045 ;
        RECT 23.130 149.875 23.350 150.745 ;
        RECT 23.575 150.625 24.270 150.815 ;
        RECT 22.850 149.495 23.350 149.875 ;
        RECT 23.520 149.825 23.930 150.445 ;
        RECT 24.100 149.655 24.270 150.625 ;
        RECT 23.575 149.485 24.270 149.655 ;
        RECT 22.510 149.030 23.340 149.200 ;
        RECT 23.575 148.985 23.745 149.485 ;
        RECT 24.460 148.985 24.685 151.105 ;
        RECT 25.355 150.815 25.525 151.105 ;
        RECT 28.000 151.025 28.255 151.185 ;
        RECT 27.915 150.855 28.255 151.025 ;
        RECT 24.860 150.645 25.525 150.815 ;
        RECT 28.000 150.655 28.255 150.855 ;
        RECT 24.860 149.655 25.090 150.645 ;
        RECT 25.260 149.825 25.610 150.475 ;
        RECT 28.000 149.795 28.180 150.655 ;
        RECT 28.900 150.455 29.150 151.105 ;
        RECT 28.350 150.125 29.150 150.455 ;
        RECT 24.860 149.485 25.525 149.655 ;
        RECT 25.355 148.985 25.525 149.485 ;
        RECT 28.000 149.125 28.255 149.795 ;
        RECT 28.900 149.535 29.150 150.125 ;
        RECT 29.350 150.770 29.670 151.100 ;
        RECT 30.710 150.975 31.560 151.145 ;
        RECT 29.350 149.875 29.540 150.770 ;
        RECT 29.860 150.445 30.520 150.715 ;
        RECT 30.190 150.385 30.520 150.445 ;
        RECT 29.710 150.215 30.040 150.275 ;
        RECT 30.710 150.215 30.880 150.975 ;
        RECT 32.640 150.725 32.890 151.155 ;
        RECT 31.050 150.555 32.300 150.725 ;
        RECT 31.050 150.435 31.380 150.555 ;
        RECT 29.710 150.045 31.610 150.215 ;
        RECT 29.350 149.705 31.270 149.875 ;
        RECT 29.350 149.685 29.670 149.705 ;
        RECT 28.900 149.025 29.230 149.535 ;
        RECT 29.500 149.075 29.670 149.685 ;
        RECT 31.440 149.535 31.610 150.045 ;
        RECT 31.780 149.975 31.960 150.385 ;
        RECT 32.130 149.795 32.300 150.555 ;
        RECT 30.400 149.365 31.610 149.535 ;
        RECT 31.780 149.485 32.300 149.795 ;
        RECT 32.470 150.385 32.890 150.725 ;
        RECT 33.760 150.985 34.775 151.185 ;
        RECT 33.180 150.385 33.590 150.715 ;
        RECT 32.470 149.615 32.660 150.385 ;
        RECT 33.760 150.255 33.930 150.985 ;
        RECT 35.075 150.815 35.245 151.145 ;
        RECT 34.100 150.435 34.450 150.805 ;
        RECT 33.760 150.215 34.180 150.255 ;
        RECT 32.830 150.045 34.180 150.215 ;
        RECT 32.830 149.885 33.080 150.045 ;
        RECT 33.590 149.615 33.840 149.875 ;
        RECT 32.470 149.365 33.840 149.615 ;
        RECT 30.400 149.075 30.640 149.365 ;
        RECT 31.440 149.285 31.610 149.365 ;
        RECT 31.440 149.035 32.070 149.285 ;
        RECT 33.040 149.075 33.210 149.365 ;
        RECT 34.010 149.200 34.180 150.045 ;
        RECT 34.630 149.875 34.850 150.745 ;
        RECT 35.075 150.625 35.770 150.815 ;
        RECT 34.350 149.495 34.850 149.875 ;
        RECT 35.020 149.825 35.430 150.445 ;
        RECT 35.600 149.655 35.770 150.625 ;
        RECT 35.075 149.485 35.770 149.655 ;
        RECT 34.010 149.030 34.840 149.200 ;
        RECT 35.075 148.985 35.245 149.485 ;
        RECT 35.960 148.985 36.185 151.105 ;
        RECT 36.855 150.815 37.025 151.105 ;
        RECT 36.360 150.645 37.025 150.815 ;
        RECT 36.360 149.655 36.590 150.645 ;
        RECT 41.170 150.585 41.670 151.195 ;
        RECT 36.760 149.825 37.110 150.475 ;
        RECT 40.965 150.125 41.315 150.375 ;
        RECT 41.500 149.955 41.670 150.585 ;
        RECT 42.300 150.715 42.630 151.195 ;
        RECT 43.195 150.715 43.525 151.195 ;
        RECT 42.300 150.545 43.525 150.715 ;
        RECT 44.135 150.565 44.475 151.195 ;
        RECT 46.565 150.795 46.735 151.145 ;
        RECT 47.435 150.795 47.605 151.145 ;
        RECT 41.840 150.175 42.170 150.375 ;
        RECT 42.340 150.175 42.670 150.375 ;
        RECT 42.840 150.175 43.260 150.375 ;
        RECT 43.435 150.205 44.130 150.375 ;
        RECT 43.435 149.955 43.605 150.205 ;
        RECT 44.300 149.955 44.475 150.565 ;
        RECT 46.030 150.125 46.380 150.695 ;
        RECT 46.565 150.625 48.175 150.795 ;
        RECT 48.345 150.690 48.615 151.035 ;
        RECT 49.325 150.795 49.495 151.145 ;
        RECT 50.195 150.795 50.365 151.145 ;
        RECT 48.005 150.455 48.175 150.625 ;
        RECT 41.170 149.785 43.605 149.955 ;
        RECT 36.360 149.485 37.025 149.655 ;
        RECT 36.855 148.985 37.025 149.485 ;
        RECT 41.170 148.985 41.500 149.785 ;
        RECT 42.300 148.985 42.630 149.785 ;
        RECT 44.135 148.985 44.475 149.955 ;
        RECT 46.030 149.665 46.350 149.955 ;
        RECT 46.550 149.835 47.260 150.455 ;
        RECT 47.430 150.125 47.835 150.455 ;
        RECT 48.005 150.125 48.275 150.455 ;
        RECT 48.005 149.955 48.175 150.125 ;
        RECT 48.445 149.955 48.615 150.690 ;
        RECT 48.790 150.125 49.140 150.695 ;
        RECT 49.325 150.625 50.935 150.795 ;
        RECT 51.105 150.690 51.375 151.035 ;
        RECT 50.765 150.455 50.935 150.625 ;
        RECT 47.450 149.785 48.175 149.955 ;
        RECT 47.450 149.665 47.620 149.785 ;
        RECT 46.030 149.495 47.620 149.665 ;
        RECT 46.030 149.035 47.685 149.325 ;
        RECT 48.345 148.985 48.615 149.955 ;
        RECT 48.790 149.665 49.110 149.955 ;
        RECT 49.310 149.835 50.020 150.455 ;
        RECT 50.190 150.125 50.595 150.455 ;
        RECT 50.765 150.125 51.035 150.455 ;
        RECT 50.765 149.955 50.935 150.125 ;
        RECT 51.205 149.955 51.375 150.690 ;
        RECT 50.210 149.785 50.935 149.955 ;
        RECT 50.210 149.665 50.380 149.785 ;
        RECT 48.790 149.495 50.380 149.665 ;
        RECT 48.790 149.035 50.445 149.325 ;
        RECT 51.105 148.985 51.375 149.955 ;
        RECT 51.545 150.565 51.885 151.195 ;
        RECT 52.495 150.715 52.825 151.195 ;
        RECT 53.390 150.715 53.720 151.195 ;
        RECT 51.545 150.005 51.720 150.565 ;
        RECT 52.495 150.545 53.720 150.715 ;
        RECT 54.350 150.585 54.850 151.195 ;
        RECT 51.890 150.205 52.585 150.375 ;
        RECT 51.545 149.955 51.775 150.005 ;
        RECT 52.415 149.955 52.585 150.205 ;
        RECT 52.760 150.175 53.180 150.375 ;
        RECT 53.350 150.175 53.680 150.375 ;
        RECT 53.850 150.175 54.180 150.375 ;
        RECT 54.350 149.955 54.520 150.585 ;
        RECT 57.800 150.555 58.045 151.160 ;
        RECT 57.525 150.385 58.755 150.555 ;
        RECT 54.705 150.125 55.055 150.375 ;
        RECT 51.545 148.985 51.885 149.955 ;
        RECT 52.415 149.785 54.850 149.955 ;
        RECT 53.390 148.985 53.720 149.785 ;
        RECT 54.520 148.985 54.850 149.785 ;
        RECT 57.525 149.575 57.865 150.385 ;
        RECT 58.035 149.820 58.785 150.010 ;
        RECT 57.525 149.165 58.040 149.575 ;
        RECT 58.615 149.155 58.785 149.820 ;
        RECT 58.955 149.835 59.145 151.195 ;
        RECT 59.315 150.345 59.590 151.195 ;
        RECT 59.780 150.830 60.310 151.195 ;
        RECT 60.135 150.795 60.310 150.830 ;
        RECT 59.315 150.175 59.595 150.345 ;
        RECT 59.315 150.035 59.590 150.175 ;
        RECT 59.795 149.835 59.965 150.635 ;
        RECT 58.955 149.665 59.965 149.835 ;
        RECT 60.135 150.625 61.065 150.795 ;
        RECT 61.235 150.625 61.490 151.195 ;
        RECT 60.135 149.495 60.305 150.625 ;
        RECT 60.895 150.455 61.065 150.625 ;
        RECT 59.180 149.325 60.305 149.495 ;
        RECT 60.475 150.125 60.670 150.455 ;
        RECT 60.895 150.125 61.150 150.455 ;
        RECT 60.475 149.155 60.645 150.125 ;
        RECT 61.320 149.955 61.490 150.625 ;
        RECT 58.615 148.985 60.645 149.155 ;
        RECT 61.155 148.985 61.490 149.955 ;
        RECT 61.665 150.690 61.925 151.195 ;
        RECT 62.615 150.815 62.785 151.195 ;
        RECT 61.665 149.890 61.835 150.690 ;
        RECT 62.120 150.645 62.785 150.815 ;
        RECT 64.055 150.815 64.225 151.195 ;
        RECT 64.055 150.645 64.720 150.815 ;
        RECT 64.915 150.690 65.175 151.195 ;
        RECT 62.120 150.390 62.290 150.645 ;
        RECT 62.005 150.060 62.290 150.390 ;
        RECT 62.525 150.095 62.855 150.465 ;
        RECT 63.985 150.095 64.315 150.465 ;
        RECT 64.550 150.390 64.720 150.645 ;
        RECT 62.120 149.915 62.290 150.060 ;
        RECT 64.550 150.060 64.835 150.390 ;
        RECT 64.550 149.915 64.720 150.060 ;
        RECT 61.665 148.985 61.935 149.890 ;
        RECT 62.120 149.745 62.785 149.915 ;
        RECT 62.615 148.985 62.785 149.745 ;
        RECT 64.055 149.745 64.720 149.915 ;
        RECT 65.005 149.890 65.175 150.690 ;
        RECT 67.735 150.815 67.905 151.195 ;
        RECT 67.735 150.645 68.450 150.815 ;
        RECT 67.645 150.095 68.000 150.465 ;
        RECT 68.280 150.455 68.450 150.645 ;
        RECT 68.620 150.620 68.875 151.195 ;
        RECT 68.280 150.125 68.535 150.455 ;
        RECT 68.280 149.915 68.450 150.125 ;
        RECT 64.055 148.985 64.225 149.745 ;
        RECT 64.905 148.985 65.175 149.890 ;
        RECT 67.735 149.745 68.450 149.915 ;
        RECT 68.705 149.890 68.875 150.620 ;
        RECT 67.735 148.985 67.905 149.745 ;
        RECT 68.620 148.985 68.875 149.890 ;
        RECT 69.925 150.620 70.180 151.195 ;
        RECT 70.895 150.815 71.065 151.195 ;
        RECT 70.350 150.645 71.065 150.815 ;
        RECT 71.835 150.715 72.095 151.105 ;
        RECT 72.695 150.715 72.990 151.105 ;
        RECT 73.615 150.865 73.915 151.195 ;
        RECT 69.925 149.890 70.095 150.620 ;
        RECT 70.350 150.455 70.520 150.645 ;
        RECT 71.340 150.545 72.990 150.715 ;
        RECT 70.265 150.125 70.520 150.455 ;
        RECT 70.350 149.915 70.520 150.125 ;
        RECT 70.800 150.095 71.155 150.465 ;
        RECT 71.340 150.035 71.745 150.545 ;
        RECT 71.915 150.205 73.055 150.375 ;
        RECT 69.925 148.985 70.180 149.890 ;
        RECT 70.350 149.745 71.065 149.915 ;
        RECT 71.340 149.865 72.095 150.035 ;
        RECT 70.895 148.985 71.065 149.745 ;
        RECT 71.835 149.615 72.095 149.865 ;
        RECT 72.885 149.955 73.055 150.205 ;
        RECT 73.225 150.125 73.575 150.695 ;
        RECT 73.745 149.955 73.915 150.865 ;
        RECT 72.885 149.785 73.915 149.955 ;
        RECT 71.835 149.445 72.955 149.615 ;
        RECT 71.835 148.985 72.095 149.445 ;
        RECT 72.695 148.985 72.955 149.445 ;
        RECT 73.605 148.985 73.915 149.785 ;
        RECT 75.005 150.865 75.305 151.195 ;
        RECT 75.005 149.955 75.175 150.865 ;
        RECT 75.930 150.715 76.225 151.105 ;
        RECT 76.825 150.715 77.085 151.105 ;
        RECT 78.305 150.795 78.475 151.145 ;
        RECT 79.175 150.795 79.345 151.145 ;
        RECT 75.345 150.125 75.695 150.695 ;
        RECT 75.930 150.545 77.580 150.715 ;
        RECT 75.865 150.205 77.005 150.375 ;
        RECT 75.865 149.955 76.035 150.205 ;
        RECT 77.175 150.035 77.580 150.545 ;
        RECT 77.770 150.125 78.120 150.695 ;
        RECT 78.305 150.625 79.915 150.795 ;
        RECT 80.085 150.690 80.355 151.035 ;
        RECT 79.745 150.455 79.915 150.625 ;
        RECT 75.005 149.785 76.035 149.955 ;
        RECT 76.825 149.865 77.580 150.035 ;
        RECT 78.290 150.005 79.000 150.455 ;
        RECT 79.170 150.125 79.575 150.455 ;
        RECT 79.745 150.125 80.015 150.455 ;
        RECT 75.005 148.985 75.315 149.785 ;
        RECT 76.825 149.615 77.085 149.865 ;
        RECT 75.965 149.445 77.085 149.615 ;
        RECT 77.770 149.665 78.090 149.955 ;
        RECT 78.285 149.835 79.000 150.005 ;
        RECT 79.745 149.955 79.915 150.125 ;
        RECT 80.185 149.955 80.355 150.690 ;
        RECT 84.940 150.555 85.185 151.160 ;
        RECT 79.190 149.785 79.915 149.955 ;
        RECT 79.190 149.665 79.360 149.785 ;
        RECT 77.770 149.495 79.360 149.665 ;
        RECT 75.965 148.985 76.225 149.445 ;
        RECT 76.825 148.985 77.085 149.445 ;
        RECT 77.770 149.035 79.425 149.325 ;
        RECT 80.085 148.985 80.355 149.955 ;
        RECT 84.665 150.385 85.895 150.555 ;
        RECT 84.665 149.575 85.005 150.385 ;
        RECT 85.175 149.820 85.925 150.010 ;
        RECT 84.665 149.165 85.180 149.575 ;
        RECT 85.755 149.155 85.925 149.820 ;
        RECT 86.095 149.835 86.285 151.195 ;
        RECT 86.455 150.345 86.730 151.195 ;
        RECT 86.920 150.830 87.450 151.195 ;
        RECT 87.275 150.795 87.450 150.830 ;
        RECT 86.455 150.175 86.735 150.345 ;
        RECT 86.455 150.035 86.730 150.175 ;
        RECT 86.935 149.835 87.105 150.635 ;
        RECT 86.095 149.665 87.105 149.835 ;
        RECT 87.275 150.625 88.205 150.795 ;
        RECT 88.375 150.625 88.630 151.195 ;
        RECT 89.355 150.815 89.525 151.105 ;
        RECT 89.355 150.645 90.020 150.815 ;
        RECT 87.275 149.495 87.445 150.625 ;
        RECT 88.035 150.455 88.205 150.625 ;
        RECT 86.320 149.325 87.445 149.495 ;
        RECT 87.615 150.125 87.810 150.455 ;
        RECT 88.035 150.125 88.290 150.455 ;
        RECT 87.615 149.155 87.785 150.125 ;
        RECT 88.460 149.955 88.630 150.625 ;
        RECT 85.755 148.985 87.785 149.155 ;
        RECT 88.295 148.985 88.630 149.955 ;
        RECT 89.270 149.825 89.620 150.475 ;
        RECT 89.790 149.655 90.020 150.645 ;
        RECT 89.355 149.485 90.020 149.655 ;
        RECT 89.355 148.985 89.525 149.485 ;
        RECT 90.195 148.985 90.420 151.105 ;
        RECT 91.135 150.815 91.305 151.145 ;
        RECT 91.605 150.985 92.620 151.185 ;
        RECT 90.610 150.625 91.305 150.815 ;
        RECT 90.610 149.655 90.780 150.625 ;
        RECT 90.950 149.825 91.360 150.445 ;
        RECT 91.530 149.875 91.750 150.745 ;
        RECT 91.930 150.435 92.280 150.805 ;
        RECT 92.450 150.255 92.620 150.985 ;
        RECT 93.490 150.725 93.740 151.155 ;
        RECT 94.820 150.975 95.670 151.145 ;
        RECT 92.790 150.385 93.200 150.715 ;
        RECT 93.490 150.385 93.910 150.725 ;
        RECT 92.200 150.215 92.620 150.255 ;
        RECT 92.200 150.045 93.550 150.215 ;
        RECT 90.610 149.485 91.305 149.655 ;
        RECT 91.530 149.495 92.030 149.875 ;
        RECT 91.135 148.985 91.305 149.485 ;
        RECT 92.200 149.200 92.370 150.045 ;
        RECT 93.300 149.885 93.550 150.045 ;
        RECT 92.540 149.615 92.790 149.875 ;
        RECT 93.720 149.615 93.910 150.385 ;
        RECT 92.540 149.365 93.910 149.615 ;
        RECT 94.080 150.555 95.330 150.725 ;
        RECT 94.080 149.795 94.250 150.555 ;
        RECT 95.000 150.435 95.330 150.555 ;
        RECT 94.420 149.975 94.600 150.385 ;
        RECT 95.500 150.215 95.670 150.975 ;
        RECT 96.710 150.770 97.030 151.100 ;
        RECT 95.860 150.445 96.520 150.715 ;
        RECT 95.860 150.385 96.190 150.445 ;
        RECT 96.340 150.215 96.670 150.275 ;
        RECT 94.770 150.045 96.670 150.215 ;
        RECT 94.080 149.485 94.600 149.795 ;
        RECT 94.770 149.535 94.940 150.045 ;
        RECT 96.840 149.875 97.030 150.770 ;
        RECT 95.110 149.705 97.030 149.875 ;
        RECT 96.710 149.685 97.030 149.705 ;
        RECT 97.230 150.455 97.480 151.105 ;
        RECT 98.125 151.025 98.380 151.185 ;
        RECT 98.125 150.855 98.465 151.025 ;
        RECT 98.125 150.655 98.380 150.855 ;
        RECT 97.230 150.125 98.030 150.455 ;
        RECT 94.770 149.365 95.980 149.535 ;
        RECT 91.540 149.030 92.370 149.200 ;
        RECT 93.170 149.075 93.340 149.365 ;
        RECT 94.770 149.285 94.940 149.365 ;
        RECT 94.310 149.035 94.940 149.285 ;
        RECT 95.740 149.075 95.980 149.365 ;
        RECT 96.710 149.075 96.880 149.685 ;
        RECT 97.230 149.535 97.480 150.125 ;
        RECT 98.200 149.795 98.380 150.655 ;
        RECT 97.150 149.025 97.480 149.535 ;
        RECT 98.125 149.125 98.380 149.795 ;
        RECT 104.445 150.690 104.715 151.035 ;
        RECT 105.455 150.795 105.625 151.145 ;
        RECT 106.325 150.795 106.495 151.145 ;
        RECT 104.445 149.955 104.615 150.690 ;
        RECT 104.885 150.625 106.495 150.795 ;
        RECT 104.885 150.455 105.055 150.625 ;
        RECT 104.785 150.125 105.055 150.455 ;
        RECT 105.225 150.125 105.630 150.455 ;
        RECT 104.885 149.955 105.055 150.125 ;
        RECT 105.800 150.005 106.510 150.455 ;
        RECT 106.680 150.125 107.030 150.695 ;
        RECT 107.205 150.565 107.545 151.195 ;
        RECT 108.155 150.715 108.485 151.195 ;
        RECT 109.050 150.715 109.380 151.195 ;
        RECT 107.205 150.515 107.435 150.565 ;
        RECT 108.155 150.545 109.380 150.715 ;
        RECT 110.010 150.585 110.510 151.195 ;
        RECT 111.000 150.735 111.285 151.195 ;
        RECT 104.445 148.985 104.715 149.955 ;
        RECT 104.885 149.785 105.610 149.955 ;
        RECT 105.800 149.835 106.515 150.005 ;
        RECT 107.205 149.955 107.380 150.515 ;
        RECT 107.550 150.205 108.245 150.375 ;
        RECT 108.075 149.955 108.245 150.205 ;
        RECT 108.420 150.175 108.840 150.375 ;
        RECT 109.010 150.175 109.340 150.375 ;
        RECT 109.510 150.175 109.840 150.375 ;
        RECT 110.010 149.955 110.180 150.585 ;
        RECT 111.000 150.565 111.955 150.735 ;
        RECT 110.365 150.125 110.715 150.375 ;
        RECT 105.440 149.665 105.610 149.785 ;
        RECT 106.710 149.665 107.030 149.955 ;
        RECT 105.440 149.495 107.030 149.665 ;
        RECT 105.375 149.035 107.030 149.325 ;
        RECT 107.205 148.985 107.545 149.955 ;
        RECT 108.075 149.785 110.510 149.955 ;
        RECT 110.885 149.835 111.575 150.395 ;
        RECT 109.050 148.985 109.380 149.785 ;
        RECT 110.180 148.985 110.510 149.785 ;
        RECT 111.745 149.665 111.955 150.565 ;
        RECT 111.000 149.445 111.955 149.665 ;
        RECT 112.125 150.395 112.525 151.195 ;
        RECT 112.715 150.735 112.995 151.195 ;
        RECT 112.715 150.565 113.840 150.735 ;
        RECT 114.010 150.625 114.395 151.195 ;
        RECT 113.390 150.455 113.840 150.565 ;
        RECT 112.125 149.835 113.220 150.395 ;
        RECT 113.390 150.125 113.945 150.455 ;
        RECT 111.000 148.985 111.285 149.445 ;
        RECT 112.125 148.985 112.525 149.835 ;
        RECT 113.390 149.665 113.840 150.125 ;
        RECT 114.115 149.955 114.395 150.625 ;
        RECT 112.715 149.445 113.840 149.665 ;
        RECT 112.715 148.985 112.995 149.445 ;
        RECT 114.010 148.985 114.395 149.955 ;
        RECT 115.950 150.655 116.205 151.185 ;
        RECT 116.925 150.985 117.995 151.155 ;
        RECT 115.950 150.005 116.160 150.655 ;
        RECT 116.925 150.630 117.245 150.985 ;
        RECT 116.920 150.455 117.245 150.630 ;
        RECT 116.330 150.155 117.245 150.455 ;
        RECT 117.415 150.415 117.655 150.815 ;
        RECT 117.825 150.755 117.995 150.985 ;
        RECT 118.525 150.915 119.475 151.195 ;
        RECT 119.695 151.005 120.045 151.175 ;
        RECT 117.825 150.585 118.355 150.755 ;
        RECT 116.330 150.125 117.070 150.155 ;
        RECT 115.950 149.125 116.205 150.005 ;
        RECT 116.900 149.535 117.070 150.125 ;
        RECT 117.415 150.045 117.955 150.415 ;
        RECT 118.135 150.305 118.355 150.585 ;
        RECT 118.525 150.135 118.695 150.915 ;
        RECT 118.290 149.965 118.695 150.135 ;
        RECT 118.865 150.125 119.215 150.745 ;
        RECT 118.290 149.875 118.460 149.965 ;
        RECT 119.385 149.955 119.595 150.745 ;
        RECT 117.240 149.705 118.460 149.875 ;
        RECT 118.920 149.795 119.595 149.955 ;
        RECT 116.900 149.365 117.700 149.535 ;
        RECT 117.530 149.075 117.700 149.365 ;
        RECT 118.290 149.325 118.460 149.705 ;
        RECT 118.630 149.785 119.595 149.795 ;
        RECT 119.785 150.615 120.045 151.005 ;
        RECT 121.460 150.975 122.315 151.145 ;
        RECT 122.520 150.975 123.015 151.145 ;
        RECT 119.785 149.925 119.955 150.615 ;
        RECT 120.125 150.265 120.295 150.445 ;
        RECT 120.465 150.435 121.255 150.685 ;
        RECT 121.460 150.265 121.630 150.975 ;
        RECT 121.800 150.465 122.155 150.685 ;
        RECT 120.125 150.095 121.815 150.265 ;
        RECT 118.630 149.495 119.090 149.785 ;
        RECT 119.785 149.755 121.285 149.925 ;
        RECT 119.785 149.615 119.955 149.755 ;
        RECT 119.395 149.445 119.955 149.615 ;
        RECT 118.290 148.985 119.160 149.325 ;
        RECT 119.395 148.985 119.565 149.445 ;
        RECT 120.400 149.415 121.475 149.585 ;
        RECT 120.400 149.075 120.570 149.415 ;
        RECT 121.305 149.075 121.475 149.415 ;
        RECT 121.645 149.315 121.815 150.095 ;
        RECT 121.985 149.875 122.155 150.465 ;
        RECT 122.325 150.065 122.675 150.685 ;
        RECT 121.985 149.485 122.450 149.875 ;
        RECT 122.845 149.615 123.015 150.975 ;
        RECT 123.185 149.785 123.645 150.835 ;
        RECT 122.620 149.445 123.015 149.615 ;
        RECT 122.620 149.315 122.790 149.445 ;
        RECT 121.645 148.985 122.325 149.315 ;
        RECT 122.540 148.985 122.790 149.315 ;
        RECT 123.380 149.000 123.705 149.785 ;
        RECT 123.875 148.985 124.045 151.105 ;
        RECT 124.715 150.815 124.970 151.105 ;
        RECT 124.220 150.645 124.970 150.815 ;
        RECT 124.220 149.655 124.450 150.645 ;
        RECT 124.620 149.825 124.970 150.475 ;
        RECT 124.220 149.485 124.970 149.655 ;
        RECT 124.715 148.985 124.970 149.485 ;
        RECT 21.355 148.305 23.385 148.475 ;
        RECT 20.265 147.885 20.780 148.295 ;
        RECT 20.265 147.075 20.605 147.885 ;
        RECT 21.355 147.640 21.525 148.305 ;
        RECT 21.920 147.965 23.045 148.135 ;
        RECT 20.775 147.450 21.525 147.640 ;
        RECT 21.695 147.625 22.705 147.795 ;
        RECT 20.265 146.905 21.495 147.075 ;
        RECT 20.540 146.300 20.785 146.905 ;
        RECT 21.695 146.265 21.885 147.625 ;
        RECT 22.055 146.605 22.330 147.425 ;
        RECT 22.535 146.825 22.705 147.625 ;
        RECT 22.875 146.835 23.045 147.965 ;
        RECT 23.215 147.335 23.385 148.305 ;
        RECT 23.895 147.505 24.230 148.475 ;
        RECT 23.215 147.005 23.410 147.335 ;
        RECT 23.635 147.005 23.890 147.335 ;
        RECT 23.635 146.835 23.805 147.005 ;
        RECT 24.060 146.835 24.230 147.505 ;
        RECT 25.765 147.495 26.095 148.475 ;
        RECT 25.345 147.085 25.675 147.335 ;
        RECT 25.845 146.895 26.095 147.495 ;
        RECT 22.875 146.665 23.805 146.835 ;
        RECT 22.875 146.630 23.050 146.665 ;
        RECT 22.055 146.435 22.335 146.605 ;
        RECT 22.055 146.265 22.330 146.435 ;
        RECT 22.520 146.265 23.050 146.630 ;
        RECT 23.975 146.265 24.230 146.835 ;
        RECT 25.765 146.265 26.095 146.895 ;
        RECT 26.705 147.570 26.975 148.475 ;
        RECT 27.655 147.715 27.825 148.475 ;
        RECT 26.705 146.770 26.875 147.570 ;
        RECT 27.160 147.545 27.825 147.715 ;
        RECT 28.175 147.715 28.345 148.475 ;
        RECT 28.175 147.545 28.840 147.715 ;
        RECT 29.025 147.570 29.295 148.475 ;
        RECT 27.160 147.400 27.330 147.545 ;
        RECT 27.045 147.070 27.330 147.400 ;
        RECT 28.670 147.400 28.840 147.545 ;
        RECT 27.160 146.815 27.330 147.070 ;
        RECT 27.565 146.995 27.895 147.365 ;
        RECT 28.105 146.995 28.435 147.365 ;
        RECT 28.670 147.070 28.955 147.400 ;
        RECT 28.670 146.815 28.840 147.070 ;
        RECT 26.705 146.265 26.965 146.770 ;
        RECT 27.160 146.645 27.825 146.815 ;
        RECT 27.655 146.265 27.825 146.645 ;
        RECT 28.175 146.645 28.840 146.815 ;
        RECT 29.125 146.770 29.295 147.570 ;
        RECT 28.175 146.265 28.345 146.645 ;
        RECT 29.035 146.265 29.295 146.770 ;
        RECT 29.470 147.505 29.805 148.475 ;
        RECT 30.315 148.305 32.345 148.475 ;
        RECT 29.470 146.835 29.640 147.505 ;
        RECT 30.315 147.335 30.485 148.305 ;
        RECT 29.810 147.005 30.065 147.335 ;
        RECT 30.290 147.005 30.485 147.335 ;
        RECT 30.655 147.965 31.780 148.135 ;
        RECT 29.895 146.835 30.065 147.005 ;
        RECT 30.655 146.835 30.825 147.965 ;
        RECT 29.470 146.265 29.725 146.835 ;
        RECT 29.895 146.665 30.825 146.835 ;
        RECT 30.995 147.625 32.005 147.795 ;
        RECT 30.995 146.825 31.165 147.625 ;
        RECT 30.650 146.630 30.825 146.665 ;
        RECT 30.650 146.265 31.180 146.630 ;
        RECT 31.370 146.605 31.645 147.425 ;
        RECT 31.365 146.435 31.645 146.605 ;
        RECT 31.370 146.265 31.645 146.435 ;
        RECT 31.815 146.265 32.005 147.625 ;
        RECT 32.175 147.640 32.345 148.305 ;
        RECT 32.920 147.885 33.435 148.295 ;
        RECT 32.175 147.450 32.925 147.640 ;
        RECT 33.095 147.075 33.435 147.885 ;
        RECT 36.110 147.675 36.440 148.475 ;
        RECT 37.240 147.675 37.570 148.475 ;
        RECT 36.110 147.505 38.545 147.675 ;
        RECT 39.075 147.505 39.415 148.475 ;
        RECT 35.905 147.085 36.255 147.335 ;
        RECT 32.205 146.905 33.435 147.075 ;
        RECT 32.915 146.300 33.160 146.905 ;
        RECT 36.440 146.875 36.610 147.505 ;
        RECT 36.780 147.085 37.110 147.285 ;
        RECT 37.280 147.085 37.610 147.285 ;
        RECT 37.780 147.085 38.200 147.285 ;
        RECT 38.375 147.255 38.545 147.505 ;
        RECT 38.375 147.085 39.070 147.255 ;
        RECT 36.110 146.265 36.610 146.875 ;
        RECT 37.240 146.745 38.465 146.915 ;
        RECT 39.240 146.895 39.415 147.505 ;
        RECT 37.240 146.265 37.570 146.745 ;
        RECT 38.135 146.265 38.465 146.745 ;
        RECT 39.075 146.265 39.415 146.895 ;
        RECT 39.585 147.505 39.925 148.475 ;
        RECT 41.430 147.675 41.760 148.475 ;
        RECT 42.560 147.675 42.890 148.475 ;
        RECT 40.455 147.505 42.890 147.675 ;
        RECT 51.550 147.505 51.885 148.475 ;
        RECT 52.395 148.305 54.425 148.475 ;
        RECT 39.585 146.895 39.760 147.505 ;
        RECT 40.455 147.255 40.625 147.505 ;
        RECT 39.930 147.085 40.625 147.255 ;
        RECT 40.800 147.085 41.220 147.285 ;
        RECT 41.390 147.085 41.720 147.285 ;
        RECT 41.890 147.085 42.220 147.285 ;
        RECT 39.585 146.265 39.925 146.895 ;
        RECT 40.535 146.745 41.760 146.915 ;
        RECT 40.535 146.265 40.865 146.745 ;
        RECT 41.430 146.265 41.760 146.745 ;
        RECT 42.390 146.875 42.560 147.505 ;
        RECT 42.745 147.085 43.095 147.335 ;
        RECT 42.390 146.265 42.890 146.875 ;
        RECT 51.550 146.835 51.720 147.505 ;
        RECT 52.395 147.335 52.565 148.305 ;
        RECT 51.890 147.005 52.145 147.335 ;
        RECT 52.370 147.005 52.565 147.335 ;
        RECT 52.735 147.965 53.860 148.135 ;
        RECT 51.975 146.835 52.145 147.005 ;
        RECT 52.735 146.835 52.905 147.965 ;
        RECT 51.550 146.265 51.805 146.835 ;
        RECT 51.975 146.665 52.905 146.835 ;
        RECT 53.075 147.625 54.085 147.795 ;
        RECT 53.075 146.825 53.245 147.625 ;
        RECT 53.450 147.285 53.725 147.425 ;
        RECT 53.445 147.115 53.725 147.285 ;
        RECT 52.730 146.630 52.905 146.665 ;
        RECT 52.730 146.265 53.260 146.630 ;
        RECT 53.450 146.265 53.725 147.115 ;
        RECT 53.895 146.265 54.085 147.625 ;
        RECT 54.255 147.640 54.425 148.305 ;
        RECT 55.000 147.885 55.515 148.295 ;
        RECT 54.255 147.450 55.005 147.640 ;
        RECT 55.175 147.075 55.515 147.885 ;
        RECT 54.285 146.905 55.515 147.075 ;
        RECT 55.685 147.505 56.025 148.475 ;
        RECT 57.530 147.675 57.860 148.475 ;
        RECT 58.660 147.675 58.990 148.475 ;
        RECT 60.915 148.305 62.945 148.475 ;
        RECT 56.555 147.505 58.990 147.675 ;
        RECT 59.825 147.885 60.340 148.295 ;
        RECT 54.995 146.300 55.240 146.905 ;
        RECT 55.685 146.895 55.860 147.505 ;
        RECT 56.555 147.255 56.725 147.505 ;
        RECT 56.030 147.085 56.725 147.255 ;
        RECT 56.900 147.085 57.320 147.285 ;
        RECT 57.490 147.085 57.820 147.285 ;
        RECT 57.990 147.085 58.320 147.285 ;
        RECT 55.685 146.265 56.025 146.895 ;
        RECT 56.635 146.745 57.860 146.915 ;
        RECT 56.635 146.265 56.965 146.745 ;
        RECT 57.530 146.265 57.860 146.745 ;
        RECT 58.490 146.875 58.660 147.505 ;
        RECT 58.845 147.085 59.195 147.335 ;
        RECT 59.825 147.075 60.165 147.885 ;
        RECT 60.915 147.640 61.085 148.305 ;
        RECT 61.480 147.965 62.605 148.135 ;
        RECT 60.335 147.450 61.085 147.640 ;
        RECT 61.255 147.625 62.265 147.795 ;
        RECT 59.825 146.905 61.055 147.075 ;
        RECT 58.490 146.265 58.990 146.875 ;
        RECT 60.100 146.300 60.345 146.905 ;
        RECT 61.255 146.265 61.445 147.625 ;
        RECT 61.615 146.945 61.890 147.425 ;
        RECT 61.615 146.775 61.895 146.945 ;
        RECT 62.095 146.825 62.265 147.625 ;
        RECT 62.435 146.835 62.605 147.965 ;
        RECT 62.775 147.335 62.945 148.305 ;
        RECT 63.455 147.505 63.790 148.475 ;
        RECT 62.775 147.005 62.970 147.335 ;
        RECT 63.195 147.005 63.450 147.335 ;
        RECT 63.195 146.835 63.365 147.005 ;
        RECT 63.620 146.835 63.790 147.505 ;
        RECT 61.615 146.265 61.890 146.775 ;
        RECT 62.435 146.665 63.365 146.835 ;
        RECT 62.435 146.630 62.610 146.665 ;
        RECT 62.080 146.265 62.610 146.630 ;
        RECT 63.535 146.265 63.790 146.835 ;
        RECT 71.305 147.570 71.560 148.475 ;
        RECT 72.275 147.715 72.445 148.475 ;
        RECT 71.305 146.840 71.475 147.570 ;
        RECT 71.730 147.545 72.445 147.715 ;
        RECT 72.795 147.715 72.965 148.475 ;
        RECT 72.795 147.545 73.510 147.715 ;
        RECT 73.680 147.570 73.935 148.475 ;
        RECT 71.730 147.335 71.900 147.545 ;
        RECT 71.645 147.005 71.900 147.335 ;
        RECT 71.305 146.265 71.560 146.840 ;
        RECT 71.730 146.815 71.900 147.005 ;
        RECT 72.180 146.995 72.535 147.365 ;
        RECT 72.705 146.995 73.060 147.365 ;
        RECT 73.340 147.335 73.510 147.545 ;
        RECT 73.340 147.005 73.595 147.335 ;
        RECT 73.340 146.815 73.510 147.005 ;
        RECT 73.765 146.840 73.935 147.570 ;
        RECT 76.590 147.675 76.920 148.475 ;
        RECT 77.720 147.675 78.050 148.475 ;
        RECT 76.590 147.505 79.025 147.675 ;
        RECT 79.555 147.505 79.895 148.475 ;
        RECT 76.385 147.085 76.735 147.335 ;
        RECT 76.920 146.875 77.090 147.505 ;
        RECT 77.260 147.085 77.590 147.285 ;
        RECT 77.760 147.085 78.090 147.285 ;
        RECT 78.260 147.085 78.680 147.285 ;
        RECT 78.855 147.255 79.025 147.505 ;
        RECT 78.855 147.085 79.550 147.255 ;
        RECT 71.730 146.645 72.445 146.815 ;
        RECT 72.275 146.265 72.445 146.645 ;
        RECT 72.795 146.645 73.510 146.815 ;
        RECT 72.795 146.265 72.965 146.645 ;
        RECT 73.680 146.265 73.935 146.840 ;
        RECT 76.590 146.265 77.090 146.875 ;
        RECT 77.720 146.745 78.945 146.915 ;
        RECT 79.720 146.895 79.895 147.505 ;
        RECT 77.720 146.265 78.050 146.745 ;
        RECT 78.615 146.265 78.945 146.745 ;
        RECT 79.555 146.265 79.895 146.895 ;
        RECT 80.065 147.505 80.405 148.475 ;
        RECT 81.910 147.675 82.240 148.475 ;
        RECT 83.040 147.675 83.370 148.475 ;
        RECT 80.935 147.505 83.370 147.675 ;
        RECT 80.065 146.895 80.240 147.505 ;
        RECT 80.935 147.255 81.105 147.505 ;
        RECT 80.410 147.085 81.105 147.255 ;
        RECT 81.280 147.085 81.700 147.285 ;
        RECT 81.870 147.085 82.200 147.285 ;
        RECT 82.370 147.085 82.700 147.285 ;
        RECT 80.065 146.265 80.405 146.895 ;
        RECT 81.015 146.745 82.240 146.915 ;
        RECT 81.015 146.265 81.345 146.745 ;
        RECT 81.910 146.265 82.240 146.745 ;
        RECT 82.870 146.875 83.040 147.505 ;
        RECT 84.185 147.495 84.515 148.475 ;
        RECT 85.500 147.665 85.755 148.335 ;
        RECT 86.400 147.925 86.730 148.435 ;
        RECT 83.225 147.085 83.575 147.335 ;
        RECT 84.185 146.895 84.435 147.495 ;
        RECT 84.605 147.085 84.935 147.335 ;
        RECT 82.870 146.265 83.370 146.875 ;
        RECT 84.185 146.265 84.515 146.895 ;
        RECT 85.500 146.805 85.680 147.665 ;
        RECT 86.400 147.335 86.650 147.925 ;
        RECT 87.000 147.775 87.170 148.385 ;
        RECT 87.900 148.095 88.140 148.385 ;
        RECT 88.940 148.175 89.570 148.425 ;
        RECT 88.940 148.095 89.110 148.175 ;
        RECT 90.540 148.095 90.710 148.385 ;
        RECT 91.510 148.260 92.340 148.430 ;
        RECT 87.900 147.925 89.110 148.095 ;
        RECT 85.850 147.005 86.650 147.335 ;
        RECT 85.500 146.605 85.755 146.805 ;
        RECT 85.415 146.435 85.755 146.605 ;
        RECT 85.500 146.275 85.755 146.435 ;
        RECT 86.400 146.355 86.650 147.005 ;
        RECT 86.850 147.755 87.170 147.775 ;
        RECT 86.850 147.585 88.770 147.755 ;
        RECT 86.850 146.690 87.040 147.585 ;
        RECT 88.940 147.415 89.110 147.925 ;
        RECT 89.280 147.665 89.800 147.975 ;
        RECT 87.210 147.245 89.110 147.415 ;
        RECT 87.210 147.185 87.540 147.245 ;
        RECT 87.690 147.015 88.020 147.075 ;
        RECT 87.360 146.745 88.020 147.015 ;
        RECT 86.850 146.360 87.170 146.690 ;
        RECT 88.210 146.485 88.380 147.245 ;
        RECT 89.280 147.075 89.460 147.485 ;
        RECT 88.550 146.905 88.880 147.025 ;
        RECT 89.630 146.905 89.800 147.665 ;
        RECT 88.550 146.735 89.800 146.905 ;
        RECT 89.970 147.845 91.340 148.095 ;
        RECT 89.970 147.075 90.160 147.845 ;
        RECT 91.090 147.585 91.340 147.845 ;
        RECT 90.330 147.415 90.580 147.575 ;
        RECT 91.510 147.415 91.680 148.260 ;
        RECT 92.575 147.975 92.745 148.475 ;
        RECT 91.850 147.585 92.350 147.965 ;
        RECT 92.575 147.805 93.270 147.975 ;
        RECT 90.330 147.245 91.680 147.415 ;
        RECT 91.260 147.205 91.680 147.245 ;
        RECT 89.970 146.735 90.390 147.075 ;
        RECT 90.680 146.745 91.090 147.075 ;
        RECT 88.210 146.315 89.060 146.485 ;
        RECT 90.140 146.305 90.390 146.735 ;
        RECT 91.260 146.475 91.430 147.205 ;
        RECT 91.600 146.655 91.950 147.025 ;
        RECT 92.130 146.715 92.350 147.585 ;
        RECT 92.520 147.015 92.930 147.635 ;
        RECT 93.100 146.835 93.270 147.805 ;
        RECT 92.575 146.645 93.270 146.835 ;
        RECT 91.260 146.275 92.275 146.475 ;
        RECT 92.575 146.315 92.745 146.645 ;
        RECT 93.460 146.355 93.685 148.475 ;
        RECT 94.355 147.975 94.525 148.475 ;
        RECT 93.860 147.805 94.525 147.975 ;
        RECT 93.860 146.815 94.090 147.805 ;
        RECT 94.260 146.985 94.610 147.635 ;
        RECT 96.145 147.495 96.475 148.475 ;
        RECT 98.175 148.305 100.205 148.475 ;
        RECT 95.725 147.085 96.055 147.335 ;
        RECT 96.225 146.895 96.475 147.495 ;
        RECT 97.085 147.885 97.600 148.295 ;
        RECT 97.085 147.075 97.425 147.885 ;
        RECT 98.175 147.640 98.345 148.305 ;
        RECT 98.740 147.965 99.865 148.135 ;
        RECT 97.595 147.450 98.345 147.640 ;
        RECT 98.515 147.625 99.525 147.795 ;
        RECT 97.085 146.905 98.315 147.075 ;
        RECT 93.860 146.645 94.525 146.815 ;
        RECT 94.355 146.355 94.525 146.645 ;
        RECT 96.145 146.265 96.475 146.895 ;
        RECT 97.360 146.300 97.605 146.905 ;
        RECT 98.515 146.265 98.705 147.625 ;
        RECT 98.875 147.285 99.150 147.425 ;
        RECT 98.875 147.115 99.155 147.285 ;
        RECT 98.875 146.265 99.150 147.115 ;
        RECT 99.355 146.825 99.525 147.625 ;
        RECT 99.695 146.835 99.865 147.965 ;
        RECT 100.035 147.335 100.205 148.305 ;
        RECT 100.715 147.505 101.050 148.475 ;
        RECT 102.235 147.715 102.405 148.475 ;
        RECT 102.235 147.545 102.900 147.715 ;
        RECT 103.085 147.570 103.355 148.475 ;
        RECT 100.035 147.005 100.230 147.335 ;
        RECT 100.455 147.005 100.710 147.335 ;
        RECT 100.455 146.835 100.625 147.005 ;
        RECT 100.880 146.835 101.050 147.505 ;
        RECT 102.730 147.400 102.900 147.545 ;
        RECT 102.165 146.995 102.495 147.365 ;
        RECT 102.730 147.070 103.015 147.400 ;
        RECT 99.695 146.665 100.625 146.835 ;
        RECT 99.695 146.630 99.870 146.665 ;
        RECT 99.340 146.265 99.870 146.630 ;
        RECT 100.795 146.265 101.050 146.835 ;
        RECT 102.730 146.815 102.900 147.070 ;
        RECT 102.235 146.645 102.900 146.815 ;
        RECT 103.185 146.770 103.355 147.570 ;
        RECT 102.235 146.265 102.405 146.645 ;
        RECT 103.095 146.265 103.355 146.770 ;
        RECT 103.985 147.505 104.255 148.475 ;
        RECT 104.915 148.135 106.570 148.425 ;
        RECT 104.980 147.795 106.570 147.965 ;
        RECT 104.980 147.675 105.150 147.795 ;
        RECT 104.425 147.505 105.150 147.675 ;
        RECT 103.985 146.770 104.155 147.505 ;
        RECT 104.425 147.335 104.595 147.505 ;
        RECT 105.340 147.455 106.055 147.625 ;
        RECT 106.250 147.505 106.570 147.795 ;
        RECT 106.745 147.505 107.085 148.475 ;
        RECT 108.590 147.675 108.920 148.475 ;
        RECT 109.720 147.675 110.050 148.475 ;
        RECT 113.355 148.305 115.385 148.475 ;
        RECT 107.615 147.505 110.050 147.675 ;
        RECT 112.265 147.885 112.780 148.295 ;
        RECT 104.325 147.005 104.595 147.335 ;
        RECT 104.765 147.005 105.170 147.335 ;
        RECT 105.340 147.005 106.050 147.455 ;
        RECT 104.425 146.835 104.595 147.005 ;
        RECT 103.985 146.425 104.255 146.770 ;
        RECT 104.425 146.665 106.035 146.835 ;
        RECT 106.220 146.765 106.570 147.335 ;
        RECT 106.745 146.945 106.920 147.505 ;
        RECT 107.615 147.255 107.785 147.505 ;
        RECT 107.090 147.085 107.785 147.255 ;
        RECT 107.960 147.085 108.380 147.285 ;
        RECT 108.550 147.085 108.880 147.285 ;
        RECT 109.050 147.085 109.380 147.285 ;
        RECT 106.745 146.895 106.975 146.945 ;
        RECT 104.995 146.315 105.165 146.665 ;
        RECT 105.865 146.315 106.035 146.665 ;
        RECT 106.745 146.265 107.085 146.895 ;
        RECT 107.695 146.745 108.920 146.915 ;
        RECT 107.695 146.265 108.025 146.745 ;
        RECT 108.590 146.265 108.920 146.745 ;
        RECT 109.550 146.875 109.720 147.505 ;
        RECT 109.905 147.085 110.255 147.335 ;
        RECT 112.265 147.075 112.605 147.885 ;
        RECT 113.355 147.640 113.525 148.305 ;
        RECT 113.920 147.965 115.045 148.135 ;
        RECT 112.775 147.450 113.525 147.640 ;
        RECT 113.695 147.625 114.705 147.795 ;
        RECT 112.265 146.905 113.495 147.075 ;
        RECT 109.550 146.265 110.050 146.875 ;
        RECT 112.540 146.300 112.785 146.905 ;
        RECT 113.695 146.265 113.885 147.625 ;
        RECT 114.055 147.285 114.330 147.425 ;
        RECT 114.055 147.115 114.335 147.285 ;
        RECT 114.055 146.265 114.330 147.115 ;
        RECT 114.535 146.825 114.705 147.625 ;
        RECT 114.875 146.835 115.045 147.965 ;
        RECT 115.215 147.335 115.385 148.305 ;
        RECT 115.895 147.505 116.230 148.475 ;
        RECT 115.215 147.005 115.410 147.335 ;
        RECT 115.635 147.005 115.890 147.335 ;
        RECT 115.635 146.835 115.805 147.005 ;
        RECT 116.060 146.835 116.230 147.505 ;
        RECT 116.780 147.665 117.035 148.335 ;
        RECT 117.680 147.925 118.010 148.435 ;
        RECT 116.780 146.945 116.960 147.665 ;
        RECT 117.680 147.335 117.930 147.925 ;
        RECT 118.280 147.775 118.450 148.385 ;
        RECT 119.180 148.095 119.420 148.385 ;
        RECT 120.220 148.175 120.850 148.425 ;
        RECT 120.220 148.095 120.390 148.175 ;
        RECT 121.820 148.095 121.990 148.385 ;
        RECT 122.790 148.260 123.620 148.430 ;
        RECT 119.180 147.925 120.390 148.095 ;
        RECT 117.130 147.005 117.930 147.335 ;
        RECT 114.875 146.665 115.805 146.835 ;
        RECT 114.875 146.630 115.050 146.665 ;
        RECT 114.520 146.265 115.050 146.630 ;
        RECT 115.975 146.265 116.230 146.835 ;
        RECT 116.695 146.805 116.960 146.945 ;
        RECT 116.695 146.775 117.035 146.805 ;
        RECT 116.780 146.275 117.035 146.775 ;
        RECT 117.680 146.355 117.930 147.005 ;
        RECT 118.130 147.755 118.450 147.775 ;
        RECT 118.130 147.585 120.050 147.755 ;
        RECT 118.130 146.690 118.320 147.585 ;
        RECT 120.220 147.415 120.390 147.925 ;
        RECT 120.560 147.665 121.080 147.975 ;
        RECT 118.490 147.245 120.390 147.415 ;
        RECT 118.490 147.185 118.820 147.245 ;
        RECT 118.970 147.015 119.300 147.075 ;
        RECT 118.640 146.745 119.300 147.015 ;
        RECT 118.130 146.360 118.450 146.690 ;
        RECT 119.490 146.485 119.660 147.245 ;
        RECT 120.560 147.075 120.740 147.485 ;
        RECT 119.830 146.905 120.160 147.025 ;
        RECT 120.910 146.905 121.080 147.665 ;
        RECT 119.830 146.735 121.080 146.905 ;
        RECT 121.250 147.845 122.620 148.095 ;
        RECT 121.250 147.075 121.440 147.845 ;
        RECT 122.370 147.585 122.620 147.845 ;
        RECT 121.610 147.415 121.860 147.575 ;
        RECT 122.790 147.415 122.960 148.260 ;
        RECT 123.855 147.975 124.025 148.475 ;
        RECT 123.130 147.585 123.630 147.965 ;
        RECT 123.855 147.805 124.550 147.975 ;
        RECT 121.610 147.245 122.960 147.415 ;
        RECT 122.540 147.205 122.960 147.245 ;
        RECT 121.250 146.735 121.670 147.075 ;
        RECT 121.960 146.745 122.370 147.075 ;
        RECT 119.490 146.315 120.340 146.485 ;
        RECT 121.420 146.305 121.670 146.735 ;
        RECT 122.540 146.475 122.710 147.205 ;
        RECT 122.880 146.655 123.230 147.025 ;
        RECT 123.410 146.715 123.630 147.585 ;
        RECT 123.800 147.015 124.210 147.635 ;
        RECT 124.380 146.835 124.550 147.805 ;
        RECT 123.855 146.645 124.550 146.835 ;
        RECT 122.540 146.275 123.555 146.475 ;
        RECT 123.855 146.315 124.025 146.645 ;
        RECT 124.740 146.355 124.965 148.475 ;
        RECT 125.635 147.975 125.805 148.475 ;
        RECT 125.140 147.805 125.805 147.975 ;
        RECT 125.140 146.815 125.370 147.805 ;
        RECT 125.540 146.985 125.890 147.635 ;
        RECT 125.140 146.645 125.805 146.815 ;
        RECT 125.635 146.355 125.805 146.645 ;
        RECT 20.705 145.125 21.035 145.755 ;
        RECT 22.480 145.585 22.735 145.745 ;
        RECT 22.395 145.415 22.735 145.585 ;
        RECT 22.480 145.215 22.735 145.415 ;
        RECT 20.705 144.525 20.955 145.125 ;
        RECT 21.125 144.685 21.455 144.935 ;
        RECT 20.705 143.545 21.035 144.525 ;
        RECT 22.480 144.355 22.660 145.215 ;
        RECT 23.380 145.015 23.630 145.665 ;
        RECT 22.830 144.685 23.630 145.015 ;
        RECT 22.480 143.685 22.735 144.355 ;
        RECT 23.380 144.095 23.630 144.685 ;
        RECT 23.830 145.330 24.150 145.660 ;
        RECT 25.190 145.535 26.040 145.705 ;
        RECT 23.830 144.435 24.020 145.330 ;
        RECT 24.340 145.005 25.000 145.275 ;
        RECT 24.670 144.945 25.000 145.005 ;
        RECT 24.190 144.775 24.520 144.835 ;
        RECT 25.190 144.775 25.360 145.535 ;
        RECT 27.120 145.285 27.370 145.715 ;
        RECT 25.530 145.115 26.780 145.285 ;
        RECT 25.530 144.995 25.860 145.115 ;
        RECT 24.190 144.605 26.090 144.775 ;
        RECT 23.830 144.265 25.750 144.435 ;
        RECT 23.830 144.245 24.150 144.265 ;
        RECT 23.380 143.585 23.710 144.095 ;
        RECT 23.980 143.635 24.150 144.245 ;
        RECT 25.920 144.095 26.090 144.605 ;
        RECT 26.260 144.535 26.440 144.945 ;
        RECT 26.610 144.355 26.780 145.115 ;
        RECT 24.880 143.925 26.090 144.095 ;
        RECT 26.260 144.045 26.780 144.355 ;
        RECT 26.950 144.945 27.370 145.285 ;
        RECT 28.240 145.545 29.255 145.745 ;
        RECT 27.660 144.945 28.070 145.275 ;
        RECT 26.950 144.175 27.140 144.945 ;
        RECT 28.240 144.815 28.410 145.545 ;
        RECT 29.555 145.375 29.725 145.705 ;
        RECT 28.580 144.995 28.930 145.365 ;
        RECT 28.240 144.775 28.660 144.815 ;
        RECT 27.310 144.605 28.660 144.775 ;
        RECT 27.310 144.445 27.560 144.605 ;
        RECT 28.070 144.175 28.320 144.435 ;
        RECT 26.950 143.925 28.320 144.175 ;
        RECT 24.880 143.635 25.120 143.925 ;
        RECT 25.920 143.845 26.090 143.925 ;
        RECT 25.920 143.595 26.550 143.845 ;
        RECT 27.520 143.635 27.690 143.925 ;
        RECT 28.490 143.760 28.660 144.605 ;
        RECT 29.110 144.435 29.330 145.305 ;
        RECT 29.555 145.185 30.250 145.375 ;
        RECT 28.830 144.055 29.330 144.435 ;
        RECT 29.500 144.385 29.910 145.005 ;
        RECT 30.080 144.215 30.250 145.185 ;
        RECT 29.555 144.045 30.250 144.215 ;
        RECT 28.490 143.590 29.320 143.760 ;
        RECT 29.555 143.545 29.725 144.045 ;
        RECT 30.440 143.545 30.665 145.665 ;
        RECT 31.335 145.375 31.505 145.665 ;
        RECT 30.840 145.205 31.505 145.375 ;
        RECT 30.840 144.215 31.070 145.205 ;
        RECT 41.405 145.125 41.735 145.755 ;
        RECT 42.435 145.375 42.605 145.665 ;
        RECT 42.435 145.205 43.100 145.375 ;
        RECT 31.240 144.385 31.590 145.035 ;
        RECT 40.985 144.685 41.315 144.935 ;
        RECT 41.485 144.525 41.735 145.125 ;
        RECT 30.840 144.045 31.505 144.215 ;
        RECT 31.335 143.545 31.505 144.045 ;
        RECT 41.405 143.545 41.735 144.525 ;
        RECT 42.350 144.385 42.700 145.035 ;
        RECT 42.870 144.215 43.100 145.205 ;
        RECT 42.435 144.045 43.100 144.215 ;
        RECT 42.435 143.545 42.605 144.045 ;
        RECT 43.275 143.545 43.500 145.665 ;
        RECT 44.215 145.375 44.385 145.705 ;
        RECT 44.685 145.545 45.700 145.745 ;
        RECT 43.690 145.185 44.385 145.375 ;
        RECT 43.690 144.215 43.860 145.185 ;
        RECT 44.030 144.385 44.440 145.005 ;
        RECT 44.610 144.435 44.830 145.305 ;
        RECT 45.010 144.995 45.360 145.365 ;
        RECT 45.530 144.815 45.700 145.545 ;
        RECT 46.570 145.285 46.820 145.715 ;
        RECT 47.900 145.535 48.750 145.705 ;
        RECT 45.870 144.945 46.280 145.275 ;
        RECT 46.570 144.945 46.990 145.285 ;
        RECT 45.280 144.775 45.700 144.815 ;
        RECT 45.280 144.605 46.630 144.775 ;
        RECT 43.690 144.045 44.385 144.215 ;
        RECT 44.610 144.055 45.110 144.435 ;
        RECT 44.215 143.545 44.385 144.045 ;
        RECT 45.280 143.760 45.450 144.605 ;
        RECT 46.380 144.445 46.630 144.605 ;
        RECT 45.620 144.175 45.870 144.435 ;
        RECT 46.800 144.175 46.990 144.945 ;
        RECT 45.620 143.925 46.990 144.175 ;
        RECT 47.160 145.115 48.410 145.285 ;
        RECT 47.160 144.355 47.330 145.115 ;
        RECT 48.080 144.995 48.410 145.115 ;
        RECT 47.500 144.535 47.680 144.945 ;
        RECT 48.580 144.775 48.750 145.535 ;
        RECT 49.790 145.330 50.110 145.660 ;
        RECT 48.940 145.005 49.600 145.275 ;
        RECT 48.940 144.945 49.270 145.005 ;
        RECT 49.420 144.775 49.750 144.835 ;
        RECT 47.850 144.605 49.750 144.775 ;
        RECT 47.160 144.045 47.680 144.355 ;
        RECT 47.850 144.095 48.020 144.605 ;
        RECT 49.920 144.435 50.110 145.330 ;
        RECT 48.190 144.265 50.110 144.435 ;
        RECT 49.790 144.245 50.110 144.265 ;
        RECT 50.310 145.015 50.560 145.665 ;
        RECT 51.205 145.215 51.460 145.745 ;
        RECT 50.310 144.685 51.110 145.015 ;
        RECT 47.850 143.925 49.060 144.095 ;
        RECT 44.620 143.590 45.450 143.760 ;
        RECT 46.250 143.635 46.420 143.925 ;
        RECT 47.850 143.845 48.020 143.925 ;
        RECT 47.390 143.595 48.020 143.845 ;
        RECT 48.820 143.635 49.060 143.925 ;
        RECT 49.790 143.635 49.960 144.245 ;
        RECT 50.310 144.095 50.560 144.685 ;
        RECT 51.280 144.355 51.460 145.215 ;
        RECT 50.230 143.585 50.560 144.095 ;
        RECT 51.205 143.885 51.460 144.355 ;
        RECT 52.005 145.250 52.265 145.755 ;
        RECT 52.955 145.375 53.125 145.755 ;
        RECT 52.005 144.450 52.175 145.250 ;
        RECT 52.460 145.205 53.125 145.375 ;
        RECT 52.460 144.950 52.630 145.205 ;
        RECT 58.885 145.125 59.215 145.755 ;
        RECT 52.345 144.620 52.630 144.950 ;
        RECT 52.865 144.655 53.195 145.025 ;
        RECT 58.465 144.685 58.795 144.935 ;
        RECT 52.460 144.475 52.630 144.620 ;
        RECT 58.965 144.525 59.215 145.125 ;
        RECT 64.240 145.115 64.485 145.720 ;
        RECT 51.205 143.715 51.545 143.885 ;
        RECT 51.205 143.685 51.460 143.715 ;
        RECT 52.005 143.545 52.275 144.450 ;
        RECT 52.460 144.305 53.125 144.475 ;
        RECT 52.955 143.545 53.125 144.305 ;
        RECT 58.885 143.545 59.215 144.525 ;
        RECT 63.965 144.945 65.195 145.115 ;
        RECT 63.965 144.135 64.305 144.945 ;
        RECT 64.475 144.380 65.225 144.570 ;
        RECT 63.965 143.725 64.480 144.135 ;
        RECT 65.055 143.715 65.225 144.380 ;
        RECT 65.395 144.395 65.585 145.755 ;
        RECT 65.755 144.905 66.030 145.755 ;
        RECT 66.220 145.390 66.750 145.755 ;
        RECT 66.575 145.355 66.750 145.390 ;
        RECT 65.755 144.735 66.035 144.905 ;
        RECT 65.755 144.595 66.030 144.735 ;
        RECT 66.235 144.395 66.405 145.195 ;
        RECT 65.395 144.225 66.405 144.395 ;
        RECT 66.575 145.185 67.505 145.355 ;
        RECT 67.675 145.185 67.930 145.755 ;
        RECT 80.145 145.355 80.315 145.705 ;
        RECT 81.015 145.355 81.185 145.705 ;
        RECT 66.575 144.055 66.745 145.185 ;
        RECT 67.335 145.015 67.505 145.185 ;
        RECT 65.620 143.885 66.745 144.055 ;
        RECT 66.915 144.685 67.110 145.015 ;
        RECT 67.335 144.685 67.590 145.015 ;
        RECT 66.915 143.715 67.085 144.685 ;
        RECT 67.760 144.515 67.930 145.185 ;
        RECT 79.610 144.685 79.960 145.255 ;
        RECT 80.145 145.185 81.755 145.355 ;
        RECT 81.925 145.250 82.195 145.595 ;
        RECT 81.585 145.015 81.755 145.185 ;
        RECT 80.130 144.565 80.840 145.015 ;
        RECT 81.010 144.685 81.415 145.015 ;
        RECT 81.585 144.685 81.855 145.015 ;
        RECT 65.055 143.545 67.085 143.715 ;
        RECT 67.595 143.545 67.930 144.515 ;
        RECT 79.610 144.225 79.930 144.515 ;
        RECT 80.125 144.395 80.840 144.565 ;
        RECT 81.585 144.515 81.755 144.685 ;
        RECT 82.025 144.515 82.195 145.250 ;
        RECT 84.940 145.115 85.185 145.720 ;
        RECT 81.030 144.345 81.755 144.515 ;
        RECT 81.030 144.225 81.200 144.345 ;
        RECT 79.610 144.055 81.200 144.225 ;
        RECT 79.610 143.595 81.265 143.885 ;
        RECT 81.925 143.545 82.195 144.515 ;
        RECT 84.665 144.945 85.895 145.115 ;
        RECT 84.665 144.135 85.005 144.945 ;
        RECT 85.175 144.380 85.925 144.570 ;
        RECT 84.665 143.725 85.180 144.135 ;
        RECT 85.755 143.715 85.925 144.380 ;
        RECT 86.095 144.395 86.285 145.755 ;
        RECT 86.455 144.905 86.730 145.755 ;
        RECT 86.920 145.390 87.450 145.755 ;
        RECT 87.275 145.355 87.450 145.390 ;
        RECT 86.455 144.735 86.735 144.905 ;
        RECT 86.455 144.595 86.730 144.735 ;
        RECT 86.935 144.395 87.105 145.195 ;
        RECT 86.095 144.225 87.105 144.395 ;
        RECT 87.275 145.185 88.205 145.355 ;
        RECT 88.375 145.185 88.630 145.755 ;
        RECT 90.275 145.375 90.445 145.755 ;
        RECT 90.275 145.205 90.940 145.375 ;
        RECT 91.135 145.250 91.395 145.755 ;
        RECT 87.275 144.055 87.445 145.185 ;
        RECT 88.035 145.015 88.205 145.185 ;
        RECT 86.320 143.885 87.445 144.055 ;
        RECT 87.615 144.685 87.810 145.015 ;
        RECT 88.035 144.685 88.290 145.015 ;
        RECT 87.615 143.715 87.785 144.685 ;
        RECT 88.460 144.515 88.630 145.185 ;
        RECT 90.205 144.655 90.535 145.025 ;
        RECT 90.770 144.950 90.940 145.205 ;
        RECT 85.755 143.545 87.785 143.715 ;
        RECT 88.295 143.545 88.630 144.515 ;
        RECT 90.770 144.620 91.055 144.950 ;
        RECT 90.770 144.475 90.940 144.620 ;
        RECT 90.275 144.305 90.940 144.475 ;
        RECT 91.225 144.450 91.395 145.250 ;
        RECT 90.275 143.545 90.445 144.305 ;
        RECT 91.125 143.545 91.395 144.450 ;
        RECT 91.565 145.250 91.825 145.755 ;
        RECT 92.515 145.375 92.685 145.755 ;
        RECT 91.565 144.450 91.735 145.250 ;
        RECT 92.020 145.205 92.685 145.375 ;
        RECT 93.060 145.295 93.345 145.755 ;
        RECT 92.020 144.950 92.190 145.205 ;
        RECT 93.060 145.125 94.015 145.295 ;
        RECT 91.905 144.620 92.190 144.950 ;
        RECT 92.425 144.655 92.755 145.025 ;
        RECT 92.020 144.475 92.190 144.620 ;
        RECT 91.565 143.545 91.835 144.450 ;
        RECT 92.020 144.305 92.685 144.475 ;
        RECT 92.945 144.395 93.635 144.955 ;
        RECT 92.515 143.545 92.685 144.305 ;
        RECT 93.805 144.225 94.015 145.125 ;
        RECT 93.060 144.005 94.015 144.225 ;
        RECT 94.185 144.955 94.585 145.755 ;
        RECT 94.775 145.295 95.055 145.755 ;
        RECT 94.775 145.125 95.900 145.295 ;
        RECT 96.070 145.185 96.455 145.755 ;
        RECT 95.450 145.015 95.900 145.125 ;
        RECT 94.185 144.395 95.280 144.955 ;
        RECT 95.450 144.685 96.005 145.015 ;
        RECT 93.060 143.545 93.345 144.005 ;
        RECT 94.185 143.545 94.585 144.395 ;
        RECT 95.450 144.225 95.900 144.685 ;
        RECT 96.175 144.515 96.455 145.185 ;
        RECT 94.775 144.005 95.900 144.225 ;
        RECT 94.775 143.545 95.055 144.005 ;
        RECT 96.070 143.545 96.455 144.515 ;
        RECT 96.630 145.215 96.885 145.745 ;
        RECT 97.605 145.545 98.675 145.715 ;
        RECT 96.630 144.565 96.840 145.215 ;
        RECT 97.605 145.190 97.925 145.545 ;
        RECT 97.600 145.015 97.925 145.190 ;
        RECT 97.010 144.715 97.925 145.015 ;
        RECT 98.095 144.975 98.335 145.375 ;
        RECT 98.505 145.315 98.675 145.545 ;
        RECT 99.205 145.475 100.155 145.755 ;
        RECT 100.375 145.565 100.725 145.735 ;
        RECT 98.505 145.145 99.035 145.315 ;
        RECT 97.010 144.685 97.750 144.715 ;
        RECT 96.630 143.685 96.885 144.565 ;
        RECT 97.580 144.095 97.750 144.685 ;
        RECT 98.095 144.605 98.635 144.975 ;
        RECT 98.815 144.865 99.035 145.145 ;
        RECT 99.205 144.695 99.375 145.475 ;
        RECT 98.970 144.525 99.375 144.695 ;
        RECT 99.545 144.685 99.895 145.305 ;
        RECT 98.970 144.435 99.140 144.525 ;
        RECT 100.065 144.515 100.275 145.305 ;
        RECT 97.920 144.265 99.140 144.435 ;
        RECT 99.600 144.355 100.275 144.515 ;
        RECT 97.580 143.925 98.380 144.095 ;
        RECT 98.210 143.635 98.380 143.925 ;
        RECT 98.970 143.885 99.140 144.265 ;
        RECT 99.310 144.345 100.275 144.355 ;
        RECT 100.465 145.175 100.725 145.565 ;
        RECT 102.140 145.535 102.995 145.705 ;
        RECT 103.200 145.535 103.695 145.705 ;
        RECT 100.465 144.485 100.635 145.175 ;
        RECT 100.805 144.825 100.975 145.005 ;
        RECT 101.145 144.995 101.935 145.245 ;
        RECT 102.140 144.825 102.310 145.535 ;
        RECT 102.480 145.025 102.835 145.245 ;
        RECT 100.805 144.655 102.495 144.825 ;
        RECT 99.310 144.055 99.770 144.345 ;
        RECT 100.465 144.315 101.965 144.485 ;
        RECT 100.465 144.175 100.635 144.315 ;
        RECT 100.075 144.005 100.635 144.175 ;
        RECT 98.970 143.545 99.840 143.885 ;
        RECT 100.075 143.545 100.245 144.005 ;
        RECT 101.080 143.975 102.155 144.145 ;
        RECT 101.080 143.635 101.250 143.975 ;
        RECT 101.985 143.635 102.155 143.975 ;
        RECT 102.325 143.875 102.495 144.655 ;
        RECT 102.665 144.435 102.835 145.025 ;
        RECT 103.005 144.625 103.355 145.245 ;
        RECT 102.665 144.045 103.130 144.435 ;
        RECT 103.525 144.175 103.695 145.535 ;
        RECT 103.865 144.345 104.325 145.395 ;
        RECT 103.300 144.005 103.695 144.175 ;
        RECT 103.300 143.875 103.470 144.005 ;
        RECT 102.325 143.545 103.005 143.875 ;
        RECT 103.220 143.545 103.470 143.875 ;
        RECT 104.060 143.560 104.385 144.345 ;
        RECT 104.555 143.545 104.725 145.665 ;
        RECT 105.395 145.375 105.650 145.665 ;
        RECT 104.900 145.205 105.650 145.375 ;
        RECT 104.900 144.215 105.130 145.205 ;
        RECT 110.170 145.145 110.670 145.755 ;
        RECT 105.300 144.385 105.650 145.035 ;
        RECT 109.965 144.685 110.315 144.935 ;
        RECT 110.500 144.515 110.670 145.145 ;
        RECT 111.300 145.275 111.630 145.755 ;
        RECT 112.195 145.275 112.525 145.755 ;
        RECT 111.300 145.105 112.525 145.275 ;
        RECT 113.135 145.125 113.475 145.755 ;
        RECT 110.840 144.735 111.170 144.935 ;
        RECT 111.340 144.735 111.670 144.935 ;
        RECT 111.840 144.735 112.260 144.935 ;
        RECT 112.435 144.765 113.130 144.935 ;
        RECT 112.435 144.515 112.605 144.765 ;
        RECT 113.300 144.515 113.475 145.125 ;
        RECT 115.760 145.115 116.005 145.720 ;
        RECT 110.170 144.345 112.605 144.515 ;
        RECT 104.900 144.045 105.650 144.215 ;
        RECT 105.395 143.545 105.650 144.045 ;
        RECT 110.170 143.545 110.500 144.345 ;
        RECT 111.300 143.545 111.630 144.345 ;
        RECT 113.135 143.545 113.475 144.515 ;
        RECT 115.485 144.945 116.715 145.115 ;
        RECT 115.485 144.135 115.825 144.945 ;
        RECT 115.995 144.380 116.745 144.570 ;
        RECT 115.485 143.725 116.000 144.135 ;
        RECT 116.575 143.715 116.745 144.380 ;
        RECT 116.915 144.395 117.105 145.755 ;
        RECT 117.275 145.585 117.550 145.755 ;
        RECT 117.275 145.415 117.555 145.585 ;
        RECT 117.275 144.595 117.550 145.415 ;
        RECT 117.740 145.390 118.270 145.755 ;
        RECT 118.095 145.355 118.270 145.390 ;
        RECT 117.755 144.395 117.925 145.195 ;
        RECT 116.915 144.225 117.925 144.395 ;
        RECT 118.095 145.185 119.025 145.355 ;
        RECT 119.195 145.185 119.450 145.755 ;
        RECT 118.095 144.055 118.265 145.185 ;
        RECT 118.855 145.015 119.025 145.185 ;
        RECT 117.140 143.885 118.265 144.055 ;
        RECT 118.435 144.685 118.630 145.015 ;
        RECT 118.855 144.685 119.110 145.015 ;
        RECT 118.435 143.715 118.605 144.685 ;
        RECT 119.280 144.515 119.450 145.185 ;
        RECT 120.065 145.125 120.395 145.755 ;
        RECT 121.555 145.375 121.725 145.755 ;
        RECT 121.555 145.205 122.220 145.375 ;
        RECT 122.415 145.250 122.675 145.755 ;
        RECT 119.645 144.685 119.975 144.935 ;
        RECT 120.145 144.525 120.395 145.125 ;
        RECT 121.485 144.655 121.815 145.025 ;
        RECT 122.050 144.950 122.220 145.205 ;
        RECT 116.575 143.545 118.605 143.715 ;
        RECT 119.115 143.545 119.450 144.515 ;
        RECT 120.065 143.545 120.395 144.525 ;
        RECT 122.050 144.620 122.335 144.950 ;
        RECT 122.050 144.475 122.220 144.620 ;
        RECT 121.555 144.305 122.220 144.475 ;
        RECT 122.505 144.450 122.675 145.250 ;
        RECT 121.555 143.545 121.725 144.305 ;
        RECT 122.405 143.545 122.675 144.450 ;
        RECT 34.525 142.065 34.795 143.035 ;
        RECT 35.455 142.695 37.110 142.985 ;
        RECT 47.410 142.695 49.065 142.985 ;
        RECT 35.520 142.355 37.110 142.525 ;
        RECT 35.520 142.235 35.690 142.355 ;
        RECT 34.965 142.065 35.690 142.235 ;
        RECT 34.525 141.330 34.695 142.065 ;
        RECT 34.965 141.895 35.135 142.065 ;
        RECT 34.865 141.565 35.135 141.895 ;
        RECT 35.305 141.565 35.710 141.895 ;
        RECT 35.880 141.565 36.590 142.185 ;
        RECT 36.790 142.065 37.110 142.355 ;
        RECT 47.410 142.355 49.000 142.525 ;
        RECT 47.410 142.065 47.730 142.355 ;
        RECT 48.830 142.235 49.000 142.355 ;
        RECT 47.925 142.015 48.640 142.185 ;
        RECT 48.830 142.065 49.555 142.235 ;
        RECT 49.725 142.065 49.995 143.035 ;
        RECT 34.965 141.395 35.135 141.565 ;
        RECT 34.525 140.985 34.795 141.330 ;
        RECT 34.965 141.225 36.575 141.395 ;
        RECT 36.760 141.325 37.110 141.895 ;
        RECT 47.410 141.325 47.760 141.895 ;
        RECT 47.930 141.565 48.640 142.015 ;
        RECT 49.385 141.895 49.555 142.065 ;
        RECT 48.810 141.565 49.215 141.895 ;
        RECT 49.385 141.565 49.655 141.895 ;
        RECT 49.385 141.395 49.555 141.565 ;
        RECT 35.535 140.875 35.705 141.225 ;
        RECT 36.405 140.875 36.575 141.225 ;
        RECT 47.945 141.225 49.555 141.395 ;
        RECT 49.825 141.330 49.995 142.065 ;
        RECT 47.945 140.875 48.115 141.225 ;
        RECT 48.815 140.875 48.985 141.225 ;
        RECT 49.725 140.985 49.995 141.330 ;
        RECT 52.465 142.065 52.805 143.035 ;
        RECT 54.310 142.235 54.640 143.035 ;
        RECT 55.440 142.235 55.770 143.035 ;
        RECT 56.260 142.575 56.545 143.035 ;
        RECT 56.260 142.355 57.215 142.575 ;
        RECT 53.335 142.065 55.770 142.235 ;
        RECT 52.465 141.505 52.640 142.065 ;
        RECT 53.335 141.815 53.505 142.065 ;
        RECT 52.810 141.645 53.505 141.815 ;
        RECT 53.675 141.675 54.100 141.845 ;
        RECT 53.680 141.645 54.100 141.675 ;
        RECT 54.270 141.645 54.600 141.845 ;
        RECT 54.770 141.645 55.100 141.845 ;
        RECT 52.465 141.455 52.695 141.505 ;
        RECT 52.465 140.825 52.805 141.455 ;
        RECT 53.415 141.305 54.640 141.475 ;
        RECT 53.415 140.825 53.745 141.305 ;
        RECT 54.310 140.825 54.640 141.305 ;
        RECT 55.270 141.435 55.440 142.065 ;
        RECT 55.625 141.645 55.975 141.895 ;
        RECT 56.145 141.625 56.835 142.185 ;
        RECT 57.005 141.455 57.215 142.355 ;
        RECT 55.270 140.825 55.770 141.435 ;
        RECT 56.260 141.285 57.215 141.455 ;
        RECT 57.385 142.185 57.785 143.035 ;
        RECT 57.975 142.575 58.255 143.035 ;
        RECT 57.975 142.355 59.100 142.575 ;
        RECT 57.385 141.625 58.480 142.185 ;
        RECT 58.650 141.895 59.100 142.355 ;
        RECT 59.270 142.065 59.655 143.035 ;
        RECT 56.260 140.825 56.545 141.285 ;
        RECT 57.385 140.825 57.785 141.625 ;
        RECT 58.650 141.565 59.205 141.895 ;
        RECT 58.650 141.455 59.100 141.565 ;
        RECT 57.975 141.285 59.100 141.455 ;
        RECT 59.375 141.395 59.655 142.065 ;
        RECT 57.975 140.825 58.255 141.285 ;
        RECT 59.270 140.825 59.655 141.395 ;
        RECT 59.830 142.015 60.085 142.895 ;
        RECT 61.410 142.655 61.580 142.945 ;
        RECT 60.780 142.485 61.580 142.655 ;
        RECT 62.170 142.695 63.040 143.035 ;
        RECT 59.830 141.365 60.040 142.015 ;
        RECT 60.780 141.895 60.950 142.485 ;
        RECT 62.170 142.315 62.340 142.695 ;
        RECT 63.275 142.575 63.445 143.035 ;
        RECT 64.280 142.605 64.450 142.945 ;
        RECT 65.185 142.605 65.355 142.945 ;
        RECT 61.120 142.145 62.340 142.315 ;
        RECT 62.510 142.235 62.970 142.525 ;
        RECT 63.275 142.405 63.835 142.575 ;
        RECT 64.280 142.435 65.355 142.605 ;
        RECT 65.525 142.705 66.205 143.035 ;
        RECT 66.420 142.705 66.670 143.035 ;
        RECT 63.665 142.265 63.835 142.405 ;
        RECT 62.510 142.225 63.475 142.235 ;
        RECT 62.170 142.055 62.340 142.145 ;
        RECT 62.800 142.065 63.475 142.225 ;
        RECT 60.210 141.865 60.950 141.895 ;
        RECT 60.210 141.565 61.125 141.865 ;
        RECT 60.800 141.390 61.125 141.565 ;
        RECT 59.830 140.835 60.085 141.365 ;
        RECT 60.805 141.035 61.125 141.390 ;
        RECT 61.295 141.605 61.835 141.975 ;
        RECT 62.170 141.885 62.575 142.055 ;
        RECT 61.295 141.205 61.535 141.605 ;
        RECT 62.015 141.435 62.235 141.715 ;
        RECT 61.705 141.265 62.235 141.435 ;
        RECT 61.705 141.035 61.875 141.265 ;
        RECT 60.805 140.865 61.875 141.035 ;
        RECT 62.405 141.105 62.575 141.885 ;
        RECT 62.745 141.275 63.095 141.895 ;
        RECT 63.265 141.275 63.475 142.065 ;
        RECT 63.665 142.095 65.165 142.265 ;
        RECT 63.665 141.405 63.835 142.095 ;
        RECT 65.525 141.925 65.695 142.705 ;
        RECT 66.500 142.575 66.670 142.705 ;
        RECT 64.005 141.755 65.695 141.925 ;
        RECT 65.865 142.145 66.330 142.535 ;
        RECT 66.500 142.405 66.895 142.575 ;
        RECT 64.005 141.575 64.175 141.755 ;
        RECT 62.405 140.825 63.355 141.105 ;
        RECT 63.665 141.015 63.925 141.405 ;
        RECT 64.345 141.335 65.135 141.585 ;
        RECT 63.575 140.845 63.925 141.015 ;
        RECT 65.340 141.045 65.510 141.755 ;
        RECT 65.865 141.555 66.035 142.145 ;
        RECT 65.680 141.335 66.035 141.555 ;
        RECT 66.205 141.335 66.555 141.955 ;
        RECT 66.725 141.045 66.895 142.405 ;
        RECT 67.260 142.235 67.585 143.020 ;
        RECT 67.065 141.185 67.525 142.235 ;
        RECT 65.340 140.875 66.195 141.045 ;
        RECT 66.400 140.875 66.895 141.045 ;
        RECT 67.755 140.915 67.925 143.035 ;
        RECT 68.595 142.535 68.850 143.035 ;
        RECT 68.100 142.365 68.850 142.535 ;
        RECT 68.100 141.375 68.330 142.365 ;
        RECT 68.500 141.545 68.850 142.195 ;
        RECT 69.025 142.130 69.295 143.035 ;
        RECT 69.975 142.275 70.145 143.035 ;
        RECT 68.100 141.205 68.850 141.375 ;
        RECT 68.595 140.915 68.850 141.205 ;
        RECT 69.025 141.330 69.195 142.130 ;
        RECT 69.480 142.105 70.145 142.275 ;
        RECT 69.480 141.960 69.650 142.105 ;
        RECT 72.225 142.055 72.555 143.035 ;
        RECT 108.590 142.695 110.245 142.985 ;
        RECT 108.590 142.355 110.180 142.525 ;
        RECT 108.590 142.065 108.910 142.355 ;
        RECT 110.010 142.235 110.180 142.355 ;
        RECT 69.365 141.630 69.650 141.960 ;
        RECT 69.480 141.375 69.650 141.630 ;
        RECT 69.885 141.555 70.215 141.925 ;
        RECT 71.805 141.645 72.135 141.895 ;
        RECT 72.305 141.455 72.555 142.055 ;
        RECT 109.105 142.015 109.820 142.185 ;
        RECT 110.010 142.065 110.735 142.235 ;
        RECT 110.905 142.065 111.175 143.035 ;
        RECT 117.035 142.865 119.065 143.035 ;
        RECT 69.025 140.825 69.285 141.330 ;
        RECT 69.480 141.205 70.145 141.375 ;
        RECT 69.975 140.825 70.145 141.205 ;
        RECT 72.225 140.825 72.555 141.455 ;
        RECT 108.590 141.325 108.940 141.895 ;
        RECT 109.110 141.565 109.820 142.015 ;
        RECT 110.565 141.895 110.735 142.065 ;
        RECT 109.990 141.565 110.395 141.895 ;
        RECT 110.565 141.565 110.835 141.895 ;
        RECT 110.565 141.395 110.735 141.565 ;
        RECT 109.125 141.225 110.735 141.395 ;
        RECT 111.005 141.330 111.175 142.065 ;
        RECT 115.945 142.445 116.460 142.855 ;
        RECT 115.945 141.635 116.285 142.445 ;
        RECT 117.035 142.200 117.205 142.865 ;
        RECT 117.600 142.525 118.725 142.695 ;
        RECT 116.455 142.010 117.205 142.200 ;
        RECT 117.375 142.185 118.385 142.355 ;
        RECT 115.945 141.465 117.175 141.635 ;
        RECT 109.125 140.875 109.295 141.225 ;
        RECT 109.995 140.875 110.165 141.225 ;
        RECT 110.905 140.985 111.175 141.330 ;
        RECT 116.220 140.860 116.465 141.465 ;
        RECT 117.375 140.825 117.565 142.185 ;
        RECT 117.735 141.845 118.010 141.985 ;
        RECT 117.735 141.675 118.015 141.845 ;
        RECT 117.735 140.825 118.010 141.675 ;
        RECT 118.215 141.385 118.385 142.185 ;
        RECT 118.555 141.395 118.725 142.525 ;
        RECT 118.895 141.895 119.065 142.865 ;
        RECT 119.575 142.065 119.910 143.035 ;
        RECT 118.895 141.565 119.090 141.895 ;
        RECT 119.315 141.565 119.570 141.895 ;
        RECT 119.315 141.395 119.485 141.565 ;
        RECT 119.740 141.395 119.910 142.065 ;
        RECT 120.525 142.055 120.855 143.035 ;
        RECT 120.105 141.645 120.435 141.895 ;
        RECT 120.605 141.455 120.855 142.055 ;
        RECT 118.555 141.225 119.485 141.395 ;
        RECT 118.555 141.190 118.730 141.225 ;
        RECT 118.200 140.825 118.730 141.190 ;
        RECT 119.655 140.825 119.910 141.395 ;
        RECT 120.525 140.825 120.855 141.455 ;
        RECT 16.500 139.775 16.755 140.305 ;
        RECT 16.500 138.915 16.680 139.775 ;
        RECT 17.400 139.575 17.650 140.225 ;
        RECT 16.850 139.245 17.650 139.575 ;
        RECT 16.500 138.445 16.755 138.915 ;
        RECT 16.415 138.275 16.755 138.445 ;
        RECT 16.500 138.245 16.755 138.275 ;
        RECT 17.400 138.655 17.650 139.245 ;
        RECT 17.850 139.890 18.170 140.220 ;
        RECT 19.210 140.095 20.060 140.265 ;
        RECT 17.850 138.995 18.040 139.890 ;
        RECT 18.360 139.565 19.020 139.835 ;
        RECT 18.690 139.505 19.020 139.565 ;
        RECT 18.210 139.335 18.540 139.395 ;
        RECT 19.210 139.335 19.380 140.095 ;
        RECT 21.140 139.845 21.390 140.275 ;
        RECT 19.550 139.675 20.800 139.845 ;
        RECT 19.550 139.555 19.880 139.675 ;
        RECT 18.210 139.165 20.110 139.335 ;
        RECT 17.850 138.825 19.770 138.995 ;
        RECT 17.850 138.805 18.170 138.825 ;
        RECT 17.400 138.145 17.730 138.655 ;
        RECT 18.000 138.195 18.170 138.805 ;
        RECT 19.940 138.655 20.110 139.165 ;
        RECT 20.280 139.095 20.460 139.505 ;
        RECT 20.630 138.915 20.800 139.675 ;
        RECT 18.900 138.485 20.110 138.655 ;
        RECT 20.280 138.605 20.800 138.915 ;
        RECT 20.970 139.505 21.390 139.845 ;
        RECT 22.260 140.105 23.275 140.305 ;
        RECT 21.680 139.505 22.090 139.835 ;
        RECT 20.970 138.735 21.160 139.505 ;
        RECT 22.260 139.375 22.430 140.105 ;
        RECT 23.575 139.935 23.745 140.265 ;
        RECT 22.600 139.555 22.950 139.925 ;
        RECT 22.260 139.335 22.680 139.375 ;
        RECT 21.330 139.165 22.680 139.335 ;
        RECT 21.330 139.005 21.580 139.165 ;
        RECT 22.090 138.735 22.340 138.995 ;
        RECT 20.970 138.485 22.340 138.735 ;
        RECT 18.900 138.195 19.140 138.485 ;
        RECT 19.940 138.405 20.110 138.485 ;
        RECT 19.940 138.155 20.570 138.405 ;
        RECT 21.540 138.195 21.710 138.485 ;
        RECT 22.510 138.320 22.680 139.165 ;
        RECT 23.130 138.995 23.350 139.865 ;
        RECT 23.575 139.745 24.270 139.935 ;
        RECT 22.850 138.615 23.350 138.995 ;
        RECT 23.520 138.945 23.930 139.565 ;
        RECT 24.100 138.775 24.270 139.745 ;
        RECT 23.575 138.605 24.270 138.775 ;
        RECT 22.510 138.150 23.340 138.320 ;
        RECT 23.575 138.105 23.745 138.605 ;
        RECT 24.460 138.105 24.685 140.225 ;
        RECT 25.355 139.935 25.525 140.225 ;
        RECT 24.860 139.765 25.525 139.935 ;
        RECT 34.265 139.855 34.595 140.215 ;
        RECT 35.635 140.025 36.195 140.315 ;
        RECT 24.860 138.775 25.090 139.765 ;
        RECT 34.265 139.665 35.655 139.855 ;
        RECT 25.260 138.945 25.610 139.595 ;
        RECT 35.485 139.575 35.655 139.665 ;
        RECT 34.080 139.245 34.755 139.495 ;
        RECT 34.975 139.245 35.315 139.495 ;
        RECT 35.485 139.245 35.775 139.575 ;
        RECT 34.080 138.885 34.345 139.245 ;
        RECT 35.485 138.995 35.655 139.245 ;
        RECT 34.715 138.825 35.655 138.995 ;
        RECT 24.860 138.605 25.525 138.775 ;
        RECT 25.355 138.105 25.525 138.605 ;
        RECT 34.715 138.275 35.015 138.825 ;
        RECT 35.945 138.655 36.195 140.025 ;
        RECT 35.735 138.105 36.195 138.655 ;
        RECT 38.665 139.810 38.935 140.155 ;
        RECT 39.675 139.915 39.845 140.265 ;
        RECT 40.545 139.915 40.715 140.265 ;
        RECT 38.665 139.075 38.835 139.810 ;
        RECT 39.105 139.745 40.715 139.915 ;
        RECT 47.485 139.915 47.655 140.265 ;
        RECT 48.355 139.915 48.525 140.265 ;
        RECT 39.105 139.575 39.275 139.745 ;
        RECT 39.005 139.245 39.275 139.575 ;
        RECT 39.445 139.245 39.850 139.575 ;
        RECT 39.105 139.075 39.275 139.245 ;
        RECT 38.665 138.105 38.935 139.075 ;
        RECT 39.105 138.905 39.830 139.075 ;
        RECT 40.020 138.955 40.730 139.575 ;
        RECT 40.900 139.245 41.250 139.815 ;
        RECT 46.950 139.245 47.300 139.815 ;
        RECT 47.485 139.745 49.095 139.915 ;
        RECT 49.265 139.810 49.535 140.155 ;
        RECT 48.925 139.575 49.095 139.745 ;
        RECT 47.470 139.125 48.180 139.575 ;
        RECT 48.350 139.245 48.755 139.575 ;
        RECT 48.925 139.245 49.195 139.575 ;
        RECT 39.660 138.785 39.830 138.905 ;
        RECT 40.930 138.785 41.250 139.075 ;
        RECT 39.660 138.615 41.250 138.785 ;
        RECT 46.950 138.785 47.270 139.075 ;
        RECT 47.465 138.955 48.180 139.125 ;
        RECT 48.925 139.075 49.095 139.245 ;
        RECT 49.365 139.075 49.535 139.810 ;
        RECT 48.370 138.905 49.095 139.075 ;
        RECT 48.370 138.785 48.540 138.905 ;
        RECT 46.950 138.615 48.540 138.785 ;
        RECT 39.595 138.155 41.250 138.445 ;
        RECT 46.950 138.155 48.605 138.445 ;
        RECT 49.265 138.105 49.535 139.075 ;
        RECT 49.705 139.685 50.045 140.315 ;
        RECT 50.655 139.835 50.985 140.315 ;
        RECT 51.550 139.835 51.880 140.315 ;
        RECT 49.705 139.635 49.935 139.685 ;
        RECT 50.655 139.665 51.880 139.835 ;
        RECT 52.510 139.705 53.010 140.315 ;
        RECT 49.705 139.075 49.880 139.635 ;
        RECT 50.050 139.325 50.745 139.495 ;
        RECT 50.575 139.075 50.745 139.325 ;
        RECT 50.920 139.295 51.340 139.495 ;
        RECT 51.510 139.295 51.840 139.495 ;
        RECT 52.010 139.295 52.340 139.495 ;
        RECT 52.510 139.075 52.680 139.705 ;
        RECT 55.665 139.685 55.995 140.315 ;
        RECT 52.865 139.245 53.215 139.495 ;
        RECT 55.245 139.245 55.575 139.495 ;
        RECT 55.745 139.085 55.995 139.685 ;
        RECT 49.705 138.105 50.045 139.075 ;
        RECT 50.575 138.905 53.010 139.075 ;
        RECT 51.550 138.105 51.880 138.905 ;
        RECT 52.680 138.105 53.010 138.905 ;
        RECT 55.665 138.105 55.995 139.085 ;
        RECT 59.365 139.685 59.705 140.315 ;
        RECT 60.315 139.835 60.645 140.315 ;
        RECT 61.210 139.835 61.540 140.315 ;
        RECT 59.365 139.075 59.540 139.685 ;
        RECT 60.315 139.665 61.540 139.835 ;
        RECT 62.170 139.705 62.670 140.315 ;
        RECT 59.710 139.325 60.405 139.495 ;
        RECT 60.235 139.075 60.405 139.325 ;
        RECT 60.580 139.295 61.000 139.495 ;
        RECT 61.170 139.295 61.500 139.495 ;
        RECT 61.670 139.295 62.000 139.495 ;
        RECT 62.170 139.075 62.340 139.705 ;
        RECT 63.965 139.685 64.305 140.315 ;
        RECT 64.915 139.835 65.245 140.315 ;
        RECT 65.810 139.835 66.140 140.315 ;
        RECT 62.525 139.245 62.875 139.495 ;
        RECT 63.965 139.075 64.140 139.685 ;
        RECT 64.915 139.665 66.140 139.835 ;
        RECT 66.770 139.705 67.270 140.315 ;
        RECT 67.735 139.935 67.905 140.225 ;
        RECT 67.735 139.765 68.400 139.935 ;
        RECT 64.310 139.325 65.005 139.495 ;
        RECT 64.835 139.075 65.005 139.325 ;
        RECT 65.180 139.295 65.600 139.495 ;
        RECT 65.770 139.295 66.100 139.495 ;
        RECT 66.270 139.295 66.600 139.495 ;
        RECT 66.770 139.075 66.940 139.705 ;
        RECT 67.125 139.245 67.475 139.495 ;
        RECT 59.365 138.105 59.705 139.075 ;
        RECT 60.235 138.905 62.670 139.075 ;
        RECT 61.210 138.105 61.540 138.905 ;
        RECT 62.340 138.105 62.670 138.905 ;
        RECT 63.965 138.105 64.305 139.075 ;
        RECT 64.835 138.905 67.270 139.075 ;
        RECT 67.650 138.945 68.000 139.595 ;
        RECT 65.810 138.105 66.140 138.905 ;
        RECT 66.940 138.105 67.270 138.905 ;
        RECT 68.170 138.775 68.400 139.765 ;
        RECT 67.735 138.605 68.400 138.775 ;
        RECT 67.735 138.105 67.905 138.605 ;
        RECT 68.575 138.105 68.800 140.225 ;
        RECT 69.515 139.935 69.685 140.265 ;
        RECT 69.985 140.105 71.000 140.305 ;
        RECT 68.990 139.745 69.685 139.935 ;
        RECT 68.990 138.775 69.160 139.745 ;
        RECT 69.330 138.945 69.740 139.565 ;
        RECT 69.910 138.995 70.130 139.865 ;
        RECT 70.310 139.555 70.660 139.925 ;
        RECT 70.830 139.375 71.000 140.105 ;
        RECT 71.870 139.845 72.120 140.275 ;
        RECT 73.200 140.095 74.050 140.265 ;
        RECT 71.170 139.505 71.580 139.835 ;
        RECT 71.870 139.505 72.290 139.845 ;
        RECT 70.580 139.335 71.000 139.375 ;
        RECT 70.580 139.165 71.930 139.335 ;
        RECT 68.990 138.605 69.685 138.775 ;
        RECT 69.910 138.615 70.410 138.995 ;
        RECT 69.515 138.105 69.685 138.605 ;
        RECT 70.580 138.320 70.750 139.165 ;
        RECT 71.680 139.005 71.930 139.165 ;
        RECT 70.920 138.735 71.170 138.995 ;
        RECT 72.100 138.735 72.290 139.505 ;
        RECT 70.920 138.485 72.290 138.735 ;
        RECT 72.460 139.675 73.710 139.845 ;
        RECT 72.460 138.915 72.630 139.675 ;
        RECT 73.380 139.555 73.710 139.675 ;
        RECT 72.800 139.095 72.980 139.505 ;
        RECT 73.880 139.335 74.050 140.095 ;
        RECT 75.090 139.890 75.410 140.220 ;
        RECT 74.240 139.565 74.900 139.835 ;
        RECT 74.240 139.505 74.570 139.565 ;
        RECT 74.720 139.335 75.050 139.395 ;
        RECT 73.150 139.165 75.050 139.335 ;
        RECT 72.460 138.605 72.980 138.915 ;
        RECT 73.150 138.655 73.320 139.165 ;
        RECT 75.220 138.995 75.410 139.890 ;
        RECT 73.490 138.825 75.410 138.995 ;
        RECT 75.090 138.805 75.410 138.825 ;
        RECT 75.610 139.575 75.860 140.225 ;
        RECT 76.505 139.775 76.760 140.305 ;
        RECT 75.610 139.245 76.410 139.575 ;
        RECT 73.150 138.485 74.360 138.655 ;
        RECT 69.920 138.150 70.750 138.320 ;
        RECT 71.550 138.195 71.720 138.485 ;
        RECT 73.150 138.405 73.320 138.485 ;
        RECT 72.690 138.155 73.320 138.405 ;
        RECT 74.120 138.195 74.360 138.485 ;
        RECT 75.090 138.195 75.260 138.805 ;
        RECT 75.610 138.655 75.860 139.245 ;
        RECT 76.580 138.915 76.760 139.775 ;
        RECT 75.530 138.145 75.860 138.655 ;
        RECT 76.505 138.445 76.760 138.915 ;
        RECT 80.065 139.685 80.405 140.315 ;
        RECT 81.015 139.835 81.345 140.315 ;
        RECT 81.910 139.835 82.240 140.315 ;
        RECT 80.065 139.075 80.240 139.685 ;
        RECT 81.015 139.665 82.240 139.835 ;
        RECT 82.870 139.705 83.370 140.315 ;
        RECT 80.410 139.325 81.105 139.495 ;
        RECT 80.935 139.075 81.105 139.325 ;
        RECT 81.280 139.295 81.700 139.495 ;
        RECT 81.870 139.295 82.200 139.495 ;
        RECT 82.370 139.295 82.700 139.495 ;
        RECT 82.870 139.075 83.040 139.705 ;
        RECT 84.940 139.675 85.185 140.280 ;
        RECT 84.665 139.505 85.895 139.675 ;
        RECT 83.225 139.245 83.575 139.495 ;
        RECT 76.505 138.275 76.845 138.445 ;
        RECT 76.505 138.245 76.760 138.275 ;
        RECT 80.065 138.105 80.405 139.075 ;
        RECT 80.935 138.905 83.370 139.075 ;
        RECT 81.910 138.105 82.240 138.905 ;
        RECT 83.040 138.105 83.370 138.905 ;
        RECT 84.665 138.695 85.005 139.505 ;
        RECT 85.175 138.940 85.925 139.130 ;
        RECT 84.665 138.285 85.180 138.695 ;
        RECT 85.755 138.275 85.925 138.940 ;
        RECT 86.095 138.955 86.285 140.315 ;
        RECT 86.455 139.465 86.730 140.315 ;
        RECT 86.920 139.950 87.450 140.315 ;
        RECT 87.275 139.915 87.450 139.950 ;
        RECT 86.455 139.295 86.735 139.465 ;
        RECT 86.455 139.155 86.730 139.295 ;
        RECT 86.935 138.955 87.105 139.755 ;
        RECT 86.095 138.785 87.105 138.955 ;
        RECT 87.275 139.745 88.205 139.915 ;
        RECT 88.375 139.745 88.630 140.315 ;
        RECT 89.815 139.935 89.985 140.315 ;
        RECT 89.815 139.765 90.480 139.935 ;
        RECT 90.675 139.810 90.935 140.315 ;
        RECT 87.275 138.615 87.445 139.745 ;
        RECT 88.035 139.575 88.205 139.745 ;
        RECT 86.320 138.445 87.445 138.615 ;
        RECT 87.615 139.245 87.810 139.575 ;
        RECT 88.035 139.245 88.290 139.575 ;
        RECT 87.615 138.275 87.785 139.245 ;
        RECT 88.460 139.075 88.630 139.745 ;
        RECT 89.745 139.215 90.075 139.585 ;
        RECT 90.310 139.510 90.480 139.765 ;
        RECT 85.755 138.105 87.785 138.275 ;
        RECT 88.295 138.105 88.630 139.075 ;
        RECT 90.310 139.180 90.595 139.510 ;
        RECT 90.310 139.035 90.480 139.180 ;
        RECT 89.815 138.865 90.480 139.035 ;
        RECT 90.765 139.010 90.935 139.810 ;
        RECT 101.665 139.685 101.995 140.315 ;
        RECT 101.245 139.245 101.575 139.495 ;
        RECT 101.745 139.085 101.995 139.685 ;
        RECT 89.815 138.105 89.985 138.865 ;
        RECT 90.665 138.105 90.935 139.010 ;
        RECT 101.665 138.105 101.995 139.085 ;
        RECT 106.285 139.685 106.625 140.315 ;
        RECT 107.235 139.835 107.565 140.315 ;
        RECT 108.130 139.835 108.460 140.315 ;
        RECT 106.285 139.635 106.515 139.685 ;
        RECT 107.235 139.665 108.460 139.835 ;
        RECT 109.090 139.705 109.590 140.315 ;
        RECT 110.170 139.705 110.670 140.315 ;
        RECT 106.285 139.075 106.460 139.635 ;
        RECT 106.630 139.325 107.325 139.495 ;
        RECT 107.155 139.075 107.325 139.325 ;
        RECT 107.500 139.295 107.920 139.495 ;
        RECT 108.090 139.295 108.420 139.495 ;
        RECT 108.590 139.295 108.920 139.495 ;
        RECT 109.090 139.075 109.260 139.705 ;
        RECT 109.445 139.245 109.795 139.495 ;
        RECT 109.965 139.245 110.315 139.495 ;
        RECT 110.500 139.075 110.670 139.705 ;
        RECT 111.300 139.835 111.630 140.315 ;
        RECT 112.195 139.835 112.525 140.315 ;
        RECT 111.300 139.665 112.525 139.835 ;
        RECT 113.135 139.685 113.475 140.315 ;
        RECT 115.925 139.685 116.255 140.315 ;
        RECT 113.245 139.635 113.475 139.685 ;
        RECT 110.840 139.295 111.170 139.495 ;
        RECT 111.340 139.295 111.670 139.495 ;
        RECT 111.840 139.295 112.260 139.495 ;
        RECT 112.435 139.325 113.130 139.495 ;
        RECT 112.435 139.075 112.605 139.325 ;
        RECT 113.300 139.075 113.475 139.635 ;
        RECT 115.505 139.245 115.835 139.495 ;
        RECT 116.005 139.085 116.255 139.685 ;
        RECT 106.285 138.105 106.625 139.075 ;
        RECT 107.155 138.905 109.590 139.075 ;
        RECT 108.130 138.105 108.460 138.905 ;
        RECT 109.260 138.105 109.590 138.905 ;
        RECT 110.170 138.905 112.605 139.075 ;
        RECT 110.170 138.105 110.500 138.905 ;
        RECT 111.300 138.105 111.630 138.905 ;
        RECT 113.135 138.105 113.475 139.075 ;
        RECT 115.925 138.105 116.255 139.085 ;
        RECT 117.240 139.775 117.495 140.305 ;
        RECT 117.240 138.915 117.420 139.775 ;
        RECT 118.140 139.575 118.390 140.225 ;
        RECT 117.590 139.245 118.390 139.575 ;
        RECT 117.240 138.785 117.495 138.915 ;
        RECT 117.155 138.615 117.495 138.785 ;
        RECT 117.240 138.245 117.495 138.615 ;
        RECT 118.140 138.655 118.390 139.245 ;
        RECT 118.590 139.890 118.910 140.220 ;
        RECT 119.950 140.095 120.800 140.265 ;
        RECT 118.590 138.995 118.780 139.890 ;
        RECT 119.100 139.565 119.760 139.835 ;
        RECT 119.430 139.505 119.760 139.565 ;
        RECT 118.950 139.335 119.280 139.395 ;
        RECT 119.950 139.335 120.120 140.095 ;
        RECT 121.880 139.845 122.130 140.275 ;
        RECT 120.290 139.675 121.540 139.845 ;
        RECT 120.290 139.555 120.620 139.675 ;
        RECT 118.950 139.165 120.850 139.335 ;
        RECT 118.590 138.825 120.510 138.995 ;
        RECT 118.590 138.805 118.910 138.825 ;
        RECT 118.140 138.145 118.470 138.655 ;
        RECT 118.740 138.195 118.910 138.805 ;
        RECT 120.680 138.655 120.850 139.165 ;
        RECT 121.020 139.095 121.200 139.505 ;
        RECT 121.370 138.915 121.540 139.675 ;
        RECT 119.640 138.485 120.850 138.655 ;
        RECT 121.020 138.605 121.540 138.915 ;
        RECT 121.710 139.505 122.130 139.845 ;
        RECT 123.000 140.105 124.015 140.305 ;
        RECT 122.420 139.505 122.830 139.835 ;
        RECT 121.710 138.735 121.900 139.505 ;
        RECT 123.000 139.375 123.170 140.105 ;
        RECT 124.315 139.935 124.485 140.265 ;
        RECT 123.340 139.555 123.690 139.925 ;
        RECT 123.000 139.335 123.420 139.375 ;
        RECT 122.070 139.165 123.420 139.335 ;
        RECT 122.070 139.005 122.320 139.165 ;
        RECT 122.830 138.735 123.080 138.995 ;
        RECT 121.710 138.485 123.080 138.735 ;
        RECT 119.640 138.195 119.880 138.485 ;
        RECT 120.680 138.405 120.850 138.485 ;
        RECT 120.680 138.155 121.310 138.405 ;
        RECT 122.280 138.195 122.450 138.485 ;
        RECT 123.250 138.320 123.420 139.165 ;
        RECT 123.870 138.995 124.090 139.865 ;
        RECT 124.315 139.745 125.010 139.935 ;
        RECT 123.590 138.615 124.090 138.995 ;
        RECT 124.260 138.945 124.670 139.565 ;
        RECT 124.840 138.775 125.010 139.745 ;
        RECT 124.315 138.605 125.010 138.775 ;
        RECT 123.250 138.150 124.080 138.320 ;
        RECT 124.315 138.105 124.485 138.605 ;
        RECT 125.200 138.105 125.425 140.225 ;
        RECT 126.095 139.935 126.265 140.225 ;
        RECT 125.600 139.765 126.265 139.935 ;
        RECT 125.600 138.775 125.830 139.765 ;
        RECT 126.000 138.945 126.350 139.595 ;
        RECT 125.600 138.605 126.265 138.775 ;
        RECT 126.095 138.105 126.265 138.605 ;
        RECT 21.735 136.835 21.905 137.595 ;
        RECT 21.735 136.665 22.400 136.835 ;
        RECT 22.585 136.690 22.855 137.595 ;
        RECT 22.230 136.520 22.400 136.665 ;
        RECT 21.665 136.115 21.995 136.485 ;
        RECT 22.230 136.190 22.515 136.520 ;
        RECT 22.230 135.935 22.400 136.190 ;
        RECT 21.735 135.765 22.400 135.935 ;
        RECT 22.685 135.890 22.855 136.690 ;
        RECT 23.465 136.615 23.795 137.595 ;
        RECT 30.095 137.425 32.125 137.595 ;
        RECT 23.045 136.205 23.375 136.455 ;
        RECT 23.545 136.015 23.795 136.615 ;
        RECT 29.005 137.005 29.520 137.415 ;
        RECT 29.005 136.195 29.345 137.005 ;
        RECT 30.095 136.760 30.265 137.425 ;
        RECT 30.660 137.085 31.785 137.255 ;
        RECT 29.515 136.570 30.265 136.760 ;
        RECT 30.435 136.745 31.445 136.915 ;
        RECT 29.005 136.025 30.235 136.195 ;
        RECT 21.735 135.385 21.905 135.765 ;
        RECT 22.595 135.385 22.855 135.890 ;
        RECT 23.465 135.385 23.795 136.015 ;
        RECT 29.280 135.420 29.525 136.025 ;
        RECT 30.435 135.385 30.625 136.745 ;
        RECT 30.795 135.725 31.070 136.545 ;
        RECT 31.275 135.945 31.445 136.745 ;
        RECT 31.615 135.955 31.785 137.085 ;
        RECT 31.955 136.455 32.125 137.425 ;
        RECT 32.635 136.625 32.970 137.595 ;
        RECT 31.955 136.125 32.150 136.455 ;
        RECT 32.375 136.125 32.630 136.455 ;
        RECT 32.375 135.955 32.545 136.125 ;
        RECT 32.800 135.955 32.970 136.625 ;
        RECT 31.615 135.785 32.545 135.955 ;
        RECT 31.615 135.750 31.790 135.785 ;
        RECT 30.795 135.555 31.075 135.725 ;
        RECT 30.795 135.385 31.070 135.555 ;
        RECT 31.260 135.385 31.790 135.750 ;
        RECT 32.715 135.385 32.970 135.955 ;
        RECT 34.985 136.625 35.255 137.595 ;
        RECT 35.915 137.255 37.570 137.545 ;
        RECT 35.980 136.915 37.570 137.085 ;
        RECT 35.980 136.795 36.150 136.915 ;
        RECT 35.425 136.625 36.150 136.795 ;
        RECT 34.985 135.890 35.155 136.625 ;
        RECT 35.425 136.455 35.595 136.625 ;
        RECT 35.325 136.125 35.595 136.455 ;
        RECT 35.765 136.125 36.170 136.455 ;
        RECT 36.340 136.125 37.050 136.745 ;
        RECT 37.250 136.625 37.570 136.915 ;
        RECT 38.395 136.875 38.695 137.425 ;
        RECT 39.415 137.045 39.875 137.595 ;
        RECT 37.760 136.455 38.025 136.815 ;
        RECT 38.395 136.705 39.335 136.875 ;
        RECT 39.165 136.455 39.335 136.705 ;
        RECT 35.425 135.955 35.595 136.125 ;
        RECT 34.985 135.545 35.255 135.890 ;
        RECT 35.425 135.785 37.035 135.955 ;
        RECT 37.220 135.885 37.570 136.455 ;
        RECT 37.760 136.205 38.435 136.455 ;
        RECT 38.655 136.205 38.995 136.455 ;
        RECT 39.165 136.125 39.455 136.455 ;
        RECT 39.165 136.035 39.335 136.125 ;
        RECT 35.995 135.435 36.165 135.785 ;
        RECT 36.865 135.435 37.035 135.785 ;
        RECT 37.945 135.845 39.335 136.035 ;
        RECT 37.945 135.485 38.275 135.845 ;
        RECT 39.625 135.675 39.875 137.045 ;
        RECT 39.315 135.385 39.875 135.675 ;
        RECT 43.725 136.625 43.995 137.595 ;
        RECT 44.655 137.255 46.310 137.545 ;
        RECT 54.015 137.425 56.045 137.595 ;
        RECT 44.720 136.915 46.310 137.085 ;
        RECT 44.720 136.795 44.890 136.915 ;
        RECT 44.165 136.625 44.890 136.795 ;
        RECT 43.725 135.890 43.895 136.625 ;
        RECT 44.165 136.455 44.335 136.625 ;
        RECT 45.080 136.575 45.795 136.745 ;
        RECT 45.990 136.625 46.310 136.915 ;
        RECT 52.925 137.005 53.440 137.415 ;
        RECT 44.065 136.125 44.335 136.455 ;
        RECT 44.505 136.125 44.910 136.455 ;
        RECT 45.080 136.125 45.790 136.575 ;
        RECT 44.165 135.955 44.335 136.125 ;
        RECT 43.725 135.545 43.995 135.890 ;
        RECT 44.165 135.785 45.775 135.955 ;
        RECT 45.960 135.885 46.310 136.455 ;
        RECT 52.925 136.195 53.265 137.005 ;
        RECT 54.015 136.760 54.185 137.425 ;
        RECT 54.580 137.085 55.705 137.255 ;
        RECT 53.435 136.570 54.185 136.760 ;
        RECT 54.355 136.745 55.365 136.915 ;
        RECT 52.925 136.025 54.155 136.195 ;
        RECT 44.735 135.435 44.905 135.785 ;
        RECT 45.605 135.435 45.775 135.785 ;
        RECT 53.200 135.420 53.445 136.025 ;
        RECT 54.355 135.385 54.545 136.745 ;
        RECT 54.715 136.405 54.990 136.545 ;
        RECT 54.715 136.235 54.995 136.405 ;
        RECT 54.715 135.385 54.990 136.235 ;
        RECT 55.195 135.945 55.365 136.745 ;
        RECT 55.535 135.955 55.705 137.085 ;
        RECT 55.875 136.455 56.045 137.425 ;
        RECT 56.555 136.625 56.890 137.595 ;
        RECT 57.615 136.835 57.785 137.595 ;
        RECT 57.615 136.665 58.280 136.835 ;
        RECT 58.465 136.690 58.735 137.595 ;
        RECT 55.875 136.125 56.070 136.455 ;
        RECT 56.295 136.125 56.550 136.455 ;
        RECT 56.295 135.955 56.465 136.125 ;
        RECT 56.720 135.955 56.890 136.625 ;
        RECT 58.110 136.520 58.280 136.665 ;
        RECT 57.545 136.115 57.875 136.485 ;
        RECT 58.110 136.190 58.395 136.520 ;
        RECT 55.535 135.785 56.465 135.955 ;
        RECT 55.535 135.750 55.710 135.785 ;
        RECT 55.180 135.385 55.710 135.750 ;
        RECT 56.635 135.385 56.890 135.955 ;
        RECT 58.110 135.935 58.280 136.190 ;
        RECT 57.615 135.765 58.280 135.935 ;
        RECT 58.565 135.890 58.735 136.690 ;
        RECT 57.615 135.385 57.785 135.765 ;
        RECT 58.475 135.385 58.735 135.890 ;
        RECT 61.205 136.625 61.545 137.595 ;
        RECT 63.050 136.795 63.380 137.595 ;
        RECT 64.180 136.795 64.510 137.595 ;
        RECT 62.075 136.625 64.510 136.795 ;
        RECT 67.185 136.915 67.445 137.595 ;
        RECT 68.115 137.215 68.365 137.595 ;
        RECT 69.895 137.375 70.230 137.595 ;
        RECT 69.495 137.215 69.725 137.255 ;
        RECT 68.115 137.015 69.725 137.215 ;
        RECT 68.115 137.005 68.950 137.015 ;
        RECT 69.540 136.925 69.725 137.015 ;
        RECT 61.205 136.065 61.380 136.625 ;
        RECT 62.075 136.375 62.245 136.625 ;
        RECT 61.550 136.205 62.245 136.375 ;
        RECT 62.420 136.205 62.840 136.405 ;
        RECT 63.010 136.205 63.340 136.405 ;
        RECT 63.510 136.205 63.840 136.405 ;
        RECT 61.205 136.015 61.435 136.065 ;
        RECT 61.205 135.385 61.545 136.015 ;
        RECT 62.155 135.865 63.380 136.035 ;
        RECT 62.155 135.385 62.485 135.865 ;
        RECT 63.050 135.385 63.380 135.865 ;
        RECT 64.010 135.995 64.180 136.625 ;
        RECT 64.365 136.205 64.715 136.455 ;
        RECT 64.010 135.385 64.510 135.995 ;
        RECT 67.185 135.715 67.355 136.915 ;
        RECT 69.055 136.815 69.385 136.845 ;
        RECT 67.585 136.755 69.385 136.815 ;
        RECT 69.975 136.755 70.230 137.375 ;
        RECT 67.525 136.645 70.230 136.755 ;
        RECT 67.525 136.610 67.725 136.645 ;
        RECT 67.525 136.035 67.695 136.610 ;
        RECT 69.055 136.585 70.230 136.645 ;
        RECT 70.405 136.625 70.790 137.595 ;
        RECT 71.805 137.135 72.085 137.595 ;
        RECT 70.960 136.915 72.085 137.135 ;
        RECT 67.925 136.170 68.335 136.475 ;
        RECT 68.505 136.205 68.835 136.415 ;
        RECT 67.525 135.915 67.795 136.035 ;
        RECT 67.525 135.870 68.370 135.915 ;
        RECT 67.615 135.745 68.370 135.870 ;
        RECT 68.625 135.805 68.835 136.205 ;
        RECT 69.080 136.205 69.555 136.415 ;
        RECT 69.745 136.205 70.235 136.405 ;
        RECT 69.080 135.805 69.300 136.205 ;
        RECT 70.405 135.955 70.685 136.625 ;
        RECT 70.960 136.455 71.410 136.915 ;
        RECT 72.275 136.745 72.675 137.595 ;
        RECT 73.515 137.135 73.800 137.595 ;
        RECT 70.855 136.125 71.410 136.455 ;
        RECT 71.580 136.185 72.675 136.745 ;
        RECT 70.960 136.015 71.410 136.125 ;
        RECT 67.185 135.385 67.445 135.715 ;
        RECT 68.200 135.595 68.370 135.745 ;
        RECT 68.200 135.385 69.500 135.595 ;
        RECT 70.405 135.385 70.790 135.955 ;
        RECT 70.960 135.845 72.085 136.015 ;
        RECT 71.805 135.385 72.085 135.845 ;
        RECT 72.275 135.385 72.675 136.185 ;
        RECT 72.845 136.915 73.800 137.135 ;
        RECT 72.845 136.015 73.055 136.915 ;
        RECT 73.225 136.185 73.915 136.745 ;
        RECT 77.305 136.625 77.575 137.595 ;
        RECT 78.235 137.255 79.890 137.545 ;
        RECT 78.300 136.915 79.890 137.085 ;
        RECT 78.300 136.795 78.470 136.915 ;
        RECT 77.745 136.625 78.470 136.795 ;
        RECT 72.845 135.845 73.800 136.015 ;
        RECT 73.515 135.385 73.800 135.845 ;
        RECT 77.305 135.890 77.475 136.625 ;
        RECT 77.745 136.455 77.915 136.625 ;
        RECT 78.660 136.575 79.375 136.745 ;
        RECT 79.570 136.625 79.890 136.915 ;
        RECT 80.065 136.625 80.405 137.595 ;
        RECT 81.910 136.795 82.240 137.595 ;
        RECT 83.040 136.795 83.370 137.595 ;
        RECT 84.120 137.425 84.375 137.455 ;
        RECT 84.035 137.255 84.375 137.425 ;
        RECT 80.935 136.625 83.370 136.795 ;
        RECT 84.120 136.785 84.375 137.255 ;
        RECT 85.020 137.045 85.350 137.555 ;
        RECT 77.645 136.125 77.915 136.455 ;
        RECT 78.085 136.125 78.490 136.455 ;
        RECT 78.660 136.125 79.370 136.575 ;
        RECT 77.745 135.955 77.915 136.125 ;
        RECT 77.305 135.545 77.575 135.890 ;
        RECT 77.745 135.785 79.355 135.955 ;
        RECT 79.540 135.885 79.890 136.455 ;
        RECT 80.065 136.015 80.240 136.625 ;
        RECT 80.935 136.375 81.105 136.625 ;
        RECT 80.410 136.205 81.105 136.375 ;
        RECT 81.280 136.205 81.700 136.405 ;
        RECT 81.870 136.205 82.200 136.405 ;
        RECT 82.370 136.205 82.700 136.405 ;
        RECT 78.315 135.435 78.485 135.785 ;
        RECT 79.185 135.435 79.355 135.785 ;
        RECT 80.065 135.385 80.405 136.015 ;
        RECT 81.015 135.865 82.240 136.035 ;
        RECT 81.015 135.385 81.345 135.865 ;
        RECT 81.910 135.385 82.240 135.865 ;
        RECT 82.870 135.995 83.040 136.625 ;
        RECT 83.225 136.205 83.575 136.455 ;
        RECT 82.870 135.385 83.370 135.995 ;
        RECT 84.120 135.925 84.300 136.785 ;
        RECT 85.020 136.455 85.270 137.045 ;
        RECT 85.620 136.895 85.790 137.505 ;
        RECT 86.520 137.215 86.760 137.505 ;
        RECT 87.560 137.295 88.190 137.545 ;
        RECT 87.560 137.215 87.730 137.295 ;
        RECT 89.160 137.215 89.330 137.505 ;
        RECT 90.130 137.380 90.960 137.550 ;
        RECT 86.520 137.045 87.730 137.215 ;
        RECT 84.470 136.125 85.270 136.455 ;
        RECT 84.120 135.395 84.375 135.925 ;
        RECT 85.020 135.475 85.270 136.125 ;
        RECT 85.470 136.875 85.790 136.895 ;
        RECT 85.470 136.705 87.390 136.875 ;
        RECT 85.470 135.810 85.660 136.705 ;
        RECT 87.560 136.535 87.730 137.045 ;
        RECT 87.900 136.785 88.420 137.095 ;
        RECT 85.830 136.365 87.730 136.535 ;
        RECT 85.830 136.305 86.160 136.365 ;
        RECT 86.310 136.135 86.640 136.195 ;
        RECT 85.980 135.865 86.640 136.135 ;
        RECT 85.470 135.480 85.790 135.810 ;
        RECT 86.830 135.605 87.000 136.365 ;
        RECT 87.900 136.195 88.080 136.605 ;
        RECT 87.170 136.025 87.500 136.145 ;
        RECT 88.250 136.025 88.420 136.785 ;
        RECT 87.170 135.855 88.420 136.025 ;
        RECT 88.590 136.965 89.960 137.215 ;
        RECT 88.590 136.195 88.780 136.965 ;
        RECT 89.710 136.705 89.960 136.965 ;
        RECT 88.950 136.535 89.200 136.695 ;
        RECT 90.130 136.535 90.300 137.380 ;
        RECT 91.195 137.095 91.365 137.595 ;
        RECT 90.470 136.705 90.970 137.085 ;
        RECT 91.195 136.925 91.890 137.095 ;
        RECT 88.950 136.365 90.300 136.535 ;
        RECT 89.880 136.325 90.300 136.365 ;
        RECT 88.590 135.855 89.010 136.195 ;
        RECT 89.300 135.865 89.710 136.195 ;
        RECT 86.830 135.435 87.680 135.605 ;
        RECT 88.760 135.425 89.010 135.855 ;
        RECT 89.880 135.595 90.050 136.325 ;
        RECT 90.220 135.775 90.570 136.145 ;
        RECT 90.750 135.835 90.970 136.705 ;
        RECT 91.140 136.135 91.550 136.755 ;
        RECT 91.720 135.955 91.890 136.925 ;
        RECT 91.195 135.765 91.890 135.955 ;
        RECT 89.880 135.395 90.895 135.595 ;
        RECT 91.195 135.435 91.365 135.765 ;
        RECT 92.080 135.475 92.305 137.595 ;
        RECT 92.975 137.095 93.145 137.595 ;
        RECT 94.495 137.425 96.525 137.595 ;
        RECT 92.480 136.925 93.145 137.095 ;
        RECT 93.405 137.005 93.920 137.415 ;
        RECT 92.480 135.935 92.710 136.925 ;
        RECT 92.880 136.105 93.230 136.755 ;
        RECT 93.405 136.195 93.745 137.005 ;
        RECT 94.495 136.760 94.665 137.425 ;
        RECT 95.060 137.085 96.185 137.255 ;
        RECT 93.915 136.570 94.665 136.760 ;
        RECT 94.835 136.745 95.845 136.915 ;
        RECT 93.405 136.025 94.635 136.195 ;
        RECT 92.480 135.765 93.145 135.935 ;
        RECT 92.975 135.475 93.145 135.765 ;
        RECT 93.680 135.420 93.925 136.025 ;
        RECT 94.835 135.385 95.025 136.745 ;
        RECT 95.195 136.405 95.470 136.545 ;
        RECT 95.195 136.235 95.475 136.405 ;
        RECT 95.195 135.385 95.470 136.235 ;
        RECT 95.675 135.945 95.845 136.745 ;
        RECT 96.015 135.955 96.185 137.085 ;
        RECT 96.355 136.455 96.525 137.425 ;
        RECT 97.035 136.625 97.370 137.595 ;
        RECT 98.210 136.795 98.540 137.595 ;
        RECT 99.340 136.795 99.670 137.595 ;
        RECT 98.210 136.625 100.645 136.795 ;
        RECT 101.175 136.625 101.515 137.595 ;
        RECT 104.155 137.425 106.185 137.595 ;
        RECT 96.355 136.125 96.550 136.455 ;
        RECT 96.775 136.125 97.030 136.455 ;
        RECT 96.775 135.955 96.945 136.125 ;
        RECT 97.200 135.955 97.370 136.625 ;
        RECT 98.005 136.205 98.355 136.455 ;
        RECT 98.540 135.995 98.710 136.625 ;
        RECT 98.880 136.205 99.210 136.405 ;
        RECT 99.380 136.205 99.710 136.405 ;
        RECT 99.880 136.205 100.300 136.405 ;
        RECT 100.475 136.375 100.645 136.625 ;
        RECT 100.475 136.205 101.170 136.375 ;
        RECT 96.015 135.785 96.945 135.955 ;
        RECT 96.015 135.750 96.190 135.785 ;
        RECT 95.660 135.385 96.190 135.750 ;
        RECT 97.115 135.385 97.370 135.955 ;
        RECT 98.210 135.385 98.710 135.995 ;
        RECT 99.340 135.865 100.565 136.035 ;
        RECT 101.340 136.015 101.515 136.625 ;
        RECT 103.065 137.005 103.580 137.415 ;
        RECT 103.065 136.195 103.405 137.005 ;
        RECT 104.155 136.760 104.325 137.425 ;
        RECT 104.720 137.085 105.845 137.255 ;
        RECT 103.575 136.570 104.325 136.760 ;
        RECT 104.495 136.745 105.505 136.915 ;
        RECT 103.065 136.025 104.295 136.195 ;
        RECT 99.340 135.385 99.670 135.865 ;
        RECT 100.235 135.385 100.565 135.865 ;
        RECT 101.175 135.385 101.515 136.015 ;
        RECT 103.340 135.420 103.585 136.025 ;
        RECT 104.495 135.385 104.685 136.745 ;
        RECT 104.855 136.065 105.130 136.545 ;
        RECT 104.855 135.895 105.135 136.065 ;
        RECT 105.335 135.945 105.505 136.745 ;
        RECT 105.675 135.955 105.845 137.085 ;
        RECT 106.015 136.455 106.185 137.425 ;
        RECT 106.695 136.625 107.030 137.595 ;
        RECT 106.015 136.125 106.210 136.455 ;
        RECT 106.435 136.125 106.690 136.455 ;
        RECT 106.435 135.955 106.605 136.125 ;
        RECT 106.860 135.955 107.030 136.625 ;
        RECT 104.855 135.385 105.130 135.895 ;
        RECT 105.675 135.785 106.605 135.955 ;
        RECT 105.675 135.750 105.850 135.785 ;
        RECT 105.320 135.385 105.850 135.750 ;
        RECT 106.775 135.385 107.030 135.955 ;
        RECT 107.205 136.690 107.475 137.595 ;
        RECT 108.155 136.835 108.325 137.595 ;
        RECT 110.595 137.425 112.625 137.595 ;
        RECT 107.205 135.890 107.375 136.690 ;
        RECT 107.660 136.665 108.325 136.835 ;
        RECT 109.505 137.005 110.020 137.415 ;
        RECT 107.660 136.520 107.830 136.665 ;
        RECT 107.545 136.190 107.830 136.520 ;
        RECT 107.660 135.935 107.830 136.190 ;
        RECT 108.065 136.115 108.395 136.485 ;
        RECT 109.505 136.195 109.845 137.005 ;
        RECT 110.595 136.760 110.765 137.425 ;
        RECT 111.160 137.085 112.285 137.255 ;
        RECT 110.015 136.570 110.765 136.760 ;
        RECT 110.935 136.745 111.945 136.915 ;
        RECT 109.505 136.025 110.735 136.195 ;
        RECT 107.205 135.385 107.465 135.890 ;
        RECT 107.660 135.765 108.325 135.935 ;
        RECT 108.155 135.385 108.325 135.765 ;
        RECT 109.780 135.420 110.025 136.025 ;
        RECT 110.935 135.385 111.125 136.745 ;
        RECT 111.295 136.405 111.570 136.545 ;
        RECT 111.295 136.235 111.575 136.405 ;
        RECT 111.295 135.385 111.570 136.235 ;
        RECT 111.775 135.945 111.945 136.745 ;
        RECT 112.115 135.955 112.285 137.085 ;
        RECT 112.455 136.455 112.625 137.425 ;
        RECT 113.135 136.625 113.470 137.595 ;
        RECT 112.455 136.125 112.650 136.455 ;
        RECT 112.875 136.125 113.130 136.455 ;
        RECT 112.875 135.955 113.045 136.125 ;
        RECT 113.300 135.955 113.470 136.625 ;
        RECT 114.020 136.785 114.275 137.455 ;
        RECT 114.920 137.045 115.250 137.555 ;
        RECT 114.020 136.065 114.200 136.785 ;
        RECT 114.920 136.455 115.170 137.045 ;
        RECT 115.520 136.895 115.690 137.505 ;
        RECT 116.420 137.215 116.660 137.505 ;
        RECT 117.460 137.295 118.090 137.545 ;
        RECT 117.460 137.215 117.630 137.295 ;
        RECT 119.060 137.215 119.230 137.505 ;
        RECT 120.030 137.380 120.860 137.550 ;
        RECT 116.420 137.045 117.630 137.215 ;
        RECT 114.370 136.125 115.170 136.455 ;
        RECT 112.115 135.785 113.045 135.955 ;
        RECT 112.115 135.750 112.290 135.785 ;
        RECT 111.760 135.385 112.290 135.750 ;
        RECT 113.215 135.385 113.470 135.955 ;
        RECT 113.935 135.925 114.200 136.065 ;
        RECT 113.935 135.895 114.275 135.925 ;
        RECT 114.020 135.395 114.275 135.895 ;
        RECT 114.920 135.475 115.170 136.125 ;
        RECT 115.370 136.875 115.690 136.895 ;
        RECT 115.370 136.705 117.290 136.875 ;
        RECT 115.370 135.810 115.560 136.705 ;
        RECT 117.460 136.535 117.630 137.045 ;
        RECT 117.800 136.785 118.320 137.095 ;
        RECT 115.730 136.365 117.630 136.535 ;
        RECT 115.730 136.305 116.060 136.365 ;
        RECT 116.210 136.135 116.540 136.195 ;
        RECT 115.880 135.865 116.540 136.135 ;
        RECT 115.370 135.480 115.690 135.810 ;
        RECT 116.730 135.605 116.900 136.365 ;
        RECT 117.800 136.195 117.980 136.605 ;
        RECT 117.070 136.025 117.400 136.145 ;
        RECT 118.150 136.025 118.320 136.785 ;
        RECT 117.070 135.855 118.320 136.025 ;
        RECT 118.490 136.965 119.860 137.215 ;
        RECT 118.490 136.195 118.680 136.965 ;
        RECT 119.610 136.705 119.860 136.965 ;
        RECT 118.850 136.535 119.100 136.695 ;
        RECT 120.030 136.535 120.200 137.380 ;
        RECT 121.095 137.095 121.265 137.595 ;
        RECT 120.370 136.705 120.870 137.085 ;
        RECT 121.095 136.925 121.790 137.095 ;
        RECT 118.850 136.365 120.200 136.535 ;
        RECT 119.780 136.325 120.200 136.365 ;
        RECT 118.490 135.855 118.910 136.195 ;
        RECT 119.200 135.865 119.610 136.195 ;
        RECT 116.730 135.435 117.580 135.605 ;
        RECT 118.660 135.425 118.910 135.855 ;
        RECT 119.780 135.595 119.950 136.325 ;
        RECT 120.120 135.775 120.470 136.145 ;
        RECT 120.650 135.835 120.870 136.705 ;
        RECT 121.040 136.135 121.450 136.755 ;
        RECT 121.620 135.955 121.790 136.925 ;
        RECT 121.095 135.765 121.790 135.955 ;
        RECT 119.780 135.395 120.795 135.595 ;
        RECT 121.095 135.435 121.265 135.765 ;
        RECT 121.980 135.475 122.205 137.595 ;
        RECT 122.875 137.095 123.045 137.595 ;
        RECT 122.380 136.925 123.045 137.095 ;
        RECT 122.380 135.935 122.610 136.925 ;
        RECT 123.395 136.835 123.565 137.595 ;
        RECT 122.780 136.105 123.130 136.755 ;
        RECT 123.395 136.665 124.060 136.835 ;
        RECT 124.245 136.690 124.515 137.595 ;
        RECT 123.890 136.520 124.060 136.665 ;
        RECT 123.325 136.115 123.655 136.485 ;
        RECT 123.890 136.190 124.175 136.520 ;
        RECT 123.890 135.935 124.060 136.190 ;
        RECT 122.380 135.765 123.045 135.935 ;
        RECT 122.875 135.475 123.045 135.765 ;
        RECT 123.395 135.765 124.060 135.935 ;
        RECT 124.345 135.890 124.515 136.690 ;
        RECT 123.395 135.385 123.565 135.765 ;
        RECT 124.255 135.385 124.515 135.890 ;
        RECT 16.565 134.245 16.895 134.875 ;
        RECT 16.565 133.645 16.815 134.245 ;
        RECT 17.780 134.235 18.025 134.840 ;
        RECT 17.505 134.065 18.735 134.235 ;
        RECT 16.985 133.805 17.315 134.055 ;
        RECT 16.565 132.665 16.895 133.645 ;
        RECT 17.505 133.255 17.845 134.065 ;
        RECT 18.015 133.500 18.765 133.690 ;
        RECT 17.505 132.845 18.020 133.255 ;
        RECT 18.595 132.835 18.765 133.500 ;
        RECT 18.935 133.515 19.125 134.875 ;
        RECT 19.295 134.705 19.570 134.875 ;
        RECT 19.295 134.535 19.575 134.705 ;
        RECT 19.295 133.715 19.570 134.535 ;
        RECT 19.760 134.510 20.290 134.875 ;
        RECT 20.115 134.475 20.290 134.510 ;
        RECT 19.775 133.515 19.945 134.315 ;
        RECT 18.935 133.345 19.945 133.515 ;
        RECT 20.115 134.305 21.045 134.475 ;
        RECT 21.215 134.305 21.470 134.875 ;
        RECT 22.020 134.365 22.275 134.865 ;
        RECT 20.115 133.175 20.285 134.305 ;
        RECT 20.875 134.135 21.045 134.305 ;
        RECT 19.160 133.005 20.285 133.175 ;
        RECT 20.455 133.805 20.650 134.135 ;
        RECT 20.875 133.805 21.130 134.135 ;
        RECT 20.455 132.835 20.625 133.805 ;
        RECT 21.300 133.635 21.470 134.305 ;
        RECT 21.935 134.335 22.275 134.365 ;
        RECT 21.935 134.195 22.200 134.335 ;
        RECT 18.595 132.665 20.625 132.835 ;
        RECT 21.135 132.665 21.470 133.635 ;
        RECT 22.020 133.475 22.200 134.195 ;
        RECT 22.920 134.135 23.170 134.785 ;
        RECT 22.370 133.805 23.170 134.135 ;
        RECT 22.020 132.805 22.275 133.475 ;
        RECT 22.920 133.215 23.170 133.805 ;
        RECT 23.370 134.450 23.690 134.780 ;
        RECT 24.730 134.655 25.580 134.825 ;
        RECT 23.370 133.555 23.560 134.450 ;
        RECT 23.880 134.125 24.540 134.395 ;
        RECT 24.210 134.065 24.540 134.125 ;
        RECT 23.730 133.895 24.060 133.955 ;
        RECT 24.730 133.895 24.900 134.655 ;
        RECT 26.660 134.405 26.910 134.835 ;
        RECT 25.070 134.235 26.320 134.405 ;
        RECT 25.070 134.115 25.400 134.235 ;
        RECT 23.730 133.725 25.630 133.895 ;
        RECT 23.370 133.385 25.290 133.555 ;
        RECT 23.370 133.365 23.690 133.385 ;
        RECT 22.920 132.705 23.250 133.215 ;
        RECT 23.520 132.755 23.690 133.365 ;
        RECT 25.460 133.215 25.630 133.725 ;
        RECT 25.800 133.655 25.980 134.065 ;
        RECT 26.150 133.475 26.320 134.235 ;
        RECT 24.420 133.045 25.630 133.215 ;
        RECT 25.800 133.165 26.320 133.475 ;
        RECT 26.490 134.065 26.910 134.405 ;
        RECT 27.780 134.665 28.795 134.865 ;
        RECT 27.200 134.065 27.610 134.395 ;
        RECT 26.490 133.295 26.680 134.065 ;
        RECT 27.780 133.935 27.950 134.665 ;
        RECT 29.095 134.495 29.265 134.825 ;
        RECT 28.120 134.115 28.470 134.485 ;
        RECT 27.780 133.895 28.200 133.935 ;
        RECT 26.850 133.725 28.200 133.895 ;
        RECT 26.850 133.565 27.100 133.725 ;
        RECT 27.610 133.295 27.860 133.555 ;
        RECT 26.490 133.045 27.860 133.295 ;
        RECT 24.420 132.755 24.660 133.045 ;
        RECT 25.460 132.965 25.630 133.045 ;
        RECT 25.460 132.715 26.090 132.965 ;
        RECT 27.060 132.755 27.230 133.045 ;
        RECT 28.030 132.880 28.200 133.725 ;
        RECT 28.650 133.555 28.870 134.425 ;
        RECT 29.095 134.305 29.790 134.495 ;
        RECT 28.370 133.175 28.870 133.555 ;
        RECT 29.040 133.505 29.450 134.125 ;
        RECT 29.620 133.335 29.790 134.305 ;
        RECT 29.095 133.165 29.790 133.335 ;
        RECT 28.030 132.710 28.860 132.880 ;
        RECT 29.095 132.665 29.265 133.165 ;
        RECT 29.980 132.665 30.205 134.785 ;
        RECT 30.875 134.495 31.045 134.785 ;
        RECT 30.380 134.325 31.045 134.495 ;
        RECT 31.305 134.370 31.565 134.875 ;
        RECT 32.255 134.495 32.425 134.875 ;
        RECT 30.380 133.335 30.610 134.325 ;
        RECT 30.780 133.505 31.130 134.155 ;
        RECT 31.305 133.570 31.475 134.370 ;
        RECT 31.760 134.325 32.425 134.495 ;
        RECT 31.760 134.070 31.930 134.325 ;
        RECT 33.420 134.235 33.665 134.840 ;
        RECT 31.645 133.740 31.930 134.070 ;
        RECT 32.165 133.775 32.495 134.145 ;
        RECT 33.145 134.065 34.375 134.235 ;
        RECT 31.760 133.595 31.930 133.740 ;
        RECT 30.380 133.165 31.045 133.335 ;
        RECT 30.875 132.665 31.045 133.165 ;
        RECT 31.305 132.665 31.575 133.570 ;
        RECT 31.760 133.425 32.425 133.595 ;
        RECT 32.255 132.665 32.425 133.425 ;
        RECT 33.145 133.255 33.485 134.065 ;
        RECT 33.655 133.500 34.405 133.690 ;
        RECT 33.145 132.845 33.660 133.255 ;
        RECT 34.235 132.835 34.405 133.500 ;
        RECT 34.575 133.515 34.765 134.875 ;
        RECT 34.935 134.365 35.210 134.875 ;
        RECT 35.400 134.510 35.930 134.875 ;
        RECT 35.755 134.475 35.930 134.510 ;
        RECT 34.935 134.195 35.215 134.365 ;
        RECT 34.935 133.715 35.210 134.195 ;
        RECT 35.415 133.515 35.585 134.315 ;
        RECT 34.575 133.345 35.585 133.515 ;
        RECT 35.755 134.305 36.685 134.475 ;
        RECT 36.855 134.305 37.110 134.875 ;
        RECT 35.755 133.175 35.925 134.305 ;
        RECT 36.515 134.135 36.685 134.305 ;
        RECT 34.800 133.005 35.925 133.175 ;
        RECT 36.095 133.805 36.290 134.135 ;
        RECT 36.515 133.805 36.770 134.135 ;
        RECT 36.095 132.835 36.265 133.805 ;
        RECT 36.940 133.635 37.110 134.305 ;
        RECT 34.235 132.665 36.265 132.835 ;
        RECT 36.775 132.665 37.110 133.635 ;
        RECT 37.745 134.370 38.015 134.715 ;
        RECT 38.755 134.475 38.925 134.825 ;
        RECT 39.625 134.475 39.795 134.825 ;
        RECT 37.745 133.635 37.915 134.370 ;
        RECT 38.185 134.305 39.795 134.475 ;
        RECT 42.425 134.475 42.595 134.825 ;
        RECT 43.295 134.475 43.465 134.825 ;
        RECT 38.185 134.135 38.355 134.305 ;
        RECT 38.085 133.805 38.355 134.135 ;
        RECT 38.525 133.805 38.930 134.135 ;
        RECT 38.185 133.635 38.355 133.805 ;
        RECT 39.100 133.685 39.810 134.135 ;
        RECT 39.980 133.805 40.330 134.375 ;
        RECT 41.890 133.805 42.240 134.375 ;
        RECT 42.425 134.305 44.035 134.475 ;
        RECT 44.205 134.370 44.475 134.715 ;
        RECT 43.865 134.135 44.035 134.305 ;
        RECT 37.745 132.665 38.015 133.635 ;
        RECT 38.185 133.465 38.910 133.635 ;
        RECT 39.100 133.515 39.815 133.685 ;
        RECT 38.740 133.345 38.910 133.465 ;
        RECT 40.010 133.345 40.330 133.635 ;
        RECT 38.740 133.175 40.330 133.345 ;
        RECT 41.890 133.345 42.210 133.635 ;
        RECT 42.410 133.515 43.120 134.135 ;
        RECT 43.290 133.805 43.695 134.135 ;
        RECT 43.865 133.805 44.135 134.135 ;
        RECT 43.865 133.635 44.035 133.805 ;
        RECT 44.305 133.635 44.475 134.370 ;
        RECT 43.310 133.465 44.035 133.635 ;
        RECT 43.310 133.345 43.480 133.465 ;
        RECT 41.890 133.175 43.480 133.345 ;
        RECT 38.675 132.715 40.330 133.005 ;
        RECT 41.890 132.715 43.545 133.005 ;
        RECT 44.205 132.665 44.475 133.635 ;
        RECT 44.645 134.245 44.985 134.875 ;
        RECT 45.595 134.395 45.925 134.875 ;
        RECT 46.490 134.395 46.820 134.875 ;
        RECT 44.645 133.635 44.820 134.245 ;
        RECT 45.595 134.225 46.820 134.395 ;
        RECT 47.450 134.265 47.950 134.875 ;
        RECT 44.990 133.885 45.685 134.055 ;
        RECT 45.515 133.635 45.685 133.885 ;
        RECT 45.860 133.855 46.280 134.055 ;
        RECT 46.450 133.855 46.780 134.055 ;
        RECT 46.950 133.855 47.280 134.055 ;
        RECT 47.450 133.635 47.620 134.265 ;
        RECT 48.325 134.245 48.665 134.875 ;
        RECT 49.275 134.395 49.605 134.875 ;
        RECT 50.170 134.395 50.500 134.875 ;
        RECT 48.325 134.195 48.555 134.245 ;
        RECT 49.275 134.225 50.500 134.395 ;
        RECT 51.130 134.265 51.630 134.875 ;
        RECT 52.380 134.335 52.635 134.865 ;
        RECT 47.805 133.805 48.155 134.055 ;
        RECT 48.325 133.635 48.500 134.195 ;
        RECT 48.670 133.885 49.365 134.055 ;
        RECT 49.195 133.635 49.365 133.885 ;
        RECT 49.540 133.855 49.960 134.055 ;
        RECT 50.130 133.855 50.460 134.055 ;
        RECT 50.630 133.855 50.960 134.055 ;
        RECT 51.130 133.635 51.300 134.265 ;
        RECT 51.485 133.805 51.835 134.055 ;
        RECT 44.645 132.665 44.985 133.635 ;
        RECT 45.515 133.465 47.950 133.635 ;
        RECT 46.490 132.665 46.820 133.465 ;
        RECT 47.620 132.665 47.950 133.465 ;
        RECT 48.325 132.665 48.665 133.635 ;
        RECT 49.195 133.465 51.630 133.635 ;
        RECT 50.170 132.665 50.500 133.465 ;
        RECT 51.300 132.665 51.630 133.465 ;
        RECT 52.380 133.475 52.560 134.335 ;
        RECT 53.280 134.135 53.530 134.785 ;
        RECT 52.730 133.805 53.530 134.135 ;
        RECT 52.380 133.005 52.635 133.475 ;
        RECT 52.295 132.835 52.635 133.005 ;
        RECT 52.380 132.805 52.635 132.835 ;
        RECT 53.280 133.215 53.530 133.805 ;
        RECT 53.730 134.450 54.050 134.780 ;
        RECT 55.090 134.655 55.940 134.825 ;
        RECT 53.730 133.555 53.920 134.450 ;
        RECT 54.240 134.125 54.900 134.395 ;
        RECT 54.570 134.065 54.900 134.125 ;
        RECT 54.090 133.895 54.420 133.955 ;
        RECT 55.090 133.895 55.260 134.655 ;
        RECT 57.020 134.405 57.270 134.835 ;
        RECT 55.430 134.235 56.680 134.405 ;
        RECT 55.430 134.115 55.760 134.235 ;
        RECT 54.090 133.725 55.990 133.895 ;
        RECT 53.730 133.385 55.650 133.555 ;
        RECT 53.730 133.365 54.050 133.385 ;
        RECT 53.280 132.705 53.610 133.215 ;
        RECT 53.880 132.755 54.050 133.365 ;
        RECT 55.820 133.215 55.990 133.725 ;
        RECT 56.160 133.655 56.340 134.065 ;
        RECT 56.510 133.475 56.680 134.235 ;
        RECT 54.780 133.045 55.990 133.215 ;
        RECT 56.160 133.165 56.680 133.475 ;
        RECT 56.850 134.065 57.270 134.405 ;
        RECT 58.140 134.665 59.155 134.865 ;
        RECT 57.560 134.065 57.970 134.395 ;
        RECT 56.850 133.295 57.040 134.065 ;
        RECT 58.140 133.935 58.310 134.665 ;
        RECT 59.455 134.495 59.625 134.825 ;
        RECT 58.480 134.115 58.830 134.485 ;
        RECT 58.140 133.895 58.560 133.935 ;
        RECT 57.210 133.725 58.560 133.895 ;
        RECT 57.210 133.565 57.460 133.725 ;
        RECT 57.970 133.295 58.220 133.555 ;
        RECT 56.850 133.045 58.220 133.295 ;
        RECT 54.780 132.755 55.020 133.045 ;
        RECT 55.820 132.965 55.990 133.045 ;
        RECT 55.820 132.715 56.450 132.965 ;
        RECT 57.420 132.755 57.590 133.045 ;
        RECT 58.390 132.880 58.560 133.725 ;
        RECT 59.010 133.555 59.230 134.425 ;
        RECT 59.455 134.305 60.150 134.495 ;
        RECT 58.730 133.175 59.230 133.555 ;
        RECT 59.400 133.505 59.810 134.125 ;
        RECT 59.980 133.335 60.150 134.305 ;
        RECT 59.455 133.165 60.150 133.335 ;
        RECT 58.390 132.710 59.220 132.880 ;
        RECT 59.455 132.665 59.625 133.165 ;
        RECT 60.340 132.665 60.565 134.785 ;
        RECT 61.235 134.495 61.405 134.785 ;
        RECT 60.740 134.325 61.405 134.495 ;
        RECT 60.740 133.335 60.970 134.325 ;
        RECT 63.505 134.245 63.845 134.875 ;
        RECT 64.455 134.395 64.785 134.875 ;
        RECT 65.350 134.395 65.680 134.875 ;
        RECT 61.140 133.505 61.490 134.155 ;
        RECT 63.505 133.635 63.680 134.245 ;
        RECT 64.455 134.225 65.680 134.395 ;
        RECT 66.310 134.265 66.810 134.875 ;
        RECT 79.685 134.475 79.855 134.825 ;
        RECT 80.555 134.475 80.725 134.825 ;
        RECT 63.850 133.885 64.545 134.055 ;
        RECT 64.375 133.635 64.545 133.885 ;
        RECT 64.720 133.855 65.140 134.055 ;
        RECT 65.310 133.855 65.640 134.055 ;
        RECT 65.810 133.855 66.140 134.055 ;
        RECT 66.310 133.635 66.480 134.265 ;
        RECT 66.665 133.805 67.015 134.055 ;
        RECT 79.150 133.805 79.500 134.375 ;
        RECT 79.685 134.305 81.295 134.475 ;
        RECT 81.465 134.370 81.735 134.715 ;
        RECT 81.125 134.135 81.295 134.305 ;
        RECT 60.740 133.165 61.405 133.335 ;
        RECT 61.235 132.665 61.405 133.165 ;
        RECT 63.505 132.665 63.845 133.635 ;
        RECT 64.375 133.465 66.810 133.635 ;
        RECT 65.350 132.665 65.680 133.465 ;
        RECT 66.480 132.665 66.810 133.465 ;
        RECT 79.150 133.345 79.470 133.635 ;
        RECT 79.670 133.515 80.380 134.135 ;
        RECT 80.550 133.805 80.955 134.135 ;
        RECT 81.125 133.805 81.395 134.135 ;
        RECT 81.125 133.635 81.295 133.805 ;
        RECT 81.565 133.635 81.735 134.370 ;
        RECT 80.570 133.465 81.295 133.635 ;
        RECT 80.570 133.345 80.740 133.465 ;
        RECT 79.150 133.175 80.740 133.345 ;
        RECT 79.150 132.715 80.805 133.005 ;
        RECT 81.465 132.665 81.735 133.635 ;
        RECT 87.865 134.245 88.195 134.875 ;
        RECT 89.640 134.705 89.895 134.865 ;
        RECT 89.555 134.535 89.895 134.705 ;
        RECT 89.640 134.335 89.895 134.535 ;
        RECT 87.865 133.645 88.115 134.245 ;
        RECT 88.285 133.805 88.615 134.055 ;
        RECT 87.865 132.665 88.195 133.645 ;
        RECT 89.640 133.475 89.820 134.335 ;
        RECT 90.540 134.135 90.790 134.785 ;
        RECT 89.990 133.805 90.790 134.135 ;
        RECT 89.640 132.805 89.895 133.475 ;
        RECT 90.540 133.215 90.790 133.805 ;
        RECT 90.990 134.450 91.310 134.780 ;
        RECT 92.350 134.655 93.200 134.825 ;
        RECT 90.990 133.555 91.180 134.450 ;
        RECT 91.500 134.125 92.160 134.395 ;
        RECT 91.830 134.065 92.160 134.125 ;
        RECT 91.350 133.895 91.680 133.955 ;
        RECT 92.350 133.895 92.520 134.655 ;
        RECT 94.280 134.405 94.530 134.835 ;
        RECT 92.690 134.235 93.940 134.405 ;
        RECT 92.690 134.115 93.020 134.235 ;
        RECT 91.350 133.725 93.250 133.895 ;
        RECT 90.990 133.385 92.910 133.555 ;
        RECT 90.990 133.365 91.310 133.385 ;
        RECT 90.540 132.705 90.870 133.215 ;
        RECT 91.140 132.755 91.310 133.365 ;
        RECT 93.080 133.215 93.250 133.725 ;
        RECT 93.420 133.655 93.600 134.065 ;
        RECT 93.770 133.475 93.940 134.235 ;
        RECT 92.040 133.045 93.250 133.215 ;
        RECT 93.420 133.165 93.940 133.475 ;
        RECT 94.110 134.065 94.530 134.405 ;
        RECT 95.400 134.665 96.415 134.865 ;
        RECT 94.820 134.065 95.230 134.395 ;
        RECT 94.110 133.295 94.300 134.065 ;
        RECT 95.400 133.935 95.570 134.665 ;
        RECT 96.715 134.495 96.885 134.825 ;
        RECT 95.740 134.115 96.090 134.485 ;
        RECT 95.400 133.895 95.820 133.935 ;
        RECT 94.470 133.725 95.820 133.895 ;
        RECT 94.470 133.565 94.720 133.725 ;
        RECT 95.230 133.295 95.480 133.555 ;
        RECT 94.110 133.045 95.480 133.295 ;
        RECT 92.040 132.755 92.280 133.045 ;
        RECT 93.080 132.965 93.250 133.045 ;
        RECT 93.080 132.715 93.710 132.965 ;
        RECT 94.680 132.755 94.850 133.045 ;
        RECT 95.650 132.880 95.820 133.725 ;
        RECT 96.270 133.555 96.490 134.425 ;
        RECT 96.715 134.305 97.410 134.495 ;
        RECT 95.990 133.175 96.490 133.555 ;
        RECT 96.660 133.505 97.070 134.125 ;
        RECT 97.240 133.335 97.410 134.305 ;
        RECT 96.715 133.165 97.410 133.335 ;
        RECT 95.650 132.710 96.480 132.880 ;
        RECT 96.715 132.665 96.885 133.165 ;
        RECT 97.600 132.665 97.825 134.785 ;
        RECT 98.495 134.495 98.665 134.785 ;
        RECT 98.000 134.325 98.665 134.495 ;
        RECT 99.300 134.335 99.555 134.865 ;
        RECT 98.000 133.335 98.230 134.325 ;
        RECT 98.400 133.505 98.750 134.155 ;
        RECT 99.300 133.475 99.480 134.335 ;
        RECT 100.200 134.135 100.450 134.785 ;
        RECT 99.650 133.805 100.450 134.135 ;
        RECT 98.000 133.165 98.665 133.335 ;
        RECT 98.495 132.665 98.665 133.165 ;
        RECT 99.300 133.005 99.555 133.475 ;
        RECT 99.215 132.835 99.555 133.005 ;
        RECT 99.300 132.805 99.555 132.835 ;
        RECT 100.200 133.215 100.450 133.805 ;
        RECT 100.650 134.450 100.970 134.780 ;
        RECT 102.010 134.655 102.860 134.825 ;
        RECT 100.650 133.555 100.840 134.450 ;
        RECT 101.160 134.125 101.820 134.395 ;
        RECT 101.490 134.065 101.820 134.125 ;
        RECT 101.010 133.895 101.340 133.955 ;
        RECT 102.010 133.895 102.180 134.655 ;
        RECT 103.940 134.405 104.190 134.835 ;
        RECT 102.350 134.235 103.600 134.405 ;
        RECT 102.350 134.115 102.680 134.235 ;
        RECT 101.010 133.725 102.910 133.895 ;
        RECT 100.650 133.385 102.570 133.555 ;
        RECT 100.650 133.365 100.970 133.385 ;
        RECT 100.200 132.705 100.530 133.215 ;
        RECT 100.800 132.755 100.970 133.365 ;
        RECT 102.740 133.215 102.910 133.725 ;
        RECT 103.080 133.655 103.260 134.065 ;
        RECT 103.430 133.475 103.600 134.235 ;
        RECT 101.700 133.045 102.910 133.215 ;
        RECT 103.080 133.165 103.600 133.475 ;
        RECT 103.770 134.065 104.190 134.405 ;
        RECT 105.060 134.665 106.075 134.865 ;
        RECT 104.480 134.065 104.890 134.395 ;
        RECT 103.770 133.295 103.960 134.065 ;
        RECT 105.060 133.935 105.230 134.665 ;
        RECT 106.375 134.495 106.545 134.825 ;
        RECT 105.400 134.115 105.750 134.485 ;
        RECT 105.060 133.895 105.480 133.935 ;
        RECT 104.130 133.725 105.480 133.895 ;
        RECT 104.130 133.565 104.380 133.725 ;
        RECT 104.890 133.295 105.140 133.555 ;
        RECT 103.770 133.045 105.140 133.295 ;
        RECT 101.700 132.755 101.940 133.045 ;
        RECT 102.740 132.965 102.910 133.045 ;
        RECT 102.740 132.715 103.370 132.965 ;
        RECT 104.340 132.755 104.510 133.045 ;
        RECT 105.310 132.880 105.480 133.725 ;
        RECT 105.930 133.555 106.150 134.425 ;
        RECT 106.375 134.305 107.070 134.495 ;
        RECT 105.650 133.175 106.150 133.555 ;
        RECT 106.320 133.505 106.730 134.125 ;
        RECT 106.900 133.335 107.070 134.305 ;
        RECT 106.375 133.165 107.070 133.335 ;
        RECT 105.310 132.710 106.140 132.880 ;
        RECT 106.375 132.665 106.545 133.165 ;
        RECT 107.260 132.665 107.485 134.785 ;
        RECT 108.155 134.495 108.325 134.785 ;
        RECT 107.660 134.325 108.325 134.495 ;
        RECT 109.125 134.475 109.295 134.825 ;
        RECT 109.995 134.475 110.165 134.825 ;
        RECT 107.660 133.335 107.890 134.325 ;
        RECT 108.060 133.505 108.410 134.155 ;
        RECT 108.590 133.805 108.940 134.375 ;
        RECT 109.125 134.305 110.735 134.475 ;
        RECT 110.905 134.370 111.175 134.715 ;
        RECT 110.565 134.135 110.735 134.305 ;
        RECT 108.590 133.345 108.910 133.635 ;
        RECT 109.110 133.515 109.820 134.135 ;
        RECT 109.990 133.805 110.395 134.135 ;
        RECT 110.565 133.805 110.835 134.135 ;
        RECT 110.565 133.635 110.735 133.805 ;
        RECT 111.005 133.635 111.175 134.370 ;
        RECT 119.255 134.495 119.425 134.875 ;
        RECT 119.255 134.325 119.920 134.495 ;
        RECT 120.115 134.370 120.375 134.875 ;
        RECT 119.185 133.775 119.515 134.145 ;
        RECT 119.750 134.070 119.920 134.325 ;
        RECT 110.010 133.465 110.735 133.635 ;
        RECT 110.010 133.345 110.180 133.465 ;
        RECT 107.660 133.165 108.325 133.335 ;
        RECT 108.590 133.175 110.180 133.345 ;
        RECT 108.155 132.665 108.325 133.165 ;
        RECT 108.590 132.715 110.245 133.005 ;
        RECT 110.905 132.665 111.175 133.635 ;
        RECT 119.750 133.740 120.035 134.070 ;
        RECT 119.750 133.595 119.920 133.740 ;
        RECT 119.255 133.425 119.920 133.595 ;
        RECT 120.205 133.570 120.375 134.370 ;
        RECT 119.255 132.665 119.425 133.425 ;
        RECT 120.105 132.665 120.375 133.570 ;
        RECT 21.355 131.985 23.385 132.155 ;
        RECT 20.265 131.565 20.780 131.975 ;
        RECT 20.265 130.755 20.605 131.565 ;
        RECT 21.355 131.320 21.525 131.985 ;
        RECT 21.920 131.645 23.045 131.815 ;
        RECT 20.775 131.130 21.525 131.320 ;
        RECT 21.695 131.305 22.705 131.475 ;
        RECT 20.265 130.585 21.495 130.755 ;
        RECT 20.540 129.980 20.785 130.585 ;
        RECT 21.695 129.945 21.885 131.305 ;
        RECT 22.055 130.625 22.330 131.105 ;
        RECT 22.055 130.455 22.335 130.625 ;
        RECT 22.535 130.505 22.705 131.305 ;
        RECT 22.875 130.515 23.045 131.645 ;
        RECT 23.215 131.015 23.385 131.985 ;
        RECT 23.895 131.185 24.230 132.155 ;
        RECT 30.760 131.985 31.015 132.015 ;
        RECT 30.675 131.815 31.015 131.985 ;
        RECT 23.215 130.685 23.410 131.015 ;
        RECT 23.635 130.685 23.890 131.015 ;
        RECT 23.635 130.515 23.805 130.685 ;
        RECT 24.060 130.515 24.230 131.185 ;
        RECT 22.055 129.945 22.330 130.455 ;
        RECT 22.875 130.345 23.805 130.515 ;
        RECT 22.875 130.310 23.050 130.345 ;
        RECT 22.520 129.945 23.050 130.310 ;
        RECT 23.975 129.945 24.230 130.515 ;
        RECT 30.760 131.345 31.015 131.815 ;
        RECT 31.660 131.605 31.990 132.115 ;
        RECT 30.760 130.485 30.940 131.345 ;
        RECT 31.660 131.015 31.910 131.605 ;
        RECT 32.260 131.455 32.430 132.065 ;
        RECT 33.160 131.775 33.400 132.065 ;
        RECT 34.200 131.855 34.830 132.105 ;
        RECT 34.200 131.775 34.370 131.855 ;
        RECT 35.800 131.775 35.970 132.065 ;
        RECT 36.770 131.940 37.600 132.110 ;
        RECT 33.160 131.605 34.370 131.775 ;
        RECT 31.110 130.685 31.910 131.015 ;
        RECT 30.760 129.955 31.015 130.485 ;
        RECT 31.660 130.035 31.910 130.685 ;
        RECT 32.110 131.435 32.430 131.455 ;
        RECT 32.110 131.265 34.030 131.435 ;
        RECT 32.110 130.370 32.300 131.265 ;
        RECT 34.200 131.095 34.370 131.605 ;
        RECT 34.540 131.345 35.060 131.655 ;
        RECT 32.470 130.925 34.370 131.095 ;
        RECT 32.470 130.865 32.800 130.925 ;
        RECT 32.950 130.695 33.280 130.755 ;
        RECT 32.620 130.425 33.280 130.695 ;
        RECT 32.110 130.040 32.430 130.370 ;
        RECT 33.470 130.165 33.640 130.925 ;
        RECT 34.540 130.755 34.720 131.165 ;
        RECT 33.810 130.585 34.140 130.705 ;
        RECT 34.890 130.585 35.060 131.345 ;
        RECT 33.810 130.415 35.060 130.585 ;
        RECT 35.230 131.525 36.600 131.775 ;
        RECT 35.230 130.755 35.420 131.525 ;
        RECT 36.350 131.265 36.600 131.525 ;
        RECT 35.590 131.095 35.840 131.255 ;
        RECT 36.770 131.095 36.940 131.940 ;
        RECT 37.835 131.655 38.005 132.155 ;
        RECT 37.110 131.265 37.610 131.645 ;
        RECT 37.835 131.485 38.530 131.655 ;
        RECT 35.590 130.925 36.940 131.095 ;
        RECT 36.520 130.885 36.940 130.925 ;
        RECT 35.230 130.415 35.650 130.755 ;
        RECT 35.940 130.425 36.350 130.755 ;
        RECT 33.470 129.995 34.320 130.165 ;
        RECT 35.400 129.985 35.650 130.415 ;
        RECT 36.520 130.155 36.690 130.885 ;
        RECT 36.860 130.335 37.210 130.705 ;
        RECT 37.390 130.395 37.610 131.265 ;
        RECT 37.780 130.695 38.190 131.315 ;
        RECT 38.360 130.515 38.530 131.485 ;
        RECT 37.835 130.325 38.530 130.515 ;
        RECT 36.520 129.955 37.535 130.155 ;
        RECT 37.835 129.995 38.005 130.325 ;
        RECT 38.720 130.035 38.945 132.155 ;
        RECT 39.615 131.655 39.785 132.155 ;
        RECT 39.120 131.485 39.785 131.655 ;
        RECT 39.120 130.495 39.350 131.485 ;
        RECT 39.520 130.665 39.870 131.315 ;
        RECT 40.045 131.250 40.315 132.155 ;
        RECT 40.995 131.395 41.165 132.155 ;
        RECT 39.120 130.325 39.785 130.495 ;
        RECT 39.615 130.035 39.785 130.325 ;
        RECT 40.045 130.450 40.215 131.250 ;
        RECT 40.500 131.225 41.165 131.395 ;
        RECT 43.455 131.435 43.755 131.985 ;
        RECT 44.475 131.605 44.935 132.155 ;
        RECT 40.500 131.080 40.670 131.225 ;
        RECT 40.385 130.750 40.670 131.080 ;
        RECT 40.500 130.495 40.670 130.750 ;
        RECT 40.905 130.675 41.235 131.045 ;
        RECT 42.820 131.015 43.085 131.375 ;
        RECT 43.455 131.265 44.395 131.435 ;
        RECT 44.225 131.015 44.395 131.265 ;
        RECT 42.820 130.765 43.495 131.015 ;
        RECT 43.715 130.765 44.055 131.015 ;
        RECT 44.225 130.685 44.515 131.015 ;
        RECT 44.225 130.595 44.395 130.685 ;
        RECT 40.045 129.945 40.305 130.450 ;
        RECT 40.500 130.325 41.165 130.495 ;
        RECT 40.995 129.945 41.165 130.325 ;
        RECT 43.005 130.405 44.395 130.595 ;
        RECT 43.005 130.045 43.335 130.405 ;
        RECT 44.685 130.235 44.935 131.605 ;
        RECT 45.755 131.435 46.055 131.985 ;
        RECT 46.775 131.605 47.235 132.155 ;
        RECT 66.435 131.985 68.465 132.155 ;
        RECT 45.120 131.015 45.385 131.375 ;
        RECT 45.755 131.265 46.695 131.435 ;
        RECT 46.525 131.015 46.695 131.265 ;
        RECT 45.120 130.765 45.795 131.015 ;
        RECT 46.015 130.765 46.355 131.015 ;
        RECT 46.525 130.685 46.815 131.015 ;
        RECT 46.525 130.595 46.695 130.685 ;
        RECT 44.375 129.945 44.935 130.235 ;
        RECT 45.305 130.405 46.695 130.595 ;
        RECT 45.305 130.045 45.635 130.405 ;
        RECT 46.985 130.235 47.235 131.605 ;
        RECT 65.345 131.565 65.860 131.975 ;
        RECT 65.345 130.755 65.685 131.565 ;
        RECT 66.435 131.320 66.605 131.985 ;
        RECT 67.000 131.645 68.125 131.815 ;
        RECT 65.855 131.130 66.605 131.320 ;
        RECT 66.775 131.305 67.785 131.475 ;
        RECT 65.345 130.585 66.575 130.755 ;
        RECT 46.675 129.945 47.235 130.235 ;
        RECT 65.620 129.980 65.865 130.585 ;
        RECT 66.775 129.945 66.965 131.305 ;
        RECT 67.135 130.625 67.410 131.105 ;
        RECT 67.135 130.455 67.415 130.625 ;
        RECT 67.615 130.505 67.785 131.305 ;
        RECT 67.955 130.515 68.125 131.645 ;
        RECT 68.295 131.015 68.465 131.985 ;
        RECT 68.975 131.185 69.310 132.155 ;
        RECT 70.455 131.720 70.640 132.125 ;
        RECT 68.295 130.685 68.490 131.015 ;
        RECT 68.715 130.685 68.970 131.015 ;
        RECT 68.715 130.515 68.885 130.685 ;
        RECT 69.140 130.515 69.310 131.185 ;
        RECT 67.135 129.945 67.410 130.455 ;
        RECT 67.955 130.345 68.885 130.515 ;
        RECT 67.955 130.310 68.130 130.345 ;
        RECT 67.600 129.945 68.130 130.310 ;
        RECT 69.055 129.945 69.310 130.515 ;
        RECT 69.975 131.545 70.640 131.720 ;
        RECT 69.975 130.515 70.315 131.545 ;
        RECT 71.345 131.355 71.615 132.125 ;
        RECT 70.485 131.185 71.615 131.355 ;
        RECT 70.485 130.685 70.735 131.185 ;
        RECT 69.975 130.345 70.660 130.515 ;
        RECT 70.915 130.435 71.275 131.015 ;
        RECT 70.455 129.945 70.660 130.345 ;
        RECT 71.445 130.275 71.615 131.185 ;
        RECT 71.355 129.945 71.615 130.275 ;
        RECT 71.785 131.605 72.245 132.155 ;
        RECT 71.785 130.235 72.035 131.605 ;
        RECT 72.965 131.435 73.265 131.985 ;
        RECT 72.325 131.265 73.265 131.435 ;
        RECT 72.325 131.015 72.495 131.265 ;
        RECT 73.635 131.015 73.900 131.375 ;
        RECT 72.205 130.685 72.495 131.015 ;
        RECT 72.665 130.765 73.005 131.015 ;
        RECT 73.225 130.765 73.900 131.015 ;
        RECT 74.085 131.355 74.355 132.125 ;
        RECT 75.060 131.720 75.245 132.125 ;
        RECT 75.060 131.545 75.725 131.720 ;
        RECT 74.085 131.185 75.215 131.355 ;
        RECT 72.325 130.595 72.495 130.685 ;
        RECT 72.325 130.405 73.715 130.595 ;
        RECT 71.785 129.945 72.345 130.235 ;
        RECT 73.385 130.045 73.715 130.405 ;
        RECT 74.085 130.275 74.255 131.185 ;
        RECT 74.425 130.435 74.785 131.015 ;
        RECT 74.965 130.685 75.215 131.185 ;
        RECT 75.385 130.515 75.725 131.545 ;
        RECT 75.040 130.345 75.725 130.515 ;
        RECT 78.685 131.605 79.145 132.155 ;
        RECT 74.085 129.945 74.345 130.275 ;
        RECT 75.040 129.945 75.245 130.345 ;
        RECT 78.685 130.235 78.935 131.605 ;
        RECT 79.865 131.435 80.165 131.985 ;
        RECT 79.225 131.265 80.165 131.435 ;
        RECT 79.225 131.015 79.395 131.265 ;
        RECT 80.535 131.015 80.800 131.375 ;
        RECT 88.325 131.175 88.655 132.155 ;
        RECT 90.355 131.985 92.385 132.155 ;
        RECT 79.105 130.685 79.395 131.015 ;
        RECT 79.565 130.765 79.905 131.015 ;
        RECT 80.125 130.765 80.800 131.015 ;
        RECT 87.905 130.765 88.235 131.015 ;
        RECT 79.225 130.595 79.395 130.685 ;
        RECT 79.225 130.405 80.615 130.595 ;
        RECT 88.405 130.575 88.655 131.175 ;
        RECT 89.265 131.565 89.780 131.975 ;
        RECT 89.265 130.755 89.605 131.565 ;
        RECT 90.355 131.320 90.525 131.985 ;
        RECT 90.920 131.645 92.045 131.815 ;
        RECT 89.775 131.130 90.525 131.320 ;
        RECT 90.695 131.305 91.705 131.475 ;
        RECT 89.265 130.585 90.495 130.755 ;
        RECT 78.685 129.945 79.245 130.235 ;
        RECT 80.285 130.045 80.615 130.405 ;
        RECT 88.325 129.945 88.655 130.575 ;
        RECT 89.540 129.980 89.785 130.585 ;
        RECT 90.695 129.945 90.885 131.305 ;
        RECT 91.055 130.285 91.330 131.105 ;
        RECT 91.535 130.505 91.705 131.305 ;
        RECT 91.875 130.515 92.045 131.645 ;
        RECT 92.215 131.015 92.385 131.985 ;
        RECT 92.895 131.185 93.230 132.155 ;
        RECT 93.955 131.395 94.125 132.155 ;
        RECT 93.955 131.225 94.620 131.395 ;
        RECT 94.805 131.250 95.075 132.155 ;
        RECT 92.215 130.685 92.410 131.015 ;
        RECT 92.635 130.685 92.890 131.015 ;
        RECT 92.635 130.515 92.805 130.685 ;
        RECT 93.060 130.515 93.230 131.185 ;
        RECT 94.450 131.080 94.620 131.225 ;
        RECT 93.885 130.675 94.215 131.045 ;
        RECT 94.450 130.750 94.735 131.080 ;
        RECT 91.875 130.345 92.805 130.515 ;
        RECT 91.875 130.310 92.050 130.345 ;
        RECT 91.055 130.115 91.335 130.285 ;
        RECT 91.055 129.945 91.330 130.115 ;
        RECT 91.520 129.945 92.050 130.310 ;
        RECT 92.975 129.945 93.230 130.515 ;
        RECT 94.450 130.495 94.620 130.750 ;
        RECT 93.955 130.325 94.620 130.495 ;
        RECT 94.905 130.450 95.075 131.250 ;
        RECT 95.335 131.395 95.505 132.155 ;
        RECT 95.335 131.225 96.000 131.395 ;
        RECT 96.185 131.250 96.455 132.155 ;
        RECT 95.830 131.080 96.000 131.225 ;
        RECT 95.265 130.675 95.595 131.045 ;
        RECT 95.830 130.750 96.115 131.080 ;
        RECT 95.830 130.495 96.000 130.750 ;
        RECT 93.955 129.945 94.125 130.325 ;
        RECT 94.815 129.945 95.075 130.450 ;
        RECT 95.335 130.325 96.000 130.495 ;
        RECT 96.285 130.450 96.455 131.250 ;
        RECT 95.335 129.945 95.505 130.325 ;
        RECT 96.195 129.945 96.455 130.450 ;
        RECT 98.005 131.185 98.275 132.155 ;
        RECT 98.935 131.815 100.590 132.105 ;
        RECT 103.990 131.815 105.645 132.105 ;
        RECT 99.000 131.475 100.590 131.645 ;
        RECT 99.000 131.355 99.170 131.475 ;
        RECT 98.445 131.185 99.170 131.355 ;
        RECT 98.005 130.450 98.175 131.185 ;
        RECT 98.445 131.015 98.615 131.185 ;
        RECT 99.360 131.135 100.075 131.305 ;
        RECT 100.270 131.185 100.590 131.475 ;
        RECT 103.990 131.475 105.580 131.645 ;
        RECT 103.990 131.185 104.310 131.475 ;
        RECT 105.410 131.355 105.580 131.475 ;
        RECT 104.505 131.135 105.220 131.305 ;
        RECT 105.410 131.185 106.135 131.355 ;
        RECT 106.305 131.185 106.575 132.155 ;
        RECT 98.345 130.685 98.615 131.015 ;
        RECT 98.785 130.685 99.190 131.015 ;
        RECT 99.360 130.685 100.070 131.135 ;
        RECT 98.445 130.515 98.615 130.685 ;
        RECT 98.005 130.105 98.275 130.450 ;
        RECT 98.445 130.345 100.055 130.515 ;
        RECT 100.240 130.445 100.590 131.015 ;
        RECT 103.990 130.445 104.340 131.015 ;
        RECT 104.510 130.685 105.220 131.135 ;
        RECT 105.965 131.015 106.135 131.185 ;
        RECT 105.390 130.685 105.795 131.015 ;
        RECT 105.965 130.685 106.235 131.015 ;
        RECT 105.965 130.515 106.135 130.685 ;
        RECT 99.015 129.995 99.185 130.345 ;
        RECT 99.885 129.995 100.055 130.345 ;
        RECT 104.525 130.345 106.135 130.515 ;
        RECT 106.405 130.450 106.575 131.185 ;
        RECT 104.525 129.995 104.695 130.345 ;
        RECT 105.395 129.995 105.565 130.345 ;
        RECT 106.305 130.105 106.575 130.450 ;
        RECT 110.425 131.605 110.885 132.155 ;
        RECT 110.425 130.235 110.675 131.605 ;
        RECT 111.605 131.435 111.905 131.985 ;
        RECT 110.965 131.265 111.905 131.435 ;
        RECT 110.965 131.015 111.135 131.265 ;
        RECT 112.275 131.015 112.540 131.375 ;
        RECT 110.845 130.685 111.135 131.015 ;
        RECT 111.305 130.765 111.645 131.015 ;
        RECT 111.865 130.765 112.540 131.015 ;
        RECT 110.965 130.595 111.135 130.685 ;
        RECT 110.965 130.405 112.355 130.595 ;
        RECT 110.425 129.945 110.985 130.235 ;
        RECT 112.025 130.045 112.355 130.405 ;
        RECT 17.420 129.265 17.675 129.425 ;
        RECT 17.335 129.095 17.675 129.265 ;
        RECT 17.420 128.895 17.675 129.095 ;
        RECT 17.420 128.035 17.600 128.895 ;
        RECT 18.320 128.695 18.570 129.345 ;
        RECT 17.770 128.365 18.570 128.695 ;
        RECT 17.420 127.365 17.675 128.035 ;
        RECT 18.320 127.775 18.570 128.365 ;
        RECT 18.770 129.010 19.090 129.340 ;
        RECT 20.130 129.215 20.980 129.385 ;
        RECT 18.770 128.115 18.960 129.010 ;
        RECT 19.280 128.685 19.940 128.955 ;
        RECT 19.610 128.625 19.940 128.685 ;
        RECT 19.130 128.455 19.460 128.515 ;
        RECT 20.130 128.455 20.300 129.215 ;
        RECT 22.060 128.965 22.310 129.395 ;
        RECT 20.470 128.795 21.720 128.965 ;
        RECT 20.470 128.675 20.800 128.795 ;
        RECT 19.130 128.285 21.030 128.455 ;
        RECT 18.770 127.945 20.690 128.115 ;
        RECT 18.770 127.925 19.090 127.945 ;
        RECT 18.320 127.265 18.650 127.775 ;
        RECT 18.920 127.315 19.090 127.925 ;
        RECT 20.860 127.775 21.030 128.285 ;
        RECT 21.200 128.215 21.380 128.625 ;
        RECT 21.550 128.035 21.720 128.795 ;
        RECT 19.820 127.605 21.030 127.775 ;
        RECT 21.200 127.725 21.720 128.035 ;
        RECT 21.890 128.625 22.310 128.965 ;
        RECT 23.180 129.225 24.195 129.425 ;
        RECT 22.600 128.625 23.010 128.955 ;
        RECT 21.890 127.855 22.080 128.625 ;
        RECT 23.180 128.495 23.350 129.225 ;
        RECT 24.495 129.055 24.665 129.385 ;
        RECT 23.520 128.675 23.870 129.045 ;
        RECT 23.180 128.455 23.600 128.495 ;
        RECT 22.250 128.285 23.600 128.455 ;
        RECT 22.250 128.125 22.500 128.285 ;
        RECT 23.010 127.855 23.260 128.115 ;
        RECT 21.890 127.605 23.260 127.855 ;
        RECT 19.820 127.315 20.060 127.605 ;
        RECT 20.860 127.525 21.030 127.605 ;
        RECT 20.860 127.275 21.490 127.525 ;
        RECT 22.460 127.315 22.630 127.605 ;
        RECT 23.430 127.440 23.600 128.285 ;
        RECT 24.050 128.115 24.270 128.985 ;
        RECT 24.495 128.865 25.190 129.055 ;
        RECT 23.770 127.735 24.270 128.115 ;
        RECT 24.440 128.065 24.850 128.685 ;
        RECT 25.020 127.895 25.190 128.865 ;
        RECT 24.495 127.725 25.190 127.895 ;
        RECT 23.430 127.270 24.260 127.440 ;
        RECT 24.495 127.225 24.665 127.725 ;
        RECT 25.380 127.225 25.605 129.345 ;
        RECT 26.275 129.055 26.445 129.345 ;
        RECT 25.780 128.885 26.445 129.055 ;
        RECT 25.780 127.895 26.010 128.885 ;
        RECT 34.045 128.805 34.375 129.435 ;
        RECT 26.180 128.065 26.530 128.715 ;
        RECT 33.625 128.365 33.955 128.615 ;
        RECT 34.125 128.205 34.375 128.805 ;
        RECT 35.185 128.975 35.515 129.335 ;
        RECT 36.555 129.145 37.115 129.435 ;
        RECT 35.185 128.785 36.575 128.975 ;
        RECT 36.405 128.695 36.575 128.785 ;
        RECT 25.780 127.725 26.445 127.895 ;
        RECT 26.275 127.225 26.445 127.725 ;
        RECT 34.045 127.225 34.375 128.205 ;
        RECT 35.000 128.365 35.675 128.615 ;
        RECT 35.895 128.365 36.235 128.615 ;
        RECT 36.405 128.365 36.695 128.695 ;
        RECT 35.000 128.005 35.265 128.365 ;
        RECT 36.405 128.115 36.575 128.365 ;
        RECT 35.635 127.945 36.575 128.115 ;
        RECT 35.635 127.395 35.935 127.945 ;
        RECT 36.865 127.775 37.115 129.145 ;
        RECT 46.685 128.975 47.015 129.335 ;
        RECT 48.055 129.145 48.615 129.435 ;
        RECT 46.685 128.785 48.075 128.975 ;
        RECT 47.905 128.695 48.075 128.785 ;
        RECT 46.500 128.365 47.175 128.615 ;
        RECT 47.395 128.365 47.735 128.615 ;
        RECT 47.905 128.365 48.195 128.695 ;
        RECT 46.500 128.005 46.765 128.365 ;
        RECT 47.905 128.115 48.075 128.365 ;
        RECT 36.655 127.225 37.115 127.775 ;
        RECT 47.135 127.945 48.075 128.115 ;
        RECT 47.135 127.395 47.435 127.945 ;
        RECT 48.365 127.775 48.615 129.145 ;
        RECT 55.040 128.795 55.285 129.400 ;
        RECT 48.155 127.225 48.615 127.775 ;
        RECT 54.765 128.625 55.995 128.795 ;
        RECT 54.765 127.815 55.105 128.625 ;
        RECT 55.275 128.060 56.025 128.250 ;
        RECT 54.765 127.405 55.280 127.815 ;
        RECT 55.855 127.395 56.025 128.060 ;
        RECT 56.195 128.075 56.385 129.435 ;
        RECT 56.555 129.265 56.830 129.435 ;
        RECT 56.555 129.095 56.835 129.265 ;
        RECT 56.555 128.275 56.830 129.095 ;
        RECT 57.020 129.070 57.550 129.435 ;
        RECT 57.375 129.035 57.550 129.070 ;
        RECT 57.035 128.075 57.205 128.875 ;
        RECT 56.195 127.905 57.205 128.075 ;
        RECT 57.375 128.865 58.305 129.035 ;
        RECT 58.475 128.865 58.730 129.435 ;
        RECT 58.995 129.055 59.165 129.435 ;
        RECT 58.995 128.885 59.660 129.055 ;
        RECT 59.855 128.930 60.115 129.435 ;
        RECT 65.260 129.265 65.515 129.425 ;
        RECT 65.175 129.095 65.515 129.265 ;
        RECT 57.375 127.735 57.545 128.865 ;
        RECT 58.135 128.695 58.305 128.865 ;
        RECT 56.420 127.565 57.545 127.735 ;
        RECT 57.715 128.365 57.910 128.695 ;
        RECT 58.135 128.365 58.390 128.695 ;
        RECT 57.715 127.395 57.885 128.365 ;
        RECT 58.560 128.195 58.730 128.865 ;
        RECT 58.925 128.335 59.255 128.705 ;
        RECT 59.490 128.630 59.660 128.885 ;
        RECT 55.855 127.225 57.885 127.395 ;
        RECT 58.395 127.225 58.730 128.195 ;
        RECT 59.490 128.300 59.775 128.630 ;
        RECT 59.490 128.155 59.660 128.300 ;
        RECT 58.995 127.985 59.660 128.155 ;
        RECT 59.945 128.130 60.115 128.930 ;
        RECT 58.995 127.225 59.165 127.985 ;
        RECT 59.845 127.225 60.115 128.130 ;
        RECT 65.260 128.895 65.515 129.095 ;
        RECT 65.260 128.035 65.440 128.895 ;
        RECT 66.160 128.695 66.410 129.345 ;
        RECT 65.610 128.365 66.410 128.695 ;
        RECT 65.260 127.365 65.515 128.035 ;
        RECT 66.160 127.775 66.410 128.365 ;
        RECT 66.610 129.010 66.930 129.340 ;
        RECT 67.970 129.215 68.820 129.385 ;
        RECT 66.610 128.115 66.800 129.010 ;
        RECT 67.120 128.685 67.780 128.955 ;
        RECT 67.450 128.625 67.780 128.685 ;
        RECT 66.970 128.455 67.300 128.515 ;
        RECT 67.970 128.455 68.140 129.215 ;
        RECT 69.900 128.965 70.150 129.395 ;
        RECT 68.310 128.795 69.560 128.965 ;
        RECT 68.310 128.675 68.640 128.795 ;
        RECT 66.970 128.285 68.870 128.455 ;
        RECT 66.610 127.945 68.530 128.115 ;
        RECT 66.610 127.925 66.930 127.945 ;
        RECT 66.160 127.265 66.490 127.775 ;
        RECT 66.760 127.315 66.930 127.925 ;
        RECT 68.700 127.775 68.870 128.285 ;
        RECT 69.040 128.215 69.220 128.625 ;
        RECT 69.390 128.035 69.560 128.795 ;
        RECT 67.660 127.605 68.870 127.775 ;
        RECT 69.040 127.725 69.560 128.035 ;
        RECT 69.730 128.625 70.150 128.965 ;
        RECT 71.020 129.225 72.035 129.425 ;
        RECT 70.440 128.625 70.850 128.955 ;
        RECT 69.730 127.855 69.920 128.625 ;
        RECT 71.020 128.495 71.190 129.225 ;
        RECT 72.335 129.055 72.505 129.385 ;
        RECT 71.360 128.675 71.710 129.045 ;
        RECT 71.020 128.455 71.440 128.495 ;
        RECT 70.090 128.285 71.440 128.455 ;
        RECT 70.090 128.125 70.340 128.285 ;
        RECT 70.850 127.855 71.100 128.115 ;
        RECT 69.730 127.605 71.100 127.855 ;
        RECT 67.660 127.315 67.900 127.605 ;
        RECT 68.700 127.525 68.870 127.605 ;
        RECT 68.700 127.275 69.330 127.525 ;
        RECT 70.300 127.315 70.470 127.605 ;
        RECT 71.270 127.440 71.440 128.285 ;
        RECT 71.890 128.115 72.110 128.985 ;
        RECT 72.335 128.865 73.030 129.055 ;
        RECT 71.610 127.735 72.110 128.115 ;
        RECT 72.280 128.065 72.690 128.685 ;
        RECT 72.860 127.895 73.030 128.865 ;
        RECT 72.335 127.725 73.030 127.895 ;
        RECT 71.270 127.270 72.100 127.440 ;
        RECT 72.335 127.225 72.505 127.725 ;
        RECT 73.220 127.225 73.445 129.345 ;
        RECT 74.115 129.055 74.285 129.345 ;
        RECT 73.620 128.885 74.285 129.055 ;
        RECT 74.745 128.975 75.075 129.335 ;
        RECT 76.115 129.145 76.675 129.435 ;
        RECT 73.620 127.895 73.850 128.885 ;
        RECT 74.745 128.785 76.135 128.975 ;
        RECT 74.020 128.065 74.370 128.715 ;
        RECT 75.965 128.695 76.135 128.785 ;
        RECT 74.560 128.365 75.235 128.615 ;
        RECT 75.455 128.365 75.795 128.615 ;
        RECT 75.965 128.365 76.255 128.695 ;
        RECT 74.560 128.005 74.825 128.365 ;
        RECT 75.965 128.115 76.135 128.365 ;
        RECT 75.195 127.945 76.135 128.115 ;
        RECT 73.620 127.725 74.285 127.895 ;
        RECT 74.115 127.225 74.285 127.725 ;
        RECT 75.195 127.395 75.495 127.945 ;
        RECT 76.425 127.775 76.675 129.145 ;
        RECT 77.045 128.975 77.375 129.335 ;
        RECT 78.415 129.145 78.975 129.435 ;
        RECT 77.045 128.785 78.435 128.975 ;
        RECT 78.265 128.695 78.435 128.785 ;
        RECT 76.860 128.365 77.535 128.615 ;
        RECT 77.755 128.365 78.095 128.615 ;
        RECT 78.265 128.365 78.555 128.695 ;
        RECT 76.860 128.005 77.125 128.365 ;
        RECT 78.265 128.115 78.435 128.365 ;
        RECT 76.215 127.225 76.675 127.775 ;
        RECT 77.495 127.945 78.435 128.115 ;
        RECT 77.495 127.395 77.795 127.945 ;
        RECT 78.725 127.775 78.975 129.145 ;
        RECT 79.420 128.795 79.665 129.400 ;
        RECT 78.515 127.225 78.975 127.775 ;
        RECT 79.145 128.625 80.375 128.795 ;
        RECT 79.145 127.815 79.485 128.625 ;
        RECT 79.655 128.060 80.405 128.250 ;
        RECT 79.145 127.405 79.660 127.815 ;
        RECT 80.235 127.395 80.405 128.060 ;
        RECT 80.575 128.075 80.765 129.435 ;
        RECT 80.935 129.265 81.210 129.435 ;
        RECT 80.935 129.095 81.215 129.265 ;
        RECT 80.935 128.275 81.210 129.095 ;
        RECT 81.400 129.070 81.930 129.435 ;
        RECT 81.755 129.035 81.930 129.070 ;
        RECT 81.415 128.075 81.585 128.875 ;
        RECT 80.575 127.905 81.585 128.075 ;
        RECT 81.755 128.865 82.685 129.035 ;
        RECT 82.855 128.865 83.110 129.435 ;
        RECT 81.755 127.735 81.925 128.865 ;
        RECT 82.515 128.695 82.685 128.865 ;
        RECT 80.800 127.565 81.925 127.735 ;
        RECT 82.095 128.365 82.290 128.695 ;
        RECT 82.515 128.365 82.770 128.695 ;
        RECT 82.095 127.395 82.265 128.365 ;
        RECT 82.940 128.195 83.110 128.865 ;
        RECT 80.235 127.225 82.265 127.395 ;
        RECT 82.775 127.225 83.110 128.195 ;
        RECT 83.285 129.145 83.845 129.435 ;
        RECT 83.285 127.775 83.535 129.145 ;
        RECT 84.885 128.975 85.215 129.335 ;
        RECT 83.825 128.785 85.215 128.975 ;
        RECT 90.100 128.895 90.355 129.425 ;
        RECT 83.825 128.695 83.995 128.785 ;
        RECT 83.705 128.365 83.995 128.695 ;
        RECT 84.165 128.365 84.505 128.615 ;
        RECT 84.725 128.365 85.400 128.615 ;
        RECT 83.825 128.115 83.995 128.365 ;
        RECT 83.825 127.945 84.765 128.115 ;
        RECT 85.135 128.005 85.400 128.365 ;
        RECT 90.100 128.035 90.280 128.895 ;
        RECT 91.000 128.695 91.250 129.345 ;
        RECT 90.450 128.365 91.250 128.695 ;
        RECT 83.285 127.225 83.745 127.775 ;
        RECT 84.465 127.395 84.765 127.945 ;
        RECT 90.100 127.565 90.355 128.035 ;
        RECT 90.015 127.395 90.355 127.565 ;
        RECT 90.100 127.365 90.355 127.395 ;
        RECT 91.000 127.775 91.250 128.365 ;
        RECT 91.450 129.010 91.770 129.340 ;
        RECT 92.810 129.215 93.660 129.385 ;
        RECT 91.450 128.115 91.640 129.010 ;
        RECT 91.960 128.685 92.620 128.955 ;
        RECT 92.290 128.625 92.620 128.685 ;
        RECT 91.810 128.455 92.140 128.515 ;
        RECT 92.810 128.455 92.980 129.215 ;
        RECT 94.740 128.965 94.990 129.395 ;
        RECT 93.150 128.795 94.400 128.965 ;
        RECT 93.150 128.675 93.480 128.795 ;
        RECT 91.810 128.285 93.710 128.455 ;
        RECT 91.450 127.945 93.370 128.115 ;
        RECT 91.450 127.925 91.770 127.945 ;
        RECT 91.000 127.265 91.330 127.775 ;
        RECT 91.600 127.315 91.770 127.925 ;
        RECT 93.540 127.775 93.710 128.285 ;
        RECT 93.880 128.215 94.060 128.625 ;
        RECT 94.230 128.035 94.400 128.795 ;
        RECT 92.500 127.605 93.710 127.775 ;
        RECT 93.880 127.725 94.400 128.035 ;
        RECT 94.570 128.625 94.990 128.965 ;
        RECT 95.860 129.225 96.875 129.425 ;
        RECT 95.280 128.625 95.690 128.955 ;
        RECT 94.570 127.855 94.760 128.625 ;
        RECT 95.860 128.495 96.030 129.225 ;
        RECT 97.175 129.055 97.345 129.385 ;
        RECT 96.200 128.675 96.550 129.045 ;
        RECT 95.860 128.455 96.280 128.495 ;
        RECT 94.930 128.285 96.280 128.455 ;
        RECT 94.930 128.125 95.180 128.285 ;
        RECT 95.690 127.855 95.940 128.115 ;
        RECT 94.570 127.605 95.940 127.855 ;
        RECT 92.500 127.315 92.740 127.605 ;
        RECT 93.540 127.525 93.710 127.605 ;
        RECT 93.540 127.275 94.170 127.525 ;
        RECT 95.140 127.315 95.310 127.605 ;
        RECT 96.110 127.440 96.280 128.285 ;
        RECT 96.730 128.115 96.950 128.985 ;
        RECT 97.175 128.865 97.870 129.055 ;
        RECT 96.450 127.735 96.950 128.115 ;
        RECT 97.120 128.065 97.530 128.685 ;
        RECT 97.700 127.895 97.870 128.865 ;
        RECT 97.175 127.725 97.870 127.895 ;
        RECT 96.110 127.270 96.940 127.440 ;
        RECT 97.175 127.225 97.345 127.725 ;
        RECT 98.060 127.225 98.285 129.345 ;
        RECT 98.955 129.055 99.125 129.345 ;
        RECT 98.460 128.885 99.125 129.055 ;
        RECT 99.585 128.975 99.915 129.335 ;
        RECT 100.955 129.145 101.515 129.435 ;
        RECT 98.460 127.895 98.690 128.885 ;
        RECT 99.585 128.785 100.975 128.975 ;
        RECT 98.860 128.065 99.210 128.715 ;
        RECT 100.805 128.695 100.975 128.785 ;
        RECT 99.400 128.365 100.075 128.615 ;
        RECT 100.295 128.365 100.635 128.615 ;
        RECT 100.805 128.365 101.095 128.695 ;
        RECT 99.400 128.005 99.665 128.365 ;
        RECT 100.805 128.115 100.975 128.365 ;
        RECT 100.035 127.945 100.975 128.115 ;
        RECT 98.460 127.725 99.125 127.895 ;
        RECT 98.955 127.225 99.125 127.725 ;
        RECT 100.035 127.395 100.335 127.945 ;
        RECT 101.265 127.775 101.515 129.145 ;
        RECT 101.055 127.225 101.515 127.775 ;
        RECT 104.445 129.145 105.005 129.435 ;
        RECT 104.445 127.775 104.695 129.145 ;
        RECT 106.045 128.975 106.375 129.335 ;
        RECT 104.985 128.785 106.375 128.975 ;
        RECT 106.745 129.145 107.305 129.435 ;
        RECT 104.985 128.695 105.155 128.785 ;
        RECT 104.865 128.365 105.155 128.695 ;
        RECT 105.325 128.365 105.665 128.615 ;
        RECT 105.885 128.365 106.560 128.615 ;
        RECT 104.985 128.115 105.155 128.365 ;
        RECT 104.985 127.945 105.925 128.115 ;
        RECT 106.295 128.005 106.560 128.365 ;
        RECT 104.445 127.225 104.905 127.775 ;
        RECT 105.625 127.395 105.925 127.945 ;
        RECT 106.745 127.775 106.995 129.145 ;
        RECT 108.345 128.975 108.675 129.335 ;
        RECT 107.285 128.785 108.675 128.975 ;
        RECT 109.045 129.145 109.605 129.435 ;
        RECT 107.285 128.695 107.455 128.785 ;
        RECT 107.165 128.365 107.455 128.695 ;
        RECT 107.625 128.365 107.965 128.615 ;
        RECT 108.185 128.365 108.860 128.615 ;
        RECT 107.285 128.115 107.455 128.365 ;
        RECT 107.285 127.945 108.225 128.115 ;
        RECT 108.595 128.005 108.860 128.365 ;
        RECT 106.745 127.225 107.205 127.775 ;
        RECT 107.925 127.395 108.225 127.945 ;
        RECT 109.045 127.775 109.295 129.145 ;
        RECT 110.645 128.975 110.975 129.335 ;
        RECT 109.585 128.785 110.975 128.975 ;
        RECT 112.315 128.955 112.575 129.345 ;
        RECT 113.175 128.955 113.470 129.345 ;
        RECT 114.095 129.105 114.395 129.435 ;
        RECT 111.820 128.785 113.470 128.955 ;
        RECT 109.585 128.695 109.755 128.785 ;
        RECT 109.465 128.365 109.755 128.695 ;
        RECT 109.925 128.365 110.265 128.615 ;
        RECT 110.485 128.365 111.160 128.615 ;
        RECT 109.585 128.115 109.755 128.365 ;
        RECT 109.585 127.945 110.525 128.115 ;
        RECT 110.895 128.005 111.160 128.365 ;
        RECT 111.820 128.275 112.225 128.785 ;
        RECT 112.395 128.445 113.535 128.615 ;
        RECT 111.820 128.105 112.575 128.275 ;
        RECT 109.045 127.225 109.505 127.775 ;
        RECT 110.225 127.395 110.525 127.945 ;
        RECT 112.315 127.855 112.575 128.105 ;
        RECT 113.365 128.195 113.535 128.445 ;
        RECT 113.705 128.365 114.055 128.935 ;
        RECT 114.225 128.195 114.395 129.105 ;
        RECT 113.365 128.025 114.395 128.195 ;
        RECT 112.315 127.685 113.435 127.855 ;
        RECT 112.315 127.225 112.575 127.685 ;
        RECT 113.175 127.225 113.435 127.685 ;
        RECT 114.085 127.225 114.395 128.025 ;
        RECT 115.025 129.145 115.585 129.435 ;
        RECT 115.025 127.775 115.275 129.145 ;
        RECT 116.625 128.975 116.955 129.335 ;
        RECT 115.565 128.785 116.955 128.975 ;
        RECT 118.685 128.805 119.015 129.435 ;
        RECT 120.175 129.055 120.345 129.435 ;
        RECT 120.175 128.885 120.840 129.055 ;
        RECT 121.035 128.930 121.295 129.435 ;
        RECT 115.565 128.695 115.735 128.785 ;
        RECT 115.445 128.365 115.735 128.695 ;
        RECT 115.905 128.365 116.245 128.615 ;
        RECT 116.465 128.365 117.140 128.615 ;
        RECT 118.265 128.365 118.595 128.615 ;
        RECT 115.565 128.115 115.735 128.365 ;
        RECT 115.565 127.945 116.505 128.115 ;
        RECT 116.875 128.005 117.140 128.365 ;
        RECT 118.765 128.205 119.015 128.805 ;
        RECT 120.105 128.335 120.435 128.705 ;
        RECT 120.670 128.630 120.840 128.885 ;
        RECT 115.025 127.225 115.485 127.775 ;
        RECT 116.205 127.395 116.505 127.945 ;
        RECT 118.685 127.225 119.015 128.205 ;
        RECT 120.670 128.300 120.955 128.630 ;
        RECT 120.670 128.155 120.840 128.300 ;
        RECT 120.175 127.985 120.840 128.155 ;
        RECT 121.125 128.130 121.295 128.930 ;
        RECT 120.175 127.225 120.345 127.985 ;
        RECT 121.025 127.225 121.295 128.130 ;
        RECT 21.165 125.735 21.495 126.715 ;
        RECT 23.115 125.955 23.285 126.715 ;
        RECT 23.115 125.785 23.780 125.955 ;
        RECT 23.965 125.810 24.235 126.715 ;
        RECT 21.165 125.135 21.415 125.735 ;
        RECT 23.610 125.640 23.780 125.785 ;
        RECT 21.585 125.325 21.915 125.575 ;
        RECT 23.045 125.235 23.375 125.605 ;
        RECT 23.610 125.310 23.895 125.640 ;
        RECT 21.165 124.505 21.495 125.135 ;
        RECT 23.610 125.055 23.780 125.310 ;
        RECT 23.115 124.885 23.780 125.055 ;
        RECT 24.065 125.010 24.235 125.810 ;
        RECT 23.115 124.505 23.285 124.885 ;
        RECT 23.975 124.505 24.235 125.010 ;
        RECT 26.250 125.745 26.585 126.715 ;
        RECT 27.095 126.545 29.125 126.715 ;
        RECT 26.250 125.075 26.420 125.745 ;
        RECT 27.095 125.575 27.265 126.545 ;
        RECT 26.590 125.245 26.845 125.575 ;
        RECT 27.070 125.245 27.265 125.575 ;
        RECT 27.435 126.205 28.560 126.375 ;
        RECT 26.675 125.075 26.845 125.245 ;
        RECT 27.435 125.075 27.605 126.205 ;
        RECT 26.250 124.505 26.505 125.075 ;
        RECT 26.675 124.905 27.605 125.075 ;
        RECT 27.775 125.865 28.785 126.035 ;
        RECT 27.775 125.065 27.945 125.865 ;
        RECT 28.150 125.525 28.425 125.665 ;
        RECT 28.145 125.355 28.425 125.525 ;
        RECT 27.430 124.870 27.605 124.905 ;
        RECT 27.430 124.505 27.960 124.870 ;
        RECT 28.150 124.505 28.425 125.355 ;
        RECT 28.595 124.505 28.785 125.865 ;
        RECT 28.955 125.880 29.125 126.545 ;
        RECT 34.235 126.545 36.265 126.715 ;
        RECT 29.700 126.125 30.215 126.535 ;
        RECT 28.955 125.690 29.705 125.880 ;
        RECT 29.875 125.315 30.215 126.125 ;
        RECT 28.985 125.145 30.215 125.315 ;
        RECT 33.145 126.125 33.660 126.535 ;
        RECT 33.145 125.315 33.485 126.125 ;
        RECT 34.235 125.880 34.405 126.545 ;
        RECT 34.800 126.205 35.925 126.375 ;
        RECT 33.655 125.690 34.405 125.880 ;
        RECT 34.575 125.865 35.585 126.035 ;
        RECT 33.145 125.145 34.375 125.315 ;
        RECT 29.695 124.540 29.940 125.145 ;
        RECT 33.420 124.540 33.665 125.145 ;
        RECT 34.575 124.505 34.765 125.865 ;
        RECT 34.935 124.845 35.210 125.665 ;
        RECT 35.415 125.065 35.585 125.865 ;
        RECT 35.755 125.075 35.925 126.205 ;
        RECT 36.095 125.575 36.265 126.545 ;
        RECT 36.775 125.745 37.110 126.715 ;
        RECT 37.935 125.995 38.235 126.545 ;
        RECT 38.955 126.165 39.415 126.715 ;
        RECT 36.095 125.245 36.290 125.575 ;
        RECT 36.515 125.245 36.770 125.575 ;
        RECT 36.515 125.075 36.685 125.245 ;
        RECT 36.940 125.075 37.110 125.745 ;
        RECT 37.300 125.575 37.565 125.935 ;
        RECT 37.935 125.825 38.875 125.995 ;
        RECT 38.705 125.575 38.875 125.825 ;
        RECT 37.300 125.325 37.975 125.575 ;
        RECT 38.195 125.325 38.535 125.575 ;
        RECT 38.705 125.245 38.995 125.575 ;
        RECT 38.705 125.155 38.875 125.245 ;
        RECT 35.755 124.905 36.685 125.075 ;
        RECT 35.755 124.870 35.930 124.905 ;
        RECT 34.935 124.675 35.215 124.845 ;
        RECT 34.935 124.505 35.210 124.675 ;
        RECT 35.400 124.505 35.930 124.870 ;
        RECT 36.855 124.505 37.110 125.075 ;
        RECT 37.485 124.965 38.875 125.155 ;
        RECT 37.485 124.605 37.815 124.965 ;
        RECT 39.165 124.795 39.415 126.165 ;
        RECT 41.155 125.995 41.455 126.545 ;
        RECT 42.175 126.165 42.635 126.715 ;
        RECT 40.520 125.575 40.785 125.935 ;
        RECT 41.155 125.825 42.095 125.995 ;
        RECT 41.925 125.575 42.095 125.825 ;
        RECT 40.520 125.325 41.195 125.575 ;
        RECT 41.415 125.325 41.755 125.575 ;
        RECT 41.925 125.245 42.215 125.575 ;
        RECT 41.925 125.155 42.095 125.245 ;
        RECT 38.855 124.505 39.415 124.795 ;
        RECT 40.705 124.965 42.095 125.155 ;
        RECT 40.705 124.605 41.035 124.965 ;
        RECT 42.385 124.795 42.635 126.165 ;
        RECT 43.455 125.995 43.755 126.545 ;
        RECT 44.475 126.165 44.935 126.715 ;
        RECT 42.820 125.575 43.085 125.935 ;
        RECT 43.455 125.825 44.395 125.995 ;
        RECT 44.225 125.575 44.395 125.825 ;
        RECT 42.820 125.325 43.495 125.575 ;
        RECT 43.715 125.325 44.055 125.575 ;
        RECT 44.225 125.245 44.515 125.575 ;
        RECT 44.225 125.155 44.395 125.245 ;
        RECT 42.075 124.505 42.635 124.795 ;
        RECT 43.005 124.965 44.395 125.155 ;
        RECT 43.005 124.605 43.335 124.965 ;
        RECT 44.685 124.795 44.935 126.165 ;
        RECT 44.375 124.505 44.935 124.795 ;
        RECT 45.105 126.165 45.565 126.715 ;
        RECT 45.105 124.795 45.355 126.165 ;
        RECT 46.285 125.995 46.585 126.545 ;
        RECT 45.645 125.825 46.585 125.995 ;
        RECT 47.915 126.255 48.175 126.715 ;
        RECT 48.775 126.255 49.035 126.715 ;
        RECT 47.915 126.085 49.035 126.255 ;
        RECT 45.645 125.575 45.815 125.825 ;
        RECT 46.955 125.575 47.220 125.935 ;
        RECT 47.915 125.835 48.175 126.085 ;
        RECT 49.685 125.915 49.995 126.715 ;
        RECT 45.525 125.245 45.815 125.575 ;
        RECT 45.985 125.325 46.325 125.575 ;
        RECT 46.545 125.325 47.220 125.575 ;
        RECT 47.420 125.665 48.175 125.835 ;
        RECT 48.965 125.745 49.995 125.915 ;
        RECT 45.645 125.155 45.815 125.245 ;
        RECT 47.420 125.155 47.825 125.665 ;
        RECT 48.965 125.495 49.135 125.745 ;
        RECT 47.995 125.325 49.135 125.495 ;
        RECT 45.645 124.965 47.035 125.155 ;
        RECT 47.420 124.985 49.070 125.155 ;
        RECT 49.305 125.005 49.655 125.575 ;
        RECT 45.105 124.505 45.665 124.795 ;
        RECT 46.705 124.605 47.035 124.965 ;
        RECT 47.915 124.595 48.175 124.985 ;
        RECT 48.775 124.595 49.070 124.985 ;
        RECT 49.825 124.835 49.995 125.745 ;
        RECT 51.570 125.575 51.815 126.715 ;
        RECT 52.430 125.575 52.680 126.710 ;
        RECT 53.280 125.985 53.540 126.710 ;
        RECT 54.140 125.985 54.400 126.710 ;
        RECT 55.000 125.985 55.260 126.710 ;
        RECT 55.860 125.985 56.120 126.710 ;
        RECT 56.705 125.985 56.965 126.710 ;
        RECT 57.565 125.985 57.825 126.710 ;
        RECT 58.425 125.985 58.685 126.710 ;
        RECT 53.280 125.970 58.685 125.985 ;
        RECT 59.295 125.970 59.585 126.710 ;
        RECT 61.375 126.545 63.405 126.715 ;
        RECT 60.285 126.125 60.800 126.535 ;
        RECT 53.280 125.745 60.025 125.970 ;
        RECT 51.085 125.015 51.400 125.575 ;
        RECT 51.570 125.325 58.690 125.575 ;
        RECT 49.695 124.505 49.995 124.835 ;
        RECT 51.570 124.515 51.820 125.325 ;
        RECT 52.430 124.515 52.680 125.325 ;
        RECT 58.860 125.155 60.025 125.745 ;
        RECT 53.280 124.985 60.025 125.155 ;
        RECT 60.285 125.315 60.625 126.125 ;
        RECT 61.375 125.880 61.545 126.545 ;
        RECT 61.940 126.205 63.065 126.375 ;
        RECT 60.795 125.690 61.545 125.880 ;
        RECT 61.715 125.865 62.725 126.035 ;
        RECT 60.285 125.145 61.515 125.315 ;
        RECT 53.280 124.530 53.540 124.985 ;
        RECT 54.140 124.530 54.400 124.985 ;
        RECT 55.000 124.530 55.260 124.985 ;
        RECT 55.845 124.530 56.120 124.985 ;
        RECT 56.705 124.530 56.965 124.985 ;
        RECT 57.565 124.530 57.825 124.985 ;
        RECT 58.425 124.530 58.685 124.985 ;
        RECT 59.295 124.530 59.555 124.985 ;
        RECT 60.560 124.540 60.805 125.145 ;
        RECT 61.715 124.505 61.905 125.865 ;
        RECT 62.075 125.525 62.350 125.665 ;
        RECT 62.075 125.355 62.355 125.525 ;
        RECT 62.075 124.505 62.350 125.355 ;
        RECT 62.555 125.065 62.725 125.865 ;
        RECT 62.895 125.075 63.065 126.205 ;
        RECT 63.235 125.575 63.405 126.545 ;
        RECT 63.915 125.745 64.250 126.715 ;
        RECT 63.235 125.245 63.430 125.575 ;
        RECT 63.655 125.245 63.910 125.575 ;
        RECT 63.655 125.075 63.825 125.245 ;
        RECT 64.080 125.075 64.250 125.745 ;
        RECT 62.895 124.905 63.825 125.075 ;
        RECT 62.895 124.870 63.070 124.905 ;
        RECT 62.540 124.505 63.070 124.870 ;
        RECT 63.995 124.505 64.250 125.075 ;
        RECT 69.005 125.735 69.335 126.715 ;
        RECT 70.035 125.955 70.205 126.715 ;
        RECT 70.035 125.785 70.700 125.955 ;
        RECT 70.885 125.810 71.155 126.715 ;
        RECT 69.005 125.135 69.255 125.735 ;
        RECT 70.530 125.640 70.700 125.785 ;
        RECT 69.425 125.325 69.755 125.575 ;
        RECT 69.965 125.235 70.295 125.605 ;
        RECT 70.530 125.310 70.815 125.640 ;
        RECT 69.005 124.505 69.335 125.135 ;
        RECT 70.530 125.055 70.700 125.310 ;
        RECT 70.035 124.885 70.700 125.055 ;
        RECT 70.985 125.010 71.155 125.810 ;
        RECT 70.035 124.505 70.205 124.885 ;
        RECT 70.895 124.505 71.155 125.010 ;
        RECT 72.705 125.915 73.015 126.715 ;
        RECT 73.665 126.255 73.925 126.715 ;
        RECT 74.525 126.255 74.785 126.715 ;
        RECT 76.760 126.545 77.015 126.575 ;
        RECT 76.675 126.375 77.015 126.545 ;
        RECT 73.665 126.085 74.785 126.255 ;
        RECT 72.705 125.745 73.735 125.915 ;
        RECT 72.705 124.835 72.875 125.745 ;
        RECT 73.045 125.005 73.395 125.575 ;
        RECT 73.565 125.495 73.735 125.745 ;
        RECT 74.525 125.835 74.785 126.085 ;
        RECT 76.760 125.905 77.015 126.375 ;
        RECT 77.660 126.165 77.990 126.675 ;
        RECT 74.525 125.665 75.280 125.835 ;
        RECT 73.565 125.325 74.705 125.495 ;
        RECT 74.875 125.155 75.280 125.665 ;
        RECT 73.630 124.985 75.280 125.155 ;
        RECT 76.760 125.045 76.940 125.905 ;
        RECT 77.660 125.575 77.910 126.165 ;
        RECT 78.260 126.015 78.430 126.625 ;
        RECT 79.160 126.335 79.400 126.625 ;
        RECT 80.200 126.415 80.830 126.665 ;
        RECT 80.200 126.335 80.370 126.415 ;
        RECT 81.800 126.335 81.970 126.625 ;
        RECT 82.770 126.500 83.600 126.670 ;
        RECT 79.160 126.165 80.370 126.335 ;
        RECT 77.110 125.245 77.910 125.575 ;
        RECT 72.705 124.505 73.005 124.835 ;
        RECT 73.630 124.595 73.925 124.985 ;
        RECT 74.525 124.595 74.785 124.985 ;
        RECT 76.760 124.515 77.015 125.045 ;
        RECT 77.660 124.595 77.910 125.245 ;
        RECT 78.110 125.995 78.430 126.015 ;
        RECT 78.110 125.825 80.030 125.995 ;
        RECT 78.110 124.930 78.300 125.825 ;
        RECT 80.200 125.655 80.370 126.165 ;
        RECT 80.540 125.905 81.060 126.215 ;
        RECT 78.470 125.485 80.370 125.655 ;
        RECT 78.470 125.425 78.800 125.485 ;
        RECT 78.950 125.255 79.280 125.315 ;
        RECT 78.620 124.985 79.280 125.255 ;
        RECT 78.110 124.600 78.430 124.930 ;
        RECT 79.470 124.725 79.640 125.485 ;
        RECT 80.540 125.315 80.720 125.725 ;
        RECT 79.810 125.145 80.140 125.265 ;
        RECT 80.890 125.145 81.060 125.905 ;
        RECT 79.810 124.975 81.060 125.145 ;
        RECT 81.230 126.085 82.600 126.335 ;
        RECT 81.230 125.315 81.420 126.085 ;
        RECT 82.350 125.825 82.600 126.085 ;
        RECT 81.590 125.655 81.840 125.815 ;
        RECT 82.770 125.655 82.940 126.500 ;
        RECT 83.835 126.215 84.005 126.715 ;
        RECT 83.110 125.825 83.610 126.205 ;
        RECT 83.835 126.045 84.530 126.215 ;
        RECT 81.590 125.485 82.940 125.655 ;
        RECT 82.520 125.445 82.940 125.485 ;
        RECT 81.230 124.975 81.650 125.315 ;
        RECT 81.940 124.985 82.350 125.315 ;
        RECT 79.470 124.555 80.320 124.725 ;
        RECT 81.400 124.545 81.650 124.975 ;
        RECT 82.520 124.715 82.690 125.445 ;
        RECT 82.860 124.895 83.210 125.265 ;
        RECT 83.390 124.955 83.610 125.825 ;
        RECT 83.780 125.255 84.190 125.875 ;
        RECT 84.360 125.075 84.530 126.045 ;
        RECT 83.835 124.885 84.530 125.075 ;
        RECT 82.520 124.515 83.535 124.715 ;
        RECT 83.835 124.555 84.005 124.885 ;
        RECT 84.720 124.595 84.945 126.715 ;
        RECT 85.615 126.215 85.785 126.715 ;
        RECT 85.120 126.045 85.785 126.215 ;
        RECT 85.120 125.055 85.350 126.045 ;
        RECT 85.520 125.225 85.870 125.875 ;
        RECT 86.495 125.865 86.825 126.715 ;
        RECT 87.335 125.865 87.665 126.715 ;
        RECT 88.175 125.865 88.505 126.715 ;
        RECT 89.015 125.865 89.345 126.715 ;
        RECT 89.855 125.865 90.185 126.715 ;
        RECT 90.695 125.865 91.025 126.715 ;
        RECT 91.535 125.865 91.865 126.715 ;
        RECT 92.375 125.865 92.705 126.715 ;
        RECT 93.215 125.865 93.545 126.715 ;
        RECT 94.055 125.865 94.385 126.715 ;
        RECT 94.895 125.865 95.225 126.715 ;
        RECT 95.735 125.865 96.065 126.715 ;
        RECT 96.575 125.865 96.905 126.715 ;
        RECT 108.295 126.545 110.325 126.715 ;
        RECT 86.045 125.695 92.705 125.865 ;
        RECT 92.875 125.695 95.225 125.865 ;
        RECT 95.395 125.695 96.905 125.865 ;
        RECT 107.205 126.125 107.720 126.535 ;
        RECT 86.045 125.155 86.320 125.695 ;
        RECT 92.875 125.525 93.050 125.695 ;
        RECT 95.395 125.525 95.565 125.695 ;
        RECT 86.490 125.325 93.050 125.525 ;
        RECT 93.255 125.325 95.565 125.525 ;
        RECT 95.735 125.325 96.910 125.525 ;
        RECT 92.875 125.155 93.050 125.325 ;
        RECT 95.395 125.155 95.565 125.325 ;
        RECT 107.205 125.315 107.545 126.125 ;
        RECT 108.295 125.880 108.465 126.545 ;
        RECT 108.860 126.205 109.985 126.375 ;
        RECT 107.715 125.690 108.465 125.880 ;
        RECT 108.635 125.865 109.645 126.035 ;
        RECT 85.120 124.885 85.785 125.055 ;
        RECT 86.045 124.985 92.705 125.155 ;
        RECT 92.875 124.985 95.225 125.155 ;
        RECT 95.395 124.985 96.905 125.155 ;
        RECT 107.205 125.145 108.435 125.315 ;
        RECT 85.615 124.595 85.785 124.885 ;
        RECT 86.495 124.510 86.825 124.985 ;
        RECT 87.335 124.510 87.665 124.985 ;
        RECT 88.175 124.510 88.505 124.985 ;
        RECT 89.015 124.510 89.345 124.985 ;
        RECT 89.855 124.510 90.185 124.985 ;
        RECT 90.695 124.510 91.025 124.985 ;
        RECT 91.535 124.510 91.865 124.985 ;
        RECT 92.375 124.510 92.705 124.985 ;
        RECT 93.215 124.510 93.545 124.985 ;
        RECT 94.055 124.510 94.385 124.985 ;
        RECT 94.895 124.510 95.225 124.985 ;
        RECT 95.735 124.510 96.065 124.985 ;
        RECT 96.575 124.510 96.905 124.985 ;
        RECT 107.480 124.540 107.725 125.145 ;
        RECT 90.775 124.505 90.945 124.510 ;
        RECT 91.615 124.505 91.785 124.510 ;
        RECT 92.455 124.505 92.705 124.510 ;
        RECT 108.635 124.505 108.825 125.865 ;
        RECT 108.995 124.845 109.270 125.665 ;
        RECT 109.475 125.065 109.645 125.865 ;
        RECT 109.815 125.075 109.985 126.205 ;
        RECT 110.155 125.575 110.325 126.545 ;
        RECT 110.835 125.745 111.170 126.715 ;
        RECT 112.435 126.545 114.465 126.715 ;
        RECT 110.155 125.245 110.350 125.575 ;
        RECT 110.575 125.245 110.830 125.575 ;
        RECT 110.575 125.075 110.745 125.245 ;
        RECT 111.000 125.075 111.170 125.745 ;
        RECT 111.345 126.125 111.860 126.535 ;
        RECT 111.345 125.315 111.685 126.125 ;
        RECT 112.435 125.880 112.605 126.545 ;
        RECT 113.000 126.205 114.125 126.375 ;
        RECT 111.855 125.690 112.605 125.880 ;
        RECT 112.775 125.865 113.785 126.035 ;
        RECT 111.345 125.145 112.575 125.315 ;
        RECT 109.815 124.905 110.745 125.075 ;
        RECT 109.815 124.870 109.990 124.905 ;
        RECT 108.995 124.675 109.275 124.845 ;
        RECT 108.995 124.505 109.270 124.675 ;
        RECT 109.460 124.505 109.990 124.870 ;
        RECT 110.915 124.505 111.170 125.075 ;
        RECT 111.620 124.540 111.865 125.145 ;
        RECT 112.775 124.505 112.965 125.865 ;
        RECT 113.135 125.185 113.410 125.665 ;
        RECT 113.135 125.015 113.415 125.185 ;
        RECT 113.615 125.065 113.785 125.865 ;
        RECT 113.955 125.075 114.125 126.205 ;
        RECT 114.295 125.575 114.465 126.545 ;
        RECT 114.975 125.745 115.310 126.715 ;
        RECT 114.295 125.245 114.490 125.575 ;
        RECT 114.715 125.245 114.970 125.575 ;
        RECT 114.715 125.075 114.885 125.245 ;
        RECT 115.140 125.075 115.310 125.745 ;
        RECT 115.860 125.905 116.115 126.575 ;
        RECT 116.760 126.165 117.090 126.675 ;
        RECT 115.860 125.185 116.040 125.905 ;
        RECT 116.760 125.575 117.010 126.165 ;
        RECT 117.360 126.015 117.530 126.625 ;
        RECT 118.260 126.335 118.500 126.625 ;
        RECT 119.300 126.415 119.930 126.665 ;
        RECT 119.300 126.335 119.470 126.415 ;
        RECT 120.900 126.335 121.070 126.625 ;
        RECT 121.870 126.500 122.700 126.670 ;
        RECT 118.260 126.165 119.470 126.335 ;
        RECT 116.210 125.245 117.010 125.575 ;
        RECT 113.135 124.505 113.410 125.015 ;
        RECT 113.955 124.905 114.885 125.075 ;
        RECT 113.955 124.870 114.130 124.905 ;
        RECT 113.600 124.505 114.130 124.870 ;
        RECT 115.055 124.505 115.310 125.075 ;
        RECT 115.775 125.045 116.040 125.185 ;
        RECT 115.775 125.015 116.115 125.045 ;
        RECT 115.860 124.515 116.115 125.015 ;
        RECT 116.760 124.595 117.010 125.245 ;
        RECT 117.210 125.995 117.530 126.015 ;
        RECT 117.210 125.825 119.130 125.995 ;
        RECT 117.210 124.930 117.400 125.825 ;
        RECT 119.300 125.655 119.470 126.165 ;
        RECT 119.640 125.905 120.160 126.215 ;
        RECT 117.570 125.485 119.470 125.655 ;
        RECT 117.570 125.425 117.900 125.485 ;
        RECT 118.050 125.255 118.380 125.315 ;
        RECT 117.720 124.985 118.380 125.255 ;
        RECT 117.210 124.600 117.530 124.930 ;
        RECT 118.570 124.725 118.740 125.485 ;
        RECT 119.640 125.315 119.820 125.725 ;
        RECT 118.910 125.145 119.240 125.265 ;
        RECT 119.990 125.145 120.160 125.905 ;
        RECT 118.910 124.975 120.160 125.145 ;
        RECT 120.330 126.085 121.700 126.335 ;
        RECT 120.330 125.315 120.520 126.085 ;
        RECT 121.450 125.825 121.700 126.085 ;
        RECT 120.690 125.655 120.940 125.815 ;
        RECT 121.870 125.655 122.040 126.500 ;
        RECT 122.935 126.215 123.105 126.715 ;
        RECT 122.210 125.825 122.710 126.205 ;
        RECT 122.935 126.045 123.630 126.215 ;
        RECT 120.690 125.485 122.040 125.655 ;
        RECT 121.620 125.445 122.040 125.485 ;
        RECT 120.330 124.975 120.750 125.315 ;
        RECT 121.040 124.985 121.450 125.315 ;
        RECT 118.570 124.555 119.420 124.725 ;
        RECT 120.500 124.545 120.750 124.975 ;
        RECT 121.620 124.715 121.790 125.445 ;
        RECT 121.960 124.895 122.310 125.265 ;
        RECT 122.490 124.955 122.710 125.825 ;
        RECT 122.880 125.255 123.290 125.875 ;
        RECT 123.460 125.075 123.630 126.045 ;
        RECT 122.935 124.885 123.630 125.075 ;
        RECT 121.620 124.515 122.635 124.715 ;
        RECT 122.935 124.555 123.105 124.885 ;
        RECT 123.820 124.595 124.045 126.715 ;
        RECT 124.715 126.215 124.885 126.715 ;
        RECT 124.220 126.045 124.885 126.215 ;
        RECT 124.220 125.055 124.450 126.045 ;
        RECT 124.620 125.225 124.970 125.875 ;
        RECT 124.220 124.885 124.885 125.055 ;
        RECT 124.715 124.595 124.885 124.885 ;
        RECT 17.045 122.925 17.360 123.485 ;
        RECT 17.530 123.175 17.780 123.985 ;
        RECT 18.390 123.175 18.640 123.985 ;
        RECT 19.240 123.515 19.500 123.970 ;
        RECT 20.100 123.515 20.360 123.970 ;
        RECT 20.960 123.515 21.220 123.970 ;
        RECT 21.805 123.515 22.080 123.970 ;
        RECT 22.665 123.515 22.925 123.970 ;
        RECT 23.525 123.515 23.785 123.970 ;
        RECT 24.385 123.515 24.645 123.970 ;
        RECT 25.255 123.515 25.515 123.970 ;
        RECT 28.645 123.515 28.905 123.970 ;
        RECT 29.515 123.515 29.775 123.970 ;
        RECT 30.375 123.515 30.635 123.970 ;
        RECT 31.235 123.515 31.495 123.970 ;
        RECT 32.080 123.515 32.355 123.970 ;
        RECT 32.940 123.515 33.200 123.970 ;
        RECT 33.800 123.515 34.060 123.970 ;
        RECT 34.660 123.515 34.920 123.970 ;
        RECT 19.240 123.345 25.985 123.515 ;
        RECT 28.175 123.485 34.920 123.515 ;
        RECT 17.530 122.925 24.650 123.175 ;
        RECT 17.530 121.785 17.775 122.925 ;
        RECT 18.390 121.790 18.640 122.925 ;
        RECT 24.820 122.755 25.985 123.345 ;
        RECT 28.145 123.345 34.920 123.485 ;
        RECT 28.145 123.315 29.340 123.345 ;
        RECT 19.240 122.530 25.985 122.755 ;
        RECT 28.175 122.755 29.340 123.315 ;
        RECT 35.520 123.175 35.770 123.985 ;
        RECT 36.380 123.175 36.630 123.985 ;
        RECT 29.510 122.925 36.630 123.175 ;
        RECT 36.800 122.925 37.115 123.485 ;
        RECT 38.020 123.355 38.265 123.960 ;
        RECT 37.745 123.185 38.975 123.355 ;
        RECT 28.175 122.530 34.920 122.755 ;
        RECT 19.240 122.515 24.645 122.530 ;
        RECT 19.240 121.790 19.500 122.515 ;
        RECT 20.100 121.790 20.360 122.515 ;
        RECT 20.960 121.790 21.220 122.515 ;
        RECT 21.820 121.790 22.080 122.515 ;
        RECT 22.665 121.790 22.925 122.515 ;
        RECT 23.525 121.790 23.785 122.515 ;
        RECT 24.385 121.790 24.645 122.515 ;
        RECT 25.255 121.790 25.545 122.530 ;
        RECT 28.615 121.790 28.905 122.530 ;
        RECT 29.515 122.515 34.920 122.530 ;
        RECT 29.515 121.790 29.775 122.515 ;
        RECT 30.375 121.790 30.635 122.515 ;
        RECT 31.235 121.790 31.495 122.515 ;
        RECT 32.080 121.790 32.340 122.515 ;
        RECT 32.940 121.790 33.200 122.515 ;
        RECT 33.800 121.790 34.060 122.515 ;
        RECT 34.660 121.790 34.920 122.515 ;
        RECT 35.520 121.790 35.770 122.925 ;
        RECT 36.385 121.785 36.630 122.925 ;
        RECT 37.745 122.375 38.085 123.185 ;
        RECT 38.255 122.620 39.005 122.810 ;
        RECT 37.745 121.965 38.260 122.375 ;
        RECT 38.835 121.955 39.005 122.620 ;
        RECT 39.175 122.635 39.365 123.995 ;
        RECT 39.535 123.145 39.810 123.995 ;
        RECT 40.000 123.630 40.530 123.995 ;
        RECT 40.355 123.595 40.530 123.630 ;
        RECT 39.535 122.975 39.815 123.145 ;
        RECT 39.535 122.835 39.810 122.975 ;
        RECT 40.015 122.635 40.185 123.435 ;
        RECT 39.175 122.465 40.185 122.635 ;
        RECT 40.355 123.425 41.285 123.595 ;
        RECT 41.455 123.425 41.710 123.995 ;
        RECT 53.300 123.825 53.555 123.985 ;
        RECT 53.215 123.655 53.555 123.825 ;
        RECT 40.355 122.295 40.525 123.425 ;
        RECT 41.115 123.255 41.285 123.425 ;
        RECT 39.400 122.125 40.525 122.295 ;
        RECT 40.695 122.925 40.890 123.255 ;
        RECT 41.115 122.925 41.370 123.255 ;
        RECT 40.695 121.955 40.865 122.925 ;
        RECT 41.540 122.755 41.710 123.425 ;
        RECT 38.835 121.785 40.865 121.955 ;
        RECT 41.375 121.785 41.710 122.755 ;
        RECT 53.300 123.455 53.555 123.655 ;
        RECT 53.300 122.595 53.480 123.455 ;
        RECT 54.200 123.255 54.450 123.905 ;
        RECT 53.650 122.925 54.450 123.255 ;
        RECT 53.300 121.925 53.555 122.595 ;
        RECT 54.200 122.335 54.450 122.925 ;
        RECT 54.650 123.570 54.970 123.900 ;
        RECT 56.010 123.775 56.860 123.945 ;
        RECT 54.650 122.675 54.840 123.570 ;
        RECT 55.160 123.245 55.820 123.515 ;
        RECT 55.490 123.185 55.820 123.245 ;
        RECT 55.010 123.015 55.340 123.075 ;
        RECT 56.010 123.015 56.180 123.775 ;
        RECT 57.940 123.525 58.190 123.955 ;
        RECT 56.350 123.355 57.600 123.525 ;
        RECT 56.350 123.235 56.680 123.355 ;
        RECT 55.010 122.845 56.910 123.015 ;
        RECT 54.650 122.505 56.570 122.675 ;
        RECT 54.650 122.485 54.970 122.505 ;
        RECT 54.200 121.825 54.530 122.335 ;
        RECT 54.800 121.875 54.970 122.485 ;
        RECT 56.740 122.335 56.910 122.845 ;
        RECT 57.080 122.775 57.260 123.185 ;
        RECT 57.430 122.595 57.600 123.355 ;
        RECT 55.700 122.165 56.910 122.335 ;
        RECT 57.080 122.285 57.600 122.595 ;
        RECT 57.770 123.185 58.190 123.525 ;
        RECT 59.060 123.785 60.075 123.985 ;
        RECT 58.480 123.185 58.890 123.515 ;
        RECT 57.770 122.415 57.960 123.185 ;
        RECT 59.060 123.055 59.230 123.785 ;
        RECT 60.375 123.615 60.545 123.945 ;
        RECT 59.400 123.235 59.750 123.605 ;
        RECT 59.060 123.015 59.480 123.055 ;
        RECT 58.130 122.845 59.480 123.015 ;
        RECT 58.130 122.685 58.380 122.845 ;
        RECT 58.890 122.415 59.140 122.675 ;
        RECT 57.770 122.165 59.140 122.415 ;
        RECT 55.700 121.875 55.940 122.165 ;
        RECT 56.740 122.085 56.910 122.165 ;
        RECT 56.740 121.835 57.370 122.085 ;
        RECT 58.340 121.875 58.510 122.165 ;
        RECT 59.310 122.000 59.480 122.845 ;
        RECT 59.930 122.675 60.150 123.545 ;
        RECT 60.375 123.425 61.070 123.615 ;
        RECT 59.650 122.295 60.150 122.675 ;
        RECT 60.320 122.625 60.730 123.245 ;
        RECT 60.900 122.455 61.070 123.425 ;
        RECT 60.375 122.285 61.070 122.455 ;
        RECT 59.310 121.830 60.140 122.000 ;
        RECT 60.375 121.785 60.545 122.285 ;
        RECT 61.260 121.785 61.485 123.905 ;
        RECT 62.155 123.615 62.325 123.905 ;
        RECT 61.660 123.445 62.325 123.615 ;
        RECT 61.660 122.455 61.890 123.445 ;
        RECT 63.780 123.355 64.025 123.960 ;
        RECT 62.060 122.625 62.410 123.275 ;
        RECT 63.505 123.185 64.735 123.355 ;
        RECT 61.660 122.285 62.325 122.455 ;
        RECT 62.155 121.785 62.325 122.285 ;
        RECT 63.505 122.375 63.845 123.185 ;
        RECT 64.015 122.620 64.765 122.810 ;
        RECT 63.505 121.965 64.020 122.375 ;
        RECT 64.595 121.955 64.765 122.620 ;
        RECT 64.935 122.635 65.125 123.995 ;
        RECT 65.295 123.825 65.570 123.995 ;
        RECT 65.295 123.655 65.575 123.825 ;
        RECT 65.295 122.835 65.570 123.655 ;
        RECT 65.760 123.630 66.290 123.995 ;
        RECT 66.115 123.595 66.290 123.630 ;
        RECT 65.775 122.635 65.945 123.435 ;
        RECT 64.935 122.465 65.945 122.635 ;
        RECT 66.115 123.425 67.045 123.595 ;
        RECT 67.215 123.425 67.470 123.995 ;
        RECT 66.115 122.295 66.285 123.425 ;
        RECT 66.875 123.255 67.045 123.425 ;
        RECT 65.160 122.125 66.285 122.295 ;
        RECT 66.455 122.925 66.650 123.255 ;
        RECT 66.875 122.925 67.130 123.255 ;
        RECT 66.455 121.955 66.625 122.925 ;
        RECT 67.300 122.755 67.470 123.425 ;
        RECT 64.595 121.785 66.625 121.955 ;
        RECT 67.135 121.785 67.470 122.755 ;
        RECT 81.885 123.365 82.215 123.995 ;
        RECT 83.375 123.615 83.545 123.995 ;
        RECT 83.375 123.445 84.040 123.615 ;
        RECT 84.235 123.490 84.495 123.995 ;
        RECT 81.885 122.765 82.135 123.365 ;
        RECT 82.305 122.925 82.635 123.175 ;
        RECT 83.305 122.895 83.635 123.265 ;
        RECT 83.870 123.190 84.040 123.445 ;
        RECT 83.870 122.860 84.155 123.190 ;
        RECT 81.885 121.785 82.215 122.765 ;
        RECT 83.870 122.715 84.040 122.860 ;
        RECT 83.375 122.545 84.040 122.715 ;
        RECT 84.325 122.690 84.495 123.490 ;
        RECT 89.265 122.925 89.580 123.485 ;
        RECT 89.750 123.175 90.000 123.985 ;
        RECT 90.610 123.175 90.860 123.985 ;
        RECT 91.460 123.515 91.720 123.970 ;
        RECT 92.320 123.515 92.580 123.970 ;
        RECT 93.180 123.515 93.440 123.970 ;
        RECT 94.025 123.515 94.300 123.970 ;
        RECT 94.885 123.515 95.145 123.970 ;
        RECT 95.745 123.515 96.005 123.970 ;
        RECT 96.605 123.515 96.865 123.970 ;
        RECT 97.475 123.515 97.735 123.970 ;
        RECT 91.460 123.345 98.205 123.515 ;
        RECT 89.750 122.925 96.870 123.175 ;
        RECT 83.375 121.785 83.545 122.545 ;
        RECT 84.225 121.785 84.495 122.690 ;
        RECT 89.750 121.785 89.995 122.925 ;
        RECT 90.610 121.790 90.860 122.925 ;
        RECT 97.040 122.805 98.205 123.345 ;
        RECT 105.365 122.925 105.680 123.485 ;
        RECT 105.850 123.175 106.100 123.985 ;
        RECT 106.710 123.175 106.960 123.985 ;
        RECT 107.560 123.515 107.820 123.970 ;
        RECT 108.420 123.515 108.680 123.970 ;
        RECT 109.280 123.515 109.540 123.970 ;
        RECT 110.125 123.515 110.400 123.970 ;
        RECT 110.985 123.515 111.245 123.970 ;
        RECT 111.845 123.515 112.105 123.970 ;
        RECT 112.705 123.515 112.965 123.970 ;
        RECT 113.575 123.515 113.835 123.970 ;
        RECT 107.560 123.345 114.305 123.515 ;
        RECT 105.850 122.925 112.970 123.175 ;
        RECT 97.040 122.755 98.235 122.805 ;
        RECT 91.460 122.635 98.235 122.755 ;
        RECT 91.460 122.530 98.205 122.635 ;
        RECT 91.460 122.515 96.865 122.530 ;
        RECT 91.460 121.790 91.720 122.515 ;
        RECT 92.320 121.790 92.580 122.515 ;
        RECT 93.180 121.790 93.440 122.515 ;
        RECT 94.040 121.790 94.300 122.515 ;
        RECT 94.885 121.790 95.145 122.515 ;
        RECT 95.745 121.790 96.005 122.515 ;
        RECT 96.605 121.790 96.865 122.515 ;
        RECT 97.475 121.790 97.765 122.530 ;
        RECT 105.850 121.785 106.095 122.925 ;
        RECT 106.710 121.790 106.960 122.925 ;
        RECT 113.140 122.755 114.305 123.345 ;
        RECT 107.560 122.530 114.305 122.755 ;
        RECT 115.860 123.455 116.115 123.985 ;
        RECT 115.860 122.595 116.040 123.455 ;
        RECT 116.760 123.255 117.010 123.905 ;
        RECT 116.210 122.925 117.010 123.255 ;
        RECT 107.560 122.515 112.965 122.530 ;
        RECT 107.560 121.790 107.820 122.515 ;
        RECT 108.420 121.790 108.680 122.515 ;
        RECT 109.280 121.790 109.540 122.515 ;
        RECT 110.140 121.790 110.400 122.515 ;
        RECT 110.985 121.790 111.245 122.515 ;
        RECT 111.845 121.790 112.105 122.515 ;
        RECT 112.705 121.790 112.965 122.515 ;
        RECT 113.575 121.790 113.865 122.530 ;
        RECT 115.860 122.125 116.115 122.595 ;
        RECT 115.775 121.955 116.115 122.125 ;
        RECT 115.860 121.925 116.115 121.955 ;
        RECT 116.760 122.335 117.010 122.925 ;
        RECT 117.210 123.570 117.530 123.900 ;
        RECT 118.570 123.775 119.420 123.945 ;
        RECT 117.210 122.675 117.400 123.570 ;
        RECT 117.720 123.245 118.380 123.515 ;
        RECT 118.050 123.185 118.380 123.245 ;
        RECT 117.570 123.015 117.900 123.075 ;
        RECT 118.570 123.015 118.740 123.775 ;
        RECT 120.500 123.525 120.750 123.955 ;
        RECT 118.910 123.355 120.160 123.525 ;
        RECT 118.910 123.235 119.240 123.355 ;
        RECT 117.570 122.845 119.470 123.015 ;
        RECT 117.210 122.505 119.130 122.675 ;
        RECT 117.210 122.485 117.530 122.505 ;
        RECT 116.760 121.825 117.090 122.335 ;
        RECT 117.360 121.875 117.530 122.485 ;
        RECT 119.300 122.335 119.470 122.845 ;
        RECT 119.640 122.775 119.820 123.185 ;
        RECT 119.990 122.595 120.160 123.355 ;
        RECT 118.260 122.165 119.470 122.335 ;
        RECT 119.640 122.285 120.160 122.595 ;
        RECT 120.330 123.185 120.750 123.525 ;
        RECT 121.620 123.785 122.635 123.985 ;
        RECT 121.040 123.185 121.450 123.515 ;
        RECT 120.330 122.415 120.520 123.185 ;
        RECT 121.620 123.055 121.790 123.785 ;
        RECT 122.935 123.615 123.105 123.945 ;
        RECT 121.960 123.235 122.310 123.605 ;
        RECT 121.620 123.015 122.040 123.055 ;
        RECT 120.690 122.845 122.040 123.015 ;
        RECT 120.690 122.685 120.940 122.845 ;
        RECT 121.450 122.415 121.700 122.675 ;
        RECT 120.330 122.165 121.700 122.415 ;
        RECT 118.260 121.875 118.500 122.165 ;
        RECT 119.300 122.085 119.470 122.165 ;
        RECT 119.300 121.835 119.930 122.085 ;
        RECT 120.900 121.875 121.070 122.165 ;
        RECT 121.870 122.000 122.040 122.845 ;
        RECT 122.490 122.675 122.710 123.545 ;
        RECT 122.935 123.425 123.630 123.615 ;
        RECT 122.210 122.295 122.710 122.675 ;
        RECT 122.880 122.625 123.290 123.245 ;
        RECT 123.460 122.455 123.630 123.425 ;
        RECT 122.935 122.285 123.630 122.455 ;
        RECT 121.870 121.830 122.700 122.000 ;
        RECT 122.935 121.785 123.105 122.285 ;
        RECT 123.820 121.785 124.045 123.905 ;
        RECT 124.715 123.615 124.885 123.905 ;
        RECT 124.220 123.445 124.885 123.615 ;
        RECT 124.220 122.455 124.450 123.445 ;
        RECT 124.620 122.625 124.970 123.275 ;
        RECT 124.220 122.285 124.885 122.455 ;
        RECT 124.715 121.785 124.885 122.285 ;
        RECT 21.355 121.105 23.385 121.275 ;
        RECT 20.265 120.685 20.780 121.095 ;
        RECT 20.265 119.875 20.605 120.685 ;
        RECT 21.355 120.440 21.525 121.105 ;
        RECT 21.920 120.765 23.045 120.935 ;
        RECT 20.775 120.250 21.525 120.440 ;
        RECT 21.695 120.425 22.705 120.595 ;
        RECT 20.265 119.705 21.495 119.875 ;
        RECT 20.540 119.100 20.785 119.705 ;
        RECT 21.695 119.065 21.885 120.425 ;
        RECT 22.055 119.405 22.330 120.225 ;
        RECT 22.535 119.625 22.705 120.425 ;
        RECT 22.875 119.635 23.045 120.765 ;
        RECT 23.215 120.135 23.385 121.105 ;
        RECT 23.895 120.305 24.230 121.275 ;
        RECT 23.215 119.805 23.410 120.135 ;
        RECT 23.635 119.805 23.890 120.135 ;
        RECT 23.635 119.635 23.805 119.805 ;
        RECT 24.060 119.635 24.230 120.305 ;
        RECT 22.875 119.465 23.805 119.635 ;
        RECT 22.875 119.430 23.050 119.465 ;
        RECT 22.055 119.235 22.335 119.405 ;
        RECT 22.055 119.065 22.330 119.235 ;
        RECT 22.520 119.065 23.050 119.430 ;
        RECT 23.975 119.065 24.230 119.635 ;
        RECT 25.785 120.370 26.055 121.275 ;
        RECT 26.735 120.515 26.905 121.275 ;
        RECT 25.785 119.570 25.955 120.370 ;
        RECT 26.240 120.345 26.905 120.515 ;
        RECT 26.240 120.200 26.410 120.345 ;
        RECT 29.905 120.295 30.235 121.275 ;
        RECT 31.285 120.295 31.615 121.275 ;
        RECT 32.600 121.105 32.855 121.135 ;
        RECT 32.515 120.935 32.855 121.105 ;
        RECT 26.125 119.870 26.410 120.200 ;
        RECT 26.240 119.615 26.410 119.870 ;
        RECT 26.645 119.795 26.975 120.165 ;
        RECT 29.485 119.885 29.815 120.135 ;
        RECT 29.985 119.695 30.235 120.295 ;
        RECT 30.865 119.885 31.195 120.135 ;
        RECT 31.365 119.695 31.615 120.295 ;
        RECT 25.785 119.065 26.045 119.570 ;
        RECT 26.240 119.445 26.905 119.615 ;
        RECT 26.735 119.065 26.905 119.445 ;
        RECT 29.905 119.065 30.235 119.695 ;
        RECT 31.285 119.065 31.615 119.695 ;
        RECT 32.600 120.465 32.855 120.935 ;
        RECT 33.500 120.725 33.830 121.235 ;
        RECT 32.600 119.605 32.780 120.465 ;
        RECT 33.500 120.135 33.750 120.725 ;
        RECT 34.100 120.575 34.270 121.185 ;
        RECT 35.000 120.895 35.240 121.185 ;
        RECT 36.040 120.975 36.670 121.225 ;
        RECT 36.040 120.895 36.210 120.975 ;
        RECT 37.640 120.895 37.810 121.185 ;
        RECT 38.610 121.060 39.440 121.230 ;
        RECT 35.000 120.725 36.210 120.895 ;
        RECT 32.950 119.805 33.750 120.135 ;
        RECT 32.600 119.075 32.855 119.605 ;
        RECT 33.500 119.155 33.750 119.805 ;
        RECT 33.950 120.555 34.270 120.575 ;
        RECT 33.950 120.385 35.870 120.555 ;
        RECT 33.950 119.490 34.140 120.385 ;
        RECT 36.040 120.215 36.210 120.725 ;
        RECT 36.380 120.465 36.900 120.775 ;
        RECT 34.310 120.045 36.210 120.215 ;
        RECT 34.310 119.985 34.640 120.045 ;
        RECT 34.790 119.815 35.120 119.875 ;
        RECT 34.460 119.545 35.120 119.815 ;
        RECT 33.950 119.160 34.270 119.490 ;
        RECT 35.310 119.285 35.480 120.045 ;
        RECT 36.380 119.875 36.560 120.285 ;
        RECT 35.650 119.705 35.980 119.825 ;
        RECT 36.730 119.705 36.900 120.465 ;
        RECT 35.650 119.535 36.900 119.705 ;
        RECT 37.070 120.645 38.440 120.895 ;
        RECT 37.070 119.875 37.260 120.645 ;
        RECT 38.190 120.385 38.440 120.645 ;
        RECT 37.430 120.215 37.680 120.375 ;
        RECT 38.610 120.215 38.780 121.060 ;
        RECT 39.675 120.775 39.845 121.275 ;
        RECT 38.950 120.385 39.450 120.765 ;
        RECT 39.675 120.605 40.370 120.775 ;
        RECT 37.430 120.045 38.780 120.215 ;
        RECT 38.360 120.005 38.780 120.045 ;
        RECT 37.070 119.535 37.490 119.875 ;
        RECT 37.780 119.545 38.190 119.875 ;
        RECT 35.310 119.115 36.160 119.285 ;
        RECT 37.240 119.105 37.490 119.535 ;
        RECT 38.360 119.275 38.530 120.005 ;
        RECT 38.700 119.455 39.050 119.825 ;
        RECT 39.230 119.515 39.450 120.385 ;
        RECT 39.620 119.815 40.030 120.435 ;
        RECT 40.200 119.635 40.370 120.605 ;
        RECT 39.675 119.445 40.370 119.635 ;
        RECT 38.360 119.075 39.375 119.275 ;
        RECT 39.675 119.115 39.845 119.445 ;
        RECT 40.560 119.155 40.785 121.275 ;
        RECT 41.455 120.775 41.625 121.275 ;
        RECT 42.975 121.105 45.005 121.275 ;
        RECT 40.960 120.605 41.625 120.775 ;
        RECT 41.885 120.685 42.400 121.095 ;
        RECT 40.960 119.615 41.190 120.605 ;
        RECT 41.360 119.785 41.710 120.435 ;
        RECT 41.885 119.875 42.225 120.685 ;
        RECT 42.975 120.440 43.145 121.105 ;
        RECT 43.540 120.765 44.665 120.935 ;
        RECT 42.395 120.250 43.145 120.440 ;
        RECT 43.315 120.425 44.325 120.595 ;
        RECT 41.885 119.705 43.115 119.875 ;
        RECT 40.960 119.445 41.625 119.615 ;
        RECT 41.455 119.155 41.625 119.445 ;
        RECT 42.160 119.100 42.405 119.705 ;
        RECT 43.315 119.065 43.505 120.425 ;
        RECT 43.675 119.405 43.950 120.225 ;
        RECT 44.155 119.625 44.325 120.425 ;
        RECT 44.495 119.635 44.665 120.765 ;
        RECT 44.835 120.135 45.005 121.105 ;
        RECT 45.515 120.305 45.850 121.275 ;
        RECT 47.115 121.105 49.145 121.275 ;
        RECT 44.835 119.805 45.030 120.135 ;
        RECT 45.255 119.805 45.510 120.135 ;
        RECT 45.255 119.635 45.425 119.805 ;
        RECT 45.680 119.635 45.850 120.305 ;
        RECT 46.025 120.685 46.540 121.095 ;
        RECT 46.025 119.875 46.365 120.685 ;
        RECT 47.115 120.440 47.285 121.105 ;
        RECT 47.680 120.765 48.805 120.935 ;
        RECT 46.535 120.250 47.285 120.440 ;
        RECT 47.455 120.425 48.465 120.595 ;
        RECT 46.025 119.705 47.255 119.875 ;
        RECT 44.495 119.465 45.425 119.635 ;
        RECT 44.495 119.430 44.670 119.465 ;
        RECT 43.675 119.235 43.955 119.405 ;
        RECT 43.675 119.065 43.950 119.235 ;
        RECT 44.140 119.065 44.670 119.430 ;
        RECT 45.595 119.065 45.850 119.635 ;
        RECT 46.300 119.100 46.545 119.705 ;
        RECT 47.455 119.065 47.645 120.425 ;
        RECT 47.815 119.745 48.090 120.225 ;
        RECT 47.815 119.575 48.095 119.745 ;
        RECT 48.295 119.625 48.465 120.425 ;
        RECT 48.635 119.635 48.805 120.765 ;
        RECT 48.975 120.135 49.145 121.105 ;
        RECT 49.655 120.305 49.990 121.275 ;
        RECT 48.975 119.805 49.170 120.135 ;
        RECT 49.395 119.805 49.650 120.135 ;
        RECT 49.395 119.635 49.565 119.805 ;
        RECT 49.820 119.635 49.990 120.305 ;
        RECT 51.065 120.295 51.395 121.275 ;
        RECT 50.645 119.885 50.975 120.135 ;
        RECT 51.145 119.695 51.395 120.295 ;
        RECT 47.815 119.065 48.090 119.575 ;
        RECT 48.635 119.465 49.565 119.635 ;
        RECT 48.635 119.430 48.810 119.465 ;
        RECT 48.280 119.065 48.810 119.430 ;
        RECT 49.735 119.065 49.990 119.635 ;
        RECT 51.065 119.065 51.395 119.695 ;
        RECT 54.035 120.425 54.205 121.275 ;
        RECT 54.875 120.425 55.045 121.275 ;
        RECT 55.635 120.465 55.965 121.275 ;
        RECT 54.035 120.255 55.045 120.425 ;
        RECT 55.250 120.295 55.965 120.465 ;
        RECT 54.035 120.085 54.530 120.255 ;
        RECT 54.035 119.915 54.535 120.085 ;
        RECT 55.250 120.055 55.420 120.295 ;
        RECT 54.035 119.715 54.530 119.915 ;
        RECT 54.920 119.885 55.420 120.055 ;
        RECT 55.590 119.885 55.970 120.125 ;
        RECT 57.265 120.105 57.595 121.275 ;
        RECT 58.325 120.105 58.685 121.275 ;
        RECT 59.740 121.105 59.995 121.135 ;
        RECT 59.655 120.935 59.995 121.105 ;
        RECT 59.740 120.465 59.995 120.935 ;
        RECT 60.640 120.725 60.970 121.235 ;
        RECT 55.250 119.715 55.420 119.885 ;
        RECT 57.265 119.825 58.685 120.105 ;
        RECT 54.035 119.545 55.045 119.715 ;
        RECT 55.250 119.545 55.885 119.715 ;
        RECT 54.035 119.065 54.205 119.545 ;
        RECT 54.875 119.065 55.045 119.545 ;
        RECT 55.715 119.065 55.885 119.545 ;
        RECT 58.325 119.490 58.685 119.825 ;
        RECT 58.855 119.555 59.195 120.135 ;
        RECT 59.740 119.605 59.920 120.465 ;
        RECT 60.640 120.135 60.890 120.725 ;
        RECT 61.240 120.575 61.410 121.185 ;
        RECT 62.140 120.895 62.380 121.185 ;
        RECT 63.180 120.975 63.810 121.225 ;
        RECT 63.180 120.895 63.350 120.975 ;
        RECT 64.780 120.895 64.950 121.185 ;
        RECT 65.750 121.060 66.580 121.230 ;
        RECT 62.140 120.725 63.350 120.895 ;
        RECT 60.090 119.805 60.890 120.135 ;
        RECT 58.065 119.065 58.685 119.490 ;
        RECT 59.740 119.075 59.995 119.605 ;
        RECT 60.640 119.155 60.890 119.805 ;
        RECT 61.090 120.555 61.410 120.575 ;
        RECT 61.090 120.385 63.010 120.555 ;
        RECT 61.090 119.490 61.280 120.385 ;
        RECT 63.180 120.215 63.350 120.725 ;
        RECT 63.520 120.465 64.040 120.775 ;
        RECT 61.450 120.045 63.350 120.215 ;
        RECT 61.450 119.985 61.780 120.045 ;
        RECT 61.930 119.815 62.260 119.875 ;
        RECT 61.600 119.545 62.260 119.815 ;
        RECT 61.090 119.160 61.410 119.490 ;
        RECT 62.450 119.285 62.620 120.045 ;
        RECT 63.520 119.875 63.700 120.285 ;
        RECT 62.790 119.705 63.120 119.825 ;
        RECT 63.870 119.705 64.040 120.465 ;
        RECT 62.790 119.535 64.040 119.705 ;
        RECT 64.210 120.645 65.580 120.895 ;
        RECT 64.210 119.875 64.400 120.645 ;
        RECT 65.330 120.385 65.580 120.645 ;
        RECT 64.570 120.215 64.820 120.375 ;
        RECT 65.750 120.215 65.920 121.060 ;
        RECT 66.815 120.775 66.985 121.275 ;
        RECT 66.090 120.385 66.590 120.765 ;
        RECT 66.815 120.605 67.510 120.775 ;
        RECT 64.570 120.045 65.920 120.215 ;
        RECT 65.500 120.005 65.920 120.045 ;
        RECT 64.210 119.535 64.630 119.875 ;
        RECT 64.920 119.545 65.330 119.875 ;
        RECT 62.450 119.115 63.300 119.285 ;
        RECT 64.380 119.105 64.630 119.535 ;
        RECT 65.500 119.275 65.670 120.005 ;
        RECT 65.840 119.455 66.190 119.825 ;
        RECT 66.370 119.515 66.590 120.385 ;
        RECT 66.760 119.815 67.170 120.435 ;
        RECT 67.340 119.635 67.510 120.605 ;
        RECT 66.815 119.445 67.510 119.635 ;
        RECT 65.500 119.075 66.515 119.275 ;
        RECT 66.815 119.115 66.985 119.445 ;
        RECT 67.700 119.155 67.925 121.275 ;
        RECT 68.595 120.775 68.765 121.275 ;
        RECT 68.100 120.605 68.765 120.775 ;
        RECT 68.100 119.615 68.330 120.605 ;
        RECT 68.500 119.785 68.850 120.435 ;
        RECT 69.025 120.370 69.295 121.275 ;
        RECT 69.975 120.515 70.145 121.275 ;
        RECT 68.100 119.445 68.765 119.615 ;
        RECT 68.595 119.155 68.765 119.445 ;
        RECT 69.025 119.570 69.195 120.370 ;
        RECT 69.480 120.345 70.145 120.515 ;
        RECT 69.480 120.200 69.650 120.345 ;
        RECT 74.985 120.295 75.315 121.275 ;
        RECT 77.935 121.105 79.965 121.275 ;
        RECT 69.365 119.870 69.650 120.200 ;
        RECT 69.480 119.615 69.650 119.870 ;
        RECT 69.885 119.795 70.215 120.165 ;
        RECT 74.565 119.885 74.895 120.135 ;
        RECT 75.065 119.695 75.315 120.295 ;
        RECT 76.845 120.685 77.360 121.095 ;
        RECT 76.845 119.875 77.185 120.685 ;
        RECT 77.935 120.440 78.105 121.105 ;
        RECT 78.500 120.765 79.625 120.935 ;
        RECT 77.355 120.250 78.105 120.440 ;
        RECT 78.275 120.425 79.285 120.595 ;
        RECT 76.845 119.705 78.075 119.875 ;
        RECT 69.025 119.065 69.285 119.570 ;
        RECT 69.480 119.445 70.145 119.615 ;
        RECT 69.975 119.065 70.145 119.445 ;
        RECT 74.985 119.065 75.315 119.695 ;
        RECT 77.120 119.100 77.365 119.705 ;
        RECT 78.275 119.065 78.465 120.425 ;
        RECT 78.635 119.405 78.910 120.225 ;
        RECT 79.115 119.625 79.285 120.425 ;
        RECT 79.455 119.635 79.625 120.765 ;
        RECT 79.795 120.135 79.965 121.105 ;
        RECT 80.475 120.305 80.810 121.275 ;
        RECT 79.795 119.805 79.990 120.135 ;
        RECT 80.215 119.805 80.470 120.135 ;
        RECT 80.215 119.635 80.385 119.805 ;
        RECT 80.640 119.635 80.810 120.305 ;
        RECT 79.455 119.465 80.385 119.635 ;
        RECT 79.455 119.430 79.630 119.465 ;
        RECT 78.635 119.235 78.915 119.405 ;
        RECT 78.635 119.065 78.910 119.235 ;
        RECT 79.100 119.065 79.630 119.430 ;
        RECT 80.555 119.065 80.810 119.635 ;
        RECT 80.985 120.370 81.255 121.275 ;
        RECT 81.935 120.515 82.105 121.275 ;
        RECT 80.985 119.570 81.155 120.370 ;
        RECT 81.440 120.345 82.105 120.515 ;
        RECT 81.440 120.200 81.610 120.345 ;
        RECT 81.325 119.870 81.610 120.200 ;
        RECT 82.805 120.295 83.135 121.275 ;
        RECT 84.295 120.515 84.465 121.275 ;
        RECT 84.295 120.345 84.960 120.515 ;
        RECT 85.145 120.370 85.415 121.275 ;
        RECT 81.440 119.615 81.610 119.870 ;
        RECT 81.845 119.795 82.175 120.165 ;
        RECT 82.805 119.695 83.055 120.295 ;
        RECT 84.790 120.200 84.960 120.345 ;
        RECT 83.225 119.885 83.555 120.135 ;
        RECT 84.225 119.795 84.555 120.165 ;
        RECT 84.790 119.870 85.075 120.200 ;
        RECT 80.985 119.065 81.245 119.570 ;
        RECT 81.440 119.445 82.105 119.615 ;
        RECT 81.935 119.065 82.105 119.445 ;
        RECT 82.805 119.065 83.135 119.695 ;
        RECT 84.790 119.615 84.960 119.870 ;
        RECT 84.295 119.445 84.960 119.615 ;
        RECT 85.245 119.570 85.415 120.370 ;
        RECT 89.705 120.295 90.035 121.275 ;
        RECT 91.085 120.295 91.415 121.275 ;
        RECT 92.400 120.465 92.655 121.135 ;
        RECT 93.300 120.725 93.630 121.235 ;
        RECT 92.400 120.425 92.580 120.465 ;
        RECT 89.285 119.885 89.615 120.135 ;
        RECT 89.785 119.695 90.035 120.295 ;
        RECT 90.665 119.885 90.995 120.135 ;
        RECT 91.165 119.695 91.415 120.295 ;
        RECT 92.315 120.255 92.580 120.425 ;
        RECT 84.295 119.065 84.465 119.445 ;
        RECT 85.155 119.065 85.415 119.570 ;
        RECT 89.705 119.065 90.035 119.695 ;
        RECT 91.085 119.065 91.415 119.695 ;
        RECT 92.400 119.605 92.580 120.255 ;
        RECT 93.300 120.135 93.550 120.725 ;
        RECT 93.900 120.575 94.070 121.185 ;
        RECT 94.800 120.895 95.040 121.185 ;
        RECT 95.840 120.975 96.470 121.225 ;
        RECT 95.840 120.895 96.010 120.975 ;
        RECT 97.440 120.895 97.610 121.185 ;
        RECT 98.410 121.060 99.240 121.230 ;
        RECT 94.800 120.725 96.010 120.895 ;
        RECT 92.750 119.805 93.550 120.135 ;
        RECT 92.400 119.075 92.655 119.605 ;
        RECT 93.300 119.155 93.550 119.805 ;
        RECT 93.750 120.555 94.070 120.575 ;
        RECT 93.750 120.385 95.670 120.555 ;
        RECT 93.750 119.490 93.940 120.385 ;
        RECT 95.840 120.215 96.010 120.725 ;
        RECT 96.180 120.465 96.700 120.775 ;
        RECT 94.110 120.045 96.010 120.215 ;
        RECT 94.110 119.985 94.440 120.045 ;
        RECT 94.590 119.815 94.920 119.875 ;
        RECT 94.260 119.545 94.920 119.815 ;
        RECT 93.750 119.160 94.070 119.490 ;
        RECT 95.110 119.285 95.280 120.045 ;
        RECT 96.180 119.875 96.360 120.285 ;
        RECT 95.450 119.705 95.780 119.825 ;
        RECT 96.530 119.705 96.700 120.465 ;
        RECT 95.450 119.535 96.700 119.705 ;
        RECT 96.870 120.645 98.240 120.895 ;
        RECT 96.870 119.875 97.060 120.645 ;
        RECT 97.990 120.385 98.240 120.645 ;
        RECT 97.230 120.215 97.480 120.375 ;
        RECT 98.410 120.215 98.580 121.060 ;
        RECT 99.475 120.775 99.645 121.275 ;
        RECT 98.750 120.385 99.250 120.765 ;
        RECT 99.475 120.605 100.170 120.775 ;
        RECT 97.230 120.045 98.580 120.215 ;
        RECT 98.160 120.005 98.580 120.045 ;
        RECT 96.870 119.535 97.290 119.875 ;
        RECT 97.580 119.545 97.990 119.875 ;
        RECT 95.110 119.115 95.960 119.285 ;
        RECT 97.040 119.105 97.290 119.535 ;
        RECT 98.160 119.275 98.330 120.005 ;
        RECT 98.500 119.455 98.850 119.825 ;
        RECT 99.030 119.515 99.250 120.385 ;
        RECT 99.420 119.815 99.830 120.435 ;
        RECT 100.000 119.635 100.170 120.605 ;
        RECT 99.475 119.445 100.170 119.635 ;
        RECT 98.160 119.075 99.175 119.275 ;
        RECT 99.475 119.115 99.645 119.445 ;
        RECT 100.360 119.155 100.585 121.275 ;
        RECT 101.255 120.775 101.425 121.275 ;
        RECT 100.760 120.605 101.425 120.775 ;
        RECT 100.760 119.615 100.990 120.605 ;
        RECT 101.160 119.785 101.510 120.435 ;
        RECT 102.145 120.370 102.415 121.275 ;
        RECT 103.095 120.515 103.265 121.275 ;
        RECT 100.760 119.445 101.425 119.615 ;
        RECT 101.255 119.155 101.425 119.445 ;
        RECT 102.145 119.570 102.315 120.370 ;
        RECT 102.600 120.345 103.265 120.515 ;
        RECT 102.600 120.200 102.770 120.345 ;
        RECT 103.965 120.295 104.295 121.275 ;
        RECT 105.995 121.105 108.025 121.275 ;
        RECT 102.485 119.870 102.770 120.200 ;
        RECT 102.600 119.615 102.770 119.870 ;
        RECT 103.005 119.795 103.335 120.165 ;
        RECT 103.545 119.885 103.875 120.135 ;
        RECT 104.045 119.695 104.295 120.295 ;
        RECT 104.905 120.685 105.420 121.095 ;
        RECT 104.905 119.875 105.245 120.685 ;
        RECT 105.995 120.440 106.165 121.105 ;
        RECT 106.560 120.765 107.685 120.935 ;
        RECT 105.415 120.250 106.165 120.440 ;
        RECT 106.335 120.425 107.345 120.595 ;
        RECT 104.905 119.705 106.135 119.875 ;
        RECT 102.145 119.065 102.405 119.570 ;
        RECT 102.600 119.445 103.265 119.615 ;
        RECT 103.095 119.065 103.265 119.445 ;
        RECT 103.965 119.065 104.295 119.695 ;
        RECT 105.180 119.100 105.425 119.705 ;
        RECT 106.335 119.065 106.525 120.425 ;
        RECT 106.695 120.085 106.970 120.225 ;
        RECT 106.695 119.915 106.975 120.085 ;
        RECT 106.695 119.065 106.970 119.915 ;
        RECT 107.175 119.625 107.345 120.425 ;
        RECT 107.515 119.635 107.685 120.765 ;
        RECT 107.855 120.135 108.025 121.105 ;
        RECT 108.535 120.305 108.870 121.275 ;
        RECT 107.855 119.805 108.050 120.135 ;
        RECT 108.275 119.805 108.530 120.135 ;
        RECT 108.275 119.635 108.445 119.805 ;
        RECT 108.700 119.635 108.870 120.305 ;
        RECT 109.420 120.465 109.675 121.135 ;
        RECT 110.320 120.725 110.650 121.235 ;
        RECT 109.420 119.745 109.600 120.465 ;
        RECT 110.320 120.135 110.570 120.725 ;
        RECT 110.920 120.575 111.090 121.185 ;
        RECT 111.820 120.895 112.060 121.185 ;
        RECT 112.860 120.975 113.490 121.225 ;
        RECT 112.860 120.895 113.030 120.975 ;
        RECT 114.460 120.895 114.630 121.185 ;
        RECT 115.430 121.060 116.260 121.230 ;
        RECT 111.820 120.725 113.030 120.895 ;
        RECT 109.770 119.805 110.570 120.135 ;
        RECT 107.515 119.465 108.445 119.635 ;
        RECT 107.515 119.430 107.690 119.465 ;
        RECT 107.160 119.065 107.690 119.430 ;
        RECT 108.615 119.065 108.870 119.635 ;
        RECT 109.335 119.605 109.600 119.745 ;
        RECT 109.335 119.575 109.675 119.605 ;
        RECT 109.420 119.075 109.675 119.575 ;
        RECT 110.320 119.155 110.570 119.805 ;
        RECT 110.770 120.555 111.090 120.575 ;
        RECT 110.770 120.385 112.690 120.555 ;
        RECT 110.770 119.490 110.960 120.385 ;
        RECT 112.860 120.215 113.030 120.725 ;
        RECT 113.200 120.465 113.720 120.775 ;
        RECT 111.130 120.045 113.030 120.215 ;
        RECT 111.130 119.985 111.460 120.045 ;
        RECT 111.610 119.815 111.940 119.875 ;
        RECT 111.280 119.545 111.940 119.815 ;
        RECT 110.770 119.160 111.090 119.490 ;
        RECT 112.130 119.285 112.300 120.045 ;
        RECT 113.200 119.875 113.380 120.285 ;
        RECT 112.470 119.705 112.800 119.825 ;
        RECT 113.550 119.705 113.720 120.465 ;
        RECT 112.470 119.535 113.720 119.705 ;
        RECT 113.890 120.645 115.260 120.895 ;
        RECT 113.890 119.875 114.080 120.645 ;
        RECT 115.010 120.385 115.260 120.645 ;
        RECT 114.250 120.215 114.500 120.375 ;
        RECT 115.430 120.215 115.600 121.060 ;
        RECT 116.495 120.775 116.665 121.275 ;
        RECT 115.770 120.385 116.270 120.765 ;
        RECT 116.495 120.605 117.190 120.775 ;
        RECT 114.250 120.045 115.600 120.215 ;
        RECT 115.180 120.005 115.600 120.045 ;
        RECT 113.890 119.535 114.310 119.875 ;
        RECT 114.600 119.545 115.010 119.875 ;
        RECT 112.130 119.115 112.980 119.285 ;
        RECT 114.060 119.105 114.310 119.535 ;
        RECT 115.180 119.275 115.350 120.005 ;
        RECT 115.520 119.455 115.870 119.825 ;
        RECT 116.050 119.515 116.270 120.385 ;
        RECT 116.440 119.815 116.850 120.435 ;
        RECT 117.020 119.635 117.190 120.605 ;
        RECT 116.495 119.445 117.190 119.635 ;
        RECT 115.180 119.075 116.195 119.275 ;
        RECT 116.495 119.115 116.665 119.445 ;
        RECT 117.380 119.155 117.605 121.275 ;
        RECT 118.275 120.775 118.445 121.275 ;
        RECT 117.780 120.605 118.445 120.775 ;
        RECT 117.780 119.615 118.010 120.605 ;
        RECT 118.180 119.785 118.530 120.435 ;
        RECT 119.145 120.295 119.475 121.275 ;
        RECT 120.635 120.515 120.805 121.275 ;
        RECT 120.635 120.345 121.300 120.515 ;
        RECT 121.485 120.370 121.755 121.275 ;
        RECT 118.725 119.885 119.055 120.135 ;
        RECT 119.225 119.695 119.475 120.295 ;
        RECT 121.130 120.200 121.300 120.345 ;
        RECT 120.565 119.795 120.895 120.165 ;
        RECT 121.130 119.870 121.415 120.200 ;
        RECT 117.780 119.445 118.445 119.615 ;
        RECT 118.275 119.155 118.445 119.445 ;
        RECT 119.145 119.065 119.475 119.695 ;
        RECT 121.130 119.615 121.300 119.870 ;
        RECT 120.635 119.445 121.300 119.615 ;
        RECT 121.585 119.570 121.755 120.370 ;
        RECT 120.635 119.065 120.805 119.445 ;
        RECT 121.495 119.065 121.755 119.570 ;
        RECT 18.340 118.385 18.595 118.545 ;
        RECT 18.255 118.215 18.595 118.385 ;
        RECT 18.340 118.015 18.595 118.215 ;
        RECT 18.340 117.155 18.520 118.015 ;
        RECT 19.240 117.815 19.490 118.465 ;
        RECT 18.690 117.485 19.490 117.815 ;
        RECT 18.340 116.485 18.595 117.155 ;
        RECT 19.240 116.895 19.490 117.485 ;
        RECT 19.690 118.130 20.010 118.460 ;
        RECT 21.050 118.335 21.900 118.505 ;
        RECT 19.690 117.235 19.880 118.130 ;
        RECT 20.200 117.805 20.860 118.075 ;
        RECT 20.530 117.745 20.860 117.805 ;
        RECT 20.050 117.575 20.380 117.635 ;
        RECT 21.050 117.575 21.220 118.335 ;
        RECT 22.980 118.085 23.230 118.515 ;
        RECT 21.390 117.915 22.640 118.085 ;
        RECT 21.390 117.795 21.720 117.915 ;
        RECT 20.050 117.405 21.950 117.575 ;
        RECT 19.690 117.065 21.610 117.235 ;
        RECT 19.690 117.045 20.010 117.065 ;
        RECT 19.240 116.385 19.570 116.895 ;
        RECT 19.840 116.435 20.010 117.045 ;
        RECT 21.780 116.895 21.950 117.405 ;
        RECT 22.120 117.335 22.300 117.745 ;
        RECT 22.470 117.155 22.640 117.915 ;
        RECT 20.740 116.725 21.950 116.895 ;
        RECT 22.120 116.845 22.640 117.155 ;
        RECT 22.810 117.745 23.230 118.085 ;
        RECT 24.100 118.345 25.115 118.545 ;
        RECT 23.520 117.745 23.930 118.075 ;
        RECT 22.810 116.975 23.000 117.745 ;
        RECT 24.100 117.615 24.270 118.345 ;
        RECT 25.415 118.175 25.585 118.505 ;
        RECT 24.440 117.795 24.790 118.165 ;
        RECT 24.100 117.575 24.520 117.615 ;
        RECT 23.170 117.405 24.520 117.575 ;
        RECT 23.170 117.245 23.420 117.405 ;
        RECT 23.930 116.975 24.180 117.235 ;
        RECT 22.810 116.725 24.180 116.975 ;
        RECT 20.740 116.435 20.980 116.725 ;
        RECT 21.780 116.645 21.950 116.725 ;
        RECT 21.780 116.395 22.410 116.645 ;
        RECT 23.380 116.435 23.550 116.725 ;
        RECT 24.350 116.560 24.520 117.405 ;
        RECT 24.970 117.235 25.190 118.105 ;
        RECT 25.415 117.985 26.110 118.175 ;
        RECT 24.690 116.855 25.190 117.235 ;
        RECT 25.360 117.185 25.770 117.805 ;
        RECT 25.940 117.015 26.110 117.985 ;
        RECT 25.415 116.845 26.110 117.015 ;
        RECT 24.350 116.390 25.180 116.560 ;
        RECT 25.415 116.345 25.585 116.845 ;
        RECT 26.300 116.345 26.525 118.465 ;
        RECT 27.195 118.175 27.365 118.465 ;
        RECT 28.000 118.385 28.255 118.545 ;
        RECT 27.915 118.215 28.255 118.385 ;
        RECT 26.700 118.005 27.365 118.175 ;
        RECT 28.000 118.015 28.255 118.215 ;
        RECT 26.700 117.015 26.930 118.005 ;
        RECT 27.100 117.185 27.450 117.835 ;
        RECT 28.000 117.155 28.180 118.015 ;
        RECT 28.900 117.815 29.150 118.465 ;
        RECT 28.350 117.485 29.150 117.815 ;
        RECT 26.700 116.845 27.365 117.015 ;
        RECT 27.195 116.345 27.365 116.845 ;
        RECT 28.000 116.485 28.255 117.155 ;
        RECT 28.900 116.895 29.150 117.485 ;
        RECT 29.350 118.130 29.670 118.460 ;
        RECT 30.710 118.335 31.560 118.505 ;
        RECT 29.350 117.235 29.540 118.130 ;
        RECT 29.860 117.805 30.520 118.075 ;
        RECT 30.190 117.745 30.520 117.805 ;
        RECT 29.710 117.575 30.040 117.635 ;
        RECT 30.710 117.575 30.880 118.335 ;
        RECT 32.640 118.085 32.890 118.515 ;
        RECT 31.050 117.915 32.300 118.085 ;
        RECT 31.050 117.795 31.380 117.915 ;
        RECT 29.710 117.405 31.610 117.575 ;
        RECT 29.350 117.065 31.270 117.235 ;
        RECT 29.350 117.045 29.670 117.065 ;
        RECT 28.900 116.385 29.230 116.895 ;
        RECT 29.500 116.435 29.670 117.045 ;
        RECT 31.440 116.895 31.610 117.405 ;
        RECT 31.780 117.335 31.960 117.745 ;
        RECT 32.130 117.155 32.300 117.915 ;
        RECT 30.400 116.725 31.610 116.895 ;
        RECT 31.780 116.845 32.300 117.155 ;
        RECT 32.470 117.745 32.890 118.085 ;
        RECT 33.760 118.345 34.775 118.545 ;
        RECT 33.180 117.745 33.590 118.075 ;
        RECT 32.470 116.975 32.660 117.745 ;
        RECT 33.760 117.615 33.930 118.345 ;
        RECT 35.075 118.175 35.245 118.505 ;
        RECT 34.100 117.795 34.450 118.165 ;
        RECT 33.760 117.575 34.180 117.615 ;
        RECT 32.830 117.405 34.180 117.575 ;
        RECT 32.830 117.245 33.080 117.405 ;
        RECT 33.590 116.975 33.840 117.235 ;
        RECT 32.470 116.725 33.840 116.975 ;
        RECT 30.400 116.435 30.640 116.725 ;
        RECT 31.440 116.645 31.610 116.725 ;
        RECT 31.440 116.395 32.070 116.645 ;
        RECT 33.040 116.435 33.210 116.725 ;
        RECT 34.010 116.560 34.180 117.405 ;
        RECT 34.630 117.235 34.850 118.105 ;
        RECT 35.075 117.985 35.770 118.175 ;
        RECT 34.350 116.855 34.850 117.235 ;
        RECT 35.020 117.185 35.430 117.805 ;
        RECT 35.600 117.015 35.770 117.985 ;
        RECT 35.075 116.845 35.770 117.015 ;
        RECT 34.010 116.390 34.840 116.560 ;
        RECT 35.075 116.345 35.245 116.845 ;
        RECT 35.960 116.345 36.185 118.465 ;
        RECT 36.855 118.175 37.025 118.465 ;
        RECT 38.120 118.385 38.375 118.545 ;
        RECT 38.035 118.215 38.375 118.385 ;
        RECT 36.360 118.005 37.025 118.175 ;
        RECT 38.120 118.015 38.375 118.215 ;
        RECT 36.360 117.015 36.590 118.005 ;
        RECT 36.760 117.185 37.110 117.835 ;
        RECT 38.120 117.155 38.300 118.015 ;
        RECT 39.020 117.815 39.270 118.465 ;
        RECT 38.470 117.485 39.270 117.815 ;
        RECT 36.360 116.845 37.025 117.015 ;
        RECT 36.855 116.345 37.025 116.845 ;
        RECT 38.120 116.485 38.375 117.155 ;
        RECT 39.020 116.895 39.270 117.485 ;
        RECT 39.470 118.130 39.790 118.460 ;
        RECT 40.830 118.335 41.680 118.505 ;
        RECT 39.470 117.235 39.660 118.130 ;
        RECT 39.980 117.805 40.640 118.075 ;
        RECT 40.310 117.745 40.640 117.805 ;
        RECT 39.830 117.575 40.160 117.635 ;
        RECT 40.830 117.575 41.000 118.335 ;
        RECT 42.760 118.085 43.010 118.515 ;
        RECT 41.170 117.915 42.420 118.085 ;
        RECT 41.170 117.795 41.500 117.915 ;
        RECT 39.830 117.405 41.730 117.575 ;
        RECT 39.470 117.065 41.390 117.235 ;
        RECT 39.470 117.045 39.790 117.065 ;
        RECT 39.020 116.385 39.350 116.895 ;
        RECT 39.620 116.435 39.790 117.045 ;
        RECT 41.560 116.895 41.730 117.405 ;
        RECT 41.900 117.335 42.080 117.745 ;
        RECT 42.250 117.155 42.420 117.915 ;
        RECT 40.520 116.725 41.730 116.895 ;
        RECT 41.900 116.845 42.420 117.155 ;
        RECT 42.590 117.745 43.010 118.085 ;
        RECT 43.880 118.345 44.895 118.545 ;
        RECT 43.300 117.745 43.710 118.075 ;
        RECT 42.590 116.975 42.780 117.745 ;
        RECT 43.880 117.615 44.050 118.345 ;
        RECT 45.195 118.175 45.365 118.505 ;
        RECT 44.220 117.795 44.570 118.165 ;
        RECT 43.880 117.575 44.300 117.615 ;
        RECT 42.950 117.405 44.300 117.575 ;
        RECT 42.950 117.245 43.200 117.405 ;
        RECT 43.710 116.975 43.960 117.235 ;
        RECT 42.590 116.725 43.960 116.975 ;
        RECT 40.520 116.435 40.760 116.725 ;
        RECT 41.560 116.645 41.730 116.725 ;
        RECT 41.560 116.395 42.190 116.645 ;
        RECT 43.160 116.435 43.330 116.725 ;
        RECT 44.130 116.560 44.300 117.405 ;
        RECT 44.750 117.235 44.970 118.105 ;
        RECT 45.195 117.985 45.890 118.175 ;
        RECT 44.470 116.855 44.970 117.235 ;
        RECT 45.140 117.185 45.550 117.805 ;
        RECT 45.720 117.015 45.890 117.985 ;
        RECT 45.195 116.845 45.890 117.015 ;
        RECT 44.130 116.390 44.960 116.560 ;
        RECT 45.195 116.345 45.365 116.845 ;
        RECT 46.080 116.345 46.305 118.465 ;
        RECT 46.975 118.175 47.145 118.465 ;
        RECT 47.780 118.385 48.035 118.545 ;
        RECT 47.695 118.215 48.035 118.385 ;
        RECT 46.480 118.005 47.145 118.175 ;
        RECT 47.780 118.015 48.035 118.215 ;
        RECT 46.480 117.015 46.710 118.005 ;
        RECT 46.880 117.185 47.230 117.835 ;
        RECT 47.780 117.155 47.960 118.015 ;
        RECT 48.680 117.815 48.930 118.465 ;
        RECT 48.130 117.485 48.930 117.815 ;
        RECT 46.480 116.845 47.145 117.015 ;
        RECT 46.975 116.345 47.145 116.845 ;
        RECT 47.780 116.485 48.035 117.155 ;
        RECT 48.680 116.895 48.930 117.485 ;
        RECT 49.130 118.130 49.450 118.460 ;
        RECT 50.490 118.335 51.340 118.505 ;
        RECT 49.130 117.235 49.320 118.130 ;
        RECT 49.640 117.805 50.300 118.075 ;
        RECT 49.970 117.745 50.300 117.805 ;
        RECT 49.490 117.575 49.820 117.635 ;
        RECT 50.490 117.575 50.660 118.335 ;
        RECT 52.420 118.085 52.670 118.515 ;
        RECT 50.830 117.915 52.080 118.085 ;
        RECT 50.830 117.795 51.160 117.915 ;
        RECT 49.490 117.405 51.390 117.575 ;
        RECT 49.130 117.065 51.050 117.235 ;
        RECT 49.130 117.045 49.450 117.065 ;
        RECT 48.680 116.385 49.010 116.895 ;
        RECT 49.280 116.435 49.450 117.045 ;
        RECT 51.220 116.895 51.390 117.405 ;
        RECT 51.560 117.335 51.740 117.745 ;
        RECT 51.910 117.155 52.080 117.915 ;
        RECT 50.180 116.725 51.390 116.895 ;
        RECT 51.560 116.845 52.080 117.155 ;
        RECT 52.250 117.745 52.670 118.085 ;
        RECT 53.540 118.345 54.555 118.545 ;
        RECT 52.960 117.745 53.370 118.075 ;
        RECT 52.250 116.975 52.440 117.745 ;
        RECT 53.540 117.615 53.710 118.345 ;
        RECT 54.855 118.175 55.025 118.505 ;
        RECT 53.880 117.795 54.230 118.165 ;
        RECT 53.540 117.575 53.960 117.615 ;
        RECT 52.610 117.405 53.960 117.575 ;
        RECT 52.610 117.245 52.860 117.405 ;
        RECT 53.370 116.975 53.620 117.235 ;
        RECT 52.250 116.725 53.620 116.975 ;
        RECT 50.180 116.435 50.420 116.725 ;
        RECT 51.220 116.645 51.390 116.725 ;
        RECT 51.220 116.395 51.850 116.645 ;
        RECT 52.820 116.435 52.990 116.725 ;
        RECT 53.790 116.560 53.960 117.405 ;
        RECT 54.410 117.235 54.630 118.105 ;
        RECT 54.855 117.985 55.550 118.175 ;
        RECT 54.130 116.855 54.630 117.235 ;
        RECT 54.800 117.185 55.210 117.805 ;
        RECT 55.380 117.015 55.550 117.985 ;
        RECT 54.855 116.845 55.550 117.015 ;
        RECT 53.790 116.390 54.620 116.560 ;
        RECT 54.855 116.345 55.025 116.845 ;
        RECT 55.740 116.345 55.965 118.465 ;
        RECT 56.635 118.175 56.805 118.465 ;
        RECT 56.140 118.005 56.805 118.175 ;
        RECT 56.140 117.015 56.370 118.005 ;
        RECT 57.505 117.925 57.835 118.555 ;
        RECT 62.105 117.925 62.435 118.555 ;
        RECT 63.880 118.385 64.135 118.545 ;
        RECT 63.795 118.215 64.135 118.385 ;
        RECT 56.540 117.185 56.890 117.835 ;
        RECT 57.505 117.325 57.755 117.925 ;
        RECT 57.925 117.485 58.255 117.735 ;
        RECT 61.685 117.485 62.015 117.735 ;
        RECT 62.185 117.325 62.435 117.925 ;
        RECT 56.140 116.845 56.805 117.015 ;
        RECT 56.635 116.345 56.805 116.845 ;
        RECT 57.505 116.345 57.835 117.325 ;
        RECT 62.105 116.345 62.435 117.325 ;
        RECT 63.880 118.015 64.135 118.215 ;
        RECT 63.880 117.155 64.060 118.015 ;
        RECT 64.780 117.815 65.030 118.465 ;
        RECT 64.230 117.485 65.030 117.815 ;
        RECT 63.880 116.485 64.135 117.155 ;
        RECT 64.780 116.895 65.030 117.485 ;
        RECT 65.230 118.130 65.550 118.460 ;
        RECT 66.590 118.335 67.440 118.505 ;
        RECT 65.230 117.235 65.420 118.130 ;
        RECT 65.740 117.805 66.400 118.075 ;
        RECT 66.070 117.745 66.400 117.805 ;
        RECT 65.590 117.575 65.920 117.635 ;
        RECT 66.590 117.575 66.760 118.335 ;
        RECT 68.520 118.085 68.770 118.515 ;
        RECT 66.930 117.915 68.180 118.085 ;
        RECT 66.930 117.795 67.260 117.915 ;
        RECT 65.590 117.405 67.490 117.575 ;
        RECT 65.230 117.065 67.150 117.235 ;
        RECT 65.230 117.045 65.550 117.065 ;
        RECT 64.780 116.385 65.110 116.895 ;
        RECT 65.380 116.435 65.550 117.045 ;
        RECT 67.320 116.895 67.490 117.405 ;
        RECT 67.660 117.335 67.840 117.745 ;
        RECT 68.010 117.155 68.180 117.915 ;
        RECT 66.280 116.725 67.490 116.895 ;
        RECT 67.660 116.845 68.180 117.155 ;
        RECT 68.350 117.745 68.770 118.085 ;
        RECT 69.640 118.345 70.655 118.545 ;
        RECT 69.060 117.745 69.470 118.075 ;
        RECT 68.350 116.975 68.540 117.745 ;
        RECT 69.640 117.615 69.810 118.345 ;
        RECT 70.955 118.175 71.125 118.505 ;
        RECT 69.980 117.795 70.330 118.165 ;
        RECT 69.640 117.575 70.060 117.615 ;
        RECT 68.710 117.405 70.060 117.575 ;
        RECT 68.710 117.245 68.960 117.405 ;
        RECT 69.470 116.975 69.720 117.235 ;
        RECT 68.350 116.725 69.720 116.975 ;
        RECT 66.280 116.435 66.520 116.725 ;
        RECT 67.320 116.645 67.490 116.725 ;
        RECT 67.320 116.395 67.950 116.645 ;
        RECT 68.920 116.435 69.090 116.725 ;
        RECT 69.890 116.560 70.060 117.405 ;
        RECT 70.510 117.235 70.730 118.105 ;
        RECT 70.955 117.985 71.650 118.175 ;
        RECT 70.230 116.855 70.730 117.235 ;
        RECT 70.900 117.185 71.310 117.805 ;
        RECT 71.480 117.015 71.650 117.985 ;
        RECT 70.955 116.845 71.650 117.015 ;
        RECT 69.890 116.390 70.720 116.560 ;
        RECT 70.955 116.345 71.125 116.845 ;
        RECT 71.840 116.345 72.065 118.465 ;
        RECT 72.735 118.175 72.905 118.465 ;
        RECT 73.540 118.385 73.795 118.545 ;
        RECT 73.455 118.215 73.795 118.385 ;
        RECT 72.240 118.005 72.905 118.175 ;
        RECT 73.540 118.015 73.795 118.215 ;
        RECT 72.240 117.015 72.470 118.005 ;
        RECT 72.640 117.185 72.990 117.835 ;
        RECT 73.540 117.155 73.720 118.015 ;
        RECT 74.440 117.815 74.690 118.465 ;
        RECT 73.890 117.485 74.690 117.815 ;
        RECT 72.240 116.845 72.905 117.015 ;
        RECT 72.735 116.345 72.905 116.845 ;
        RECT 73.540 116.485 73.795 117.155 ;
        RECT 74.440 116.895 74.690 117.485 ;
        RECT 74.890 118.130 75.210 118.460 ;
        RECT 76.250 118.335 77.100 118.505 ;
        RECT 74.890 117.235 75.080 118.130 ;
        RECT 75.400 117.805 76.060 118.075 ;
        RECT 75.730 117.745 76.060 117.805 ;
        RECT 75.250 117.575 75.580 117.635 ;
        RECT 76.250 117.575 76.420 118.335 ;
        RECT 78.180 118.085 78.430 118.515 ;
        RECT 76.590 117.915 77.840 118.085 ;
        RECT 76.590 117.795 76.920 117.915 ;
        RECT 75.250 117.405 77.150 117.575 ;
        RECT 74.890 117.065 76.810 117.235 ;
        RECT 74.890 117.045 75.210 117.065 ;
        RECT 74.440 116.385 74.770 116.895 ;
        RECT 75.040 116.435 75.210 117.045 ;
        RECT 76.980 116.895 77.150 117.405 ;
        RECT 77.320 117.335 77.500 117.745 ;
        RECT 77.670 117.155 77.840 117.915 ;
        RECT 75.940 116.725 77.150 116.895 ;
        RECT 77.320 116.845 77.840 117.155 ;
        RECT 78.010 117.745 78.430 118.085 ;
        RECT 79.300 118.345 80.315 118.545 ;
        RECT 78.720 117.745 79.130 118.075 ;
        RECT 78.010 116.975 78.200 117.745 ;
        RECT 79.300 117.615 79.470 118.345 ;
        RECT 80.615 118.175 80.785 118.505 ;
        RECT 79.640 117.795 79.990 118.165 ;
        RECT 79.300 117.575 79.720 117.615 ;
        RECT 78.370 117.405 79.720 117.575 ;
        RECT 78.370 117.245 78.620 117.405 ;
        RECT 79.130 116.975 79.380 117.235 ;
        RECT 78.010 116.725 79.380 116.975 ;
        RECT 75.940 116.435 76.180 116.725 ;
        RECT 76.980 116.645 77.150 116.725 ;
        RECT 76.980 116.395 77.610 116.645 ;
        RECT 78.580 116.435 78.750 116.725 ;
        RECT 79.550 116.560 79.720 117.405 ;
        RECT 80.170 117.235 80.390 118.105 ;
        RECT 80.615 117.985 81.310 118.175 ;
        RECT 79.890 116.855 80.390 117.235 ;
        RECT 80.560 117.185 80.970 117.805 ;
        RECT 81.140 117.015 81.310 117.985 ;
        RECT 80.615 116.845 81.310 117.015 ;
        RECT 79.550 116.390 80.380 116.560 ;
        RECT 80.615 116.345 80.785 116.845 ;
        RECT 81.500 116.345 81.725 118.465 ;
        RECT 82.395 118.175 82.565 118.465 ;
        RECT 81.900 118.005 82.565 118.175 ;
        RECT 81.900 117.015 82.130 118.005 ;
        RECT 82.830 117.985 83.085 118.555 ;
        RECT 84.010 118.190 84.540 118.555 ;
        RECT 84.010 118.155 84.185 118.190 ;
        RECT 83.255 117.985 84.185 118.155 ;
        RECT 84.730 118.045 85.005 118.555 ;
        RECT 82.300 117.185 82.650 117.835 ;
        RECT 82.830 117.315 83.000 117.985 ;
        RECT 83.255 117.815 83.425 117.985 ;
        RECT 83.170 117.485 83.425 117.815 ;
        RECT 83.650 117.485 83.845 117.815 ;
        RECT 81.900 116.845 82.565 117.015 ;
        RECT 82.395 116.345 82.565 116.845 ;
        RECT 82.830 116.345 83.165 117.315 ;
        RECT 83.675 116.515 83.845 117.485 ;
        RECT 84.015 116.855 84.185 117.985 ;
        RECT 84.355 117.195 84.525 117.995 ;
        RECT 84.725 117.875 85.005 118.045 ;
        RECT 84.730 117.395 85.005 117.875 ;
        RECT 85.175 117.195 85.365 118.555 ;
        RECT 86.275 117.915 86.520 118.520 ;
        RECT 87.865 117.925 88.195 118.555 ;
        RECT 89.640 118.385 89.895 118.545 ;
        RECT 89.555 118.215 89.895 118.385 ;
        RECT 85.565 117.745 86.795 117.915 ;
        RECT 84.355 117.025 85.365 117.195 ;
        RECT 85.535 117.180 86.285 117.370 ;
        RECT 84.015 116.685 85.140 116.855 ;
        RECT 85.535 116.515 85.705 117.180 ;
        RECT 86.455 116.935 86.795 117.745 ;
        RECT 87.445 117.485 87.775 117.735 ;
        RECT 87.945 117.325 88.195 117.925 ;
        RECT 86.280 116.525 86.795 116.935 ;
        RECT 83.675 116.345 85.705 116.515 ;
        RECT 87.865 116.345 88.195 117.325 ;
        RECT 89.640 118.015 89.895 118.215 ;
        RECT 89.640 117.155 89.820 118.015 ;
        RECT 90.540 117.815 90.790 118.465 ;
        RECT 89.990 117.485 90.790 117.815 ;
        RECT 89.640 116.485 89.895 117.155 ;
        RECT 90.540 116.895 90.790 117.485 ;
        RECT 90.990 118.130 91.310 118.460 ;
        RECT 92.350 118.335 93.200 118.505 ;
        RECT 90.990 117.235 91.180 118.130 ;
        RECT 91.500 117.805 92.160 118.075 ;
        RECT 91.830 117.745 92.160 117.805 ;
        RECT 91.350 117.575 91.680 117.635 ;
        RECT 92.350 117.575 92.520 118.335 ;
        RECT 94.280 118.085 94.530 118.515 ;
        RECT 92.690 117.915 93.940 118.085 ;
        RECT 92.690 117.795 93.020 117.915 ;
        RECT 91.350 117.405 93.250 117.575 ;
        RECT 90.990 117.065 92.910 117.235 ;
        RECT 90.990 117.045 91.310 117.065 ;
        RECT 90.540 116.385 90.870 116.895 ;
        RECT 91.140 116.435 91.310 117.045 ;
        RECT 93.080 116.895 93.250 117.405 ;
        RECT 93.420 117.335 93.600 117.745 ;
        RECT 93.770 117.155 93.940 117.915 ;
        RECT 92.040 116.725 93.250 116.895 ;
        RECT 93.420 116.845 93.940 117.155 ;
        RECT 94.110 117.745 94.530 118.085 ;
        RECT 95.400 118.345 96.415 118.545 ;
        RECT 94.820 117.745 95.230 118.075 ;
        RECT 94.110 116.975 94.300 117.745 ;
        RECT 95.400 117.615 95.570 118.345 ;
        RECT 96.715 118.175 96.885 118.505 ;
        RECT 95.740 117.795 96.090 118.165 ;
        RECT 95.400 117.575 95.820 117.615 ;
        RECT 94.470 117.405 95.820 117.575 ;
        RECT 94.470 117.245 94.720 117.405 ;
        RECT 95.230 116.975 95.480 117.235 ;
        RECT 94.110 116.725 95.480 116.975 ;
        RECT 92.040 116.435 92.280 116.725 ;
        RECT 93.080 116.645 93.250 116.725 ;
        RECT 93.080 116.395 93.710 116.645 ;
        RECT 94.680 116.435 94.850 116.725 ;
        RECT 95.650 116.560 95.820 117.405 ;
        RECT 96.270 117.235 96.490 118.105 ;
        RECT 96.715 117.985 97.410 118.175 ;
        RECT 95.990 116.855 96.490 117.235 ;
        RECT 96.660 117.185 97.070 117.805 ;
        RECT 97.240 117.015 97.410 117.985 ;
        RECT 96.715 116.845 97.410 117.015 ;
        RECT 95.650 116.390 96.480 116.560 ;
        RECT 96.715 116.345 96.885 116.845 ;
        RECT 97.600 116.345 97.825 118.465 ;
        RECT 98.495 118.175 98.665 118.465 ;
        RECT 98.000 118.005 98.665 118.175 ;
        RECT 98.925 118.050 99.185 118.555 ;
        RECT 99.875 118.175 100.045 118.555 ;
        RECT 101.600 118.385 101.855 118.545 ;
        RECT 101.515 118.215 101.855 118.385 ;
        RECT 98.000 117.015 98.230 118.005 ;
        RECT 98.400 117.185 98.750 117.835 ;
        RECT 98.925 117.250 99.095 118.050 ;
        RECT 99.380 118.005 100.045 118.175 ;
        RECT 101.600 118.015 101.855 118.215 ;
        RECT 99.380 117.750 99.550 118.005 ;
        RECT 99.265 117.420 99.550 117.750 ;
        RECT 99.785 117.455 100.115 117.825 ;
        RECT 99.380 117.275 99.550 117.420 ;
        RECT 98.000 116.845 98.665 117.015 ;
        RECT 98.495 116.345 98.665 116.845 ;
        RECT 98.925 116.345 99.195 117.250 ;
        RECT 99.380 117.105 100.045 117.275 ;
        RECT 99.875 116.345 100.045 117.105 ;
        RECT 101.600 117.155 101.780 118.015 ;
        RECT 102.500 117.815 102.750 118.465 ;
        RECT 101.950 117.485 102.750 117.815 ;
        RECT 101.600 116.485 101.855 117.155 ;
        RECT 102.500 116.895 102.750 117.485 ;
        RECT 102.950 118.130 103.270 118.460 ;
        RECT 104.310 118.335 105.160 118.505 ;
        RECT 102.950 117.235 103.140 118.130 ;
        RECT 103.460 117.805 104.120 118.075 ;
        RECT 103.790 117.745 104.120 117.805 ;
        RECT 103.310 117.575 103.640 117.635 ;
        RECT 104.310 117.575 104.480 118.335 ;
        RECT 106.240 118.085 106.490 118.515 ;
        RECT 104.650 117.915 105.900 118.085 ;
        RECT 104.650 117.795 104.980 117.915 ;
        RECT 103.310 117.405 105.210 117.575 ;
        RECT 102.950 117.065 104.870 117.235 ;
        RECT 102.950 117.045 103.270 117.065 ;
        RECT 102.500 116.385 102.830 116.895 ;
        RECT 103.100 116.435 103.270 117.045 ;
        RECT 105.040 116.895 105.210 117.405 ;
        RECT 105.380 117.335 105.560 117.745 ;
        RECT 105.730 117.155 105.900 117.915 ;
        RECT 104.000 116.725 105.210 116.895 ;
        RECT 105.380 116.845 105.900 117.155 ;
        RECT 106.070 117.745 106.490 118.085 ;
        RECT 107.360 118.345 108.375 118.545 ;
        RECT 106.780 117.745 107.190 118.075 ;
        RECT 106.070 116.975 106.260 117.745 ;
        RECT 107.360 117.615 107.530 118.345 ;
        RECT 108.675 118.175 108.845 118.505 ;
        RECT 107.700 117.795 108.050 118.165 ;
        RECT 107.360 117.575 107.780 117.615 ;
        RECT 106.430 117.405 107.780 117.575 ;
        RECT 106.430 117.245 106.680 117.405 ;
        RECT 107.190 116.975 107.440 117.235 ;
        RECT 106.070 116.725 107.440 116.975 ;
        RECT 104.000 116.435 104.240 116.725 ;
        RECT 105.040 116.645 105.210 116.725 ;
        RECT 105.040 116.395 105.670 116.645 ;
        RECT 106.640 116.435 106.810 116.725 ;
        RECT 107.610 116.560 107.780 117.405 ;
        RECT 108.230 117.235 108.450 118.105 ;
        RECT 108.675 117.985 109.370 118.175 ;
        RECT 107.950 116.855 108.450 117.235 ;
        RECT 108.620 117.185 109.030 117.805 ;
        RECT 109.200 117.015 109.370 117.985 ;
        RECT 108.675 116.845 109.370 117.015 ;
        RECT 107.610 116.390 108.440 116.560 ;
        RECT 108.675 116.345 108.845 116.845 ;
        RECT 109.560 116.345 109.785 118.465 ;
        RECT 110.455 118.175 110.625 118.465 ;
        RECT 109.960 118.005 110.625 118.175 ;
        RECT 110.885 118.050 111.145 118.555 ;
        RECT 111.835 118.175 112.005 118.555 ;
        RECT 109.960 117.015 110.190 118.005 ;
        RECT 110.360 117.185 110.710 117.835 ;
        RECT 110.885 117.250 111.055 118.050 ;
        RECT 111.340 118.005 112.005 118.175 ;
        RECT 111.340 117.750 111.510 118.005 ;
        RECT 113.165 117.925 113.495 118.555 ;
        RECT 115.575 118.175 115.745 118.555 ;
        RECT 115.575 118.005 116.240 118.175 ;
        RECT 116.435 118.050 116.695 118.555 ;
        RECT 111.225 117.420 111.510 117.750 ;
        RECT 111.745 117.455 112.075 117.825 ;
        RECT 111.340 117.275 111.510 117.420 ;
        RECT 113.165 117.325 113.415 117.925 ;
        RECT 113.585 117.485 113.915 117.735 ;
        RECT 115.505 117.455 115.835 117.825 ;
        RECT 116.070 117.750 116.240 118.005 ;
        RECT 116.070 117.420 116.355 117.750 ;
        RECT 109.960 116.845 110.625 117.015 ;
        RECT 110.455 116.345 110.625 116.845 ;
        RECT 110.885 116.345 111.155 117.250 ;
        RECT 111.340 117.105 112.005 117.275 ;
        RECT 111.835 116.345 112.005 117.105 ;
        RECT 113.165 116.345 113.495 117.325 ;
        RECT 116.070 117.275 116.240 117.420 ;
        RECT 115.575 117.105 116.240 117.275 ;
        RECT 116.525 117.250 116.695 118.050 ;
        RECT 117.325 117.485 117.640 118.045 ;
        RECT 117.810 117.735 118.060 118.545 ;
        RECT 118.670 117.735 118.920 118.545 ;
        RECT 119.520 118.075 119.780 118.530 ;
        RECT 120.380 118.075 120.640 118.530 ;
        RECT 121.240 118.075 121.500 118.530 ;
        RECT 122.085 118.075 122.360 118.530 ;
        RECT 122.945 118.075 123.205 118.530 ;
        RECT 123.805 118.075 124.065 118.530 ;
        RECT 124.665 118.075 124.925 118.530 ;
        RECT 125.535 118.075 125.795 118.530 ;
        RECT 119.520 117.905 126.265 118.075 ;
        RECT 117.810 117.485 124.930 117.735 ;
        RECT 115.575 116.345 115.745 117.105 ;
        RECT 116.425 116.345 116.695 117.250 ;
        RECT 117.810 116.345 118.055 117.485 ;
        RECT 118.670 116.350 118.920 117.485 ;
        RECT 125.100 117.365 126.265 117.905 ;
        RECT 125.100 117.315 126.295 117.365 ;
        RECT 119.520 117.195 126.295 117.315 ;
        RECT 119.520 117.090 126.265 117.195 ;
        RECT 119.520 117.075 124.925 117.090 ;
        RECT 119.520 116.350 119.780 117.075 ;
        RECT 120.380 116.350 120.640 117.075 ;
        RECT 121.240 116.350 121.500 117.075 ;
        RECT 122.100 116.350 122.360 117.075 ;
        RECT 122.945 116.350 123.205 117.075 ;
        RECT 123.805 116.350 124.065 117.075 ;
        RECT 124.665 116.350 124.925 117.075 ;
        RECT 125.535 116.350 125.825 117.090 ;
        RECT 20.705 114.855 21.035 115.835 ;
        RECT 20.285 114.445 20.615 114.695 ;
        RECT 20.785 114.255 21.035 114.855 ;
        RECT 20.705 113.625 21.035 114.255 ;
        RECT 22.085 114.855 22.415 115.835 ;
        RECT 23.115 115.075 23.285 115.835 ;
        RECT 23.115 114.905 23.780 115.075 ;
        RECT 23.965 114.930 24.235 115.835 ;
        RECT 22.085 114.255 22.335 114.855 ;
        RECT 23.610 114.760 23.780 114.905 ;
        RECT 22.505 114.445 22.835 114.695 ;
        RECT 23.045 114.355 23.375 114.725 ;
        RECT 23.610 114.430 23.895 114.760 ;
        RECT 22.085 113.625 22.415 114.255 ;
        RECT 23.610 114.175 23.780 114.430 ;
        RECT 23.115 114.005 23.780 114.175 ;
        RECT 24.065 114.130 24.235 114.930 ;
        RECT 25.350 114.695 25.595 115.835 ;
        RECT 26.210 114.695 26.460 115.830 ;
        RECT 27.060 115.105 27.320 115.830 ;
        RECT 27.920 115.105 28.180 115.830 ;
        RECT 28.780 115.105 29.040 115.830 ;
        RECT 29.640 115.105 29.900 115.830 ;
        RECT 30.485 115.105 30.745 115.830 ;
        RECT 31.345 115.105 31.605 115.830 ;
        RECT 32.205 115.105 32.465 115.830 ;
        RECT 27.060 115.090 32.465 115.105 ;
        RECT 33.075 115.090 33.365 115.830 ;
        RECT 34.595 115.090 34.885 115.830 ;
        RECT 35.495 115.105 35.755 115.830 ;
        RECT 36.355 115.105 36.615 115.830 ;
        RECT 37.215 115.105 37.475 115.830 ;
        RECT 38.060 115.105 38.320 115.830 ;
        RECT 38.920 115.105 39.180 115.830 ;
        RECT 39.780 115.105 40.040 115.830 ;
        RECT 40.640 115.105 40.900 115.830 ;
        RECT 35.495 115.090 40.900 115.105 ;
        RECT 27.060 114.865 33.805 115.090 ;
        RECT 34.155 114.985 40.900 115.090 ;
        RECT 24.865 114.135 25.180 114.695 ;
        RECT 25.350 114.445 32.470 114.695 ;
        RECT 23.115 113.625 23.285 114.005 ;
        RECT 23.975 113.625 24.235 114.130 ;
        RECT 25.350 113.635 25.600 114.445 ;
        RECT 26.210 113.635 26.460 114.445 ;
        RECT 32.640 114.275 33.805 114.865 ;
        RECT 34.125 114.865 40.900 114.985 ;
        RECT 34.125 114.815 35.320 114.865 ;
        RECT 27.060 114.105 33.805 114.275 ;
        RECT 34.155 114.275 35.320 114.815 ;
        RECT 41.500 114.695 41.750 115.830 ;
        RECT 42.365 114.695 42.610 115.835 ;
        RECT 43.265 114.930 43.535 115.835 ;
        RECT 44.215 115.075 44.385 115.835 ;
        RECT 35.490 114.445 42.610 114.695 ;
        RECT 34.155 114.105 40.900 114.275 ;
        RECT 27.060 113.650 27.320 114.105 ;
        RECT 27.920 113.650 28.180 114.105 ;
        RECT 28.780 113.650 29.040 114.105 ;
        RECT 29.625 113.650 29.900 114.105 ;
        RECT 30.485 113.650 30.745 114.105 ;
        RECT 31.345 113.650 31.605 114.105 ;
        RECT 32.205 113.650 32.465 114.105 ;
        RECT 33.075 113.650 33.335 114.105 ;
        RECT 34.625 113.650 34.885 114.105 ;
        RECT 35.495 113.650 35.755 114.105 ;
        RECT 36.355 113.650 36.615 114.105 ;
        RECT 37.215 113.650 37.475 114.105 ;
        RECT 38.060 113.650 38.335 114.105 ;
        RECT 38.920 113.650 39.180 114.105 ;
        RECT 39.780 113.650 40.040 114.105 ;
        RECT 40.640 113.650 40.900 114.105 ;
        RECT 41.500 113.635 41.750 114.445 ;
        RECT 42.360 113.635 42.610 114.445 ;
        RECT 42.780 114.135 43.095 114.695 ;
        RECT 43.265 114.130 43.435 114.930 ;
        RECT 43.720 114.905 44.385 115.075 ;
        RECT 43.720 114.760 43.890 114.905 ;
        RECT 43.605 114.430 43.890 114.760 ;
        RECT 45.085 114.855 45.415 115.835 ;
        RECT 47.865 114.930 48.135 115.835 ;
        RECT 48.815 115.075 48.985 115.835 ;
        RECT 43.720 114.175 43.890 114.430 ;
        RECT 44.125 114.355 44.455 114.725 ;
        RECT 45.085 114.255 45.335 114.855 ;
        RECT 45.505 114.445 45.835 114.695 ;
        RECT 43.265 113.625 43.525 114.130 ;
        RECT 43.720 114.005 44.385 114.175 ;
        RECT 44.215 113.625 44.385 114.005 ;
        RECT 45.085 113.625 45.415 114.255 ;
        RECT 47.865 114.130 48.035 114.930 ;
        RECT 48.320 114.905 48.985 115.075 ;
        RECT 52.555 115.075 52.725 115.835 ;
        RECT 52.555 114.905 53.220 115.075 ;
        RECT 53.405 114.930 53.675 115.835 ;
        RECT 48.320 114.760 48.490 114.905 ;
        RECT 48.205 114.430 48.490 114.760 ;
        RECT 53.050 114.760 53.220 114.905 ;
        RECT 48.320 114.175 48.490 114.430 ;
        RECT 48.725 114.355 49.055 114.725 ;
        RECT 52.485 114.355 52.815 114.725 ;
        RECT 53.050 114.430 53.335 114.760 ;
        RECT 53.050 114.175 53.220 114.430 ;
        RECT 47.865 113.625 48.125 114.130 ;
        RECT 48.320 114.005 48.985 114.175 ;
        RECT 48.815 113.625 48.985 114.005 ;
        RECT 52.555 114.005 53.220 114.175 ;
        RECT 53.505 114.130 53.675 114.930 ;
        RECT 66.245 114.855 66.575 115.835 ;
        RECT 68.195 115.075 68.365 115.835 ;
        RECT 68.195 114.905 68.860 115.075 ;
        RECT 69.045 114.930 69.315 115.835 ;
        RECT 77.680 115.665 77.935 115.695 ;
        RECT 77.595 115.495 77.935 115.665 ;
        RECT 65.825 114.445 66.155 114.695 ;
        RECT 66.325 114.255 66.575 114.855 ;
        RECT 68.690 114.760 68.860 114.905 ;
        RECT 68.125 114.355 68.455 114.725 ;
        RECT 68.690 114.430 68.975 114.760 ;
        RECT 52.555 113.625 52.725 114.005 ;
        RECT 53.415 113.625 53.675 114.130 ;
        RECT 66.245 113.625 66.575 114.255 ;
        RECT 68.690 114.175 68.860 114.430 ;
        RECT 68.195 114.005 68.860 114.175 ;
        RECT 69.145 114.130 69.315 114.930 ;
        RECT 68.195 113.625 68.365 114.005 ;
        RECT 69.055 113.625 69.315 114.130 ;
        RECT 77.680 115.025 77.935 115.495 ;
        RECT 78.580 115.285 78.910 115.795 ;
        RECT 77.680 114.165 77.860 115.025 ;
        RECT 78.580 114.695 78.830 115.285 ;
        RECT 79.180 115.135 79.350 115.745 ;
        RECT 80.080 115.455 80.320 115.745 ;
        RECT 81.120 115.535 81.750 115.785 ;
        RECT 81.120 115.455 81.290 115.535 ;
        RECT 82.720 115.455 82.890 115.745 ;
        RECT 83.690 115.620 84.520 115.790 ;
        RECT 80.080 115.285 81.290 115.455 ;
        RECT 78.030 114.365 78.830 114.695 ;
        RECT 77.680 113.635 77.935 114.165 ;
        RECT 78.580 113.715 78.830 114.365 ;
        RECT 79.030 115.115 79.350 115.135 ;
        RECT 79.030 114.945 80.950 115.115 ;
        RECT 79.030 114.050 79.220 114.945 ;
        RECT 81.120 114.775 81.290 115.285 ;
        RECT 81.460 115.025 81.980 115.335 ;
        RECT 79.390 114.605 81.290 114.775 ;
        RECT 79.390 114.545 79.720 114.605 ;
        RECT 79.870 114.375 80.200 114.435 ;
        RECT 79.540 114.105 80.200 114.375 ;
        RECT 79.030 113.720 79.350 114.050 ;
        RECT 80.390 113.845 80.560 114.605 ;
        RECT 81.460 114.435 81.640 114.845 ;
        RECT 80.730 114.265 81.060 114.385 ;
        RECT 81.810 114.265 81.980 115.025 ;
        RECT 80.730 114.095 81.980 114.265 ;
        RECT 82.150 115.205 83.520 115.455 ;
        RECT 82.150 114.435 82.340 115.205 ;
        RECT 83.270 114.945 83.520 115.205 ;
        RECT 82.510 114.775 82.760 114.935 ;
        RECT 83.690 114.775 83.860 115.620 ;
        RECT 84.755 115.335 84.925 115.835 ;
        RECT 84.030 114.945 84.530 115.325 ;
        RECT 84.755 115.165 85.450 115.335 ;
        RECT 82.510 114.605 83.860 114.775 ;
        RECT 83.440 114.565 83.860 114.605 ;
        RECT 82.150 114.095 82.570 114.435 ;
        RECT 82.860 114.105 83.270 114.435 ;
        RECT 80.390 113.675 81.240 113.845 ;
        RECT 82.320 113.665 82.570 114.095 ;
        RECT 83.440 113.835 83.610 114.565 ;
        RECT 83.780 114.015 84.130 114.385 ;
        RECT 84.310 114.075 84.530 114.945 ;
        RECT 84.700 114.375 85.110 114.995 ;
        RECT 85.280 114.195 85.450 115.165 ;
        RECT 84.755 114.005 85.450 114.195 ;
        RECT 83.440 113.635 84.455 113.835 ;
        RECT 84.755 113.675 84.925 114.005 ;
        RECT 85.640 113.715 85.865 115.835 ;
        RECT 86.535 115.335 86.705 115.835 ;
        RECT 92.195 115.665 94.225 115.835 ;
        RECT 86.040 115.165 86.705 115.335 ;
        RECT 91.105 115.245 91.620 115.655 ;
        RECT 86.040 114.175 86.270 115.165 ;
        RECT 86.440 114.345 86.790 114.995 ;
        RECT 91.105 114.435 91.445 115.245 ;
        RECT 92.195 115.000 92.365 115.665 ;
        RECT 92.760 115.325 93.885 115.495 ;
        RECT 91.615 114.810 92.365 115.000 ;
        RECT 92.535 114.985 93.545 115.155 ;
        RECT 91.105 114.265 92.335 114.435 ;
        RECT 86.040 114.005 86.705 114.175 ;
        RECT 86.535 113.715 86.705 114.005 ;
        RECT 91.380 113.660 91.625 114.265 ;
        RECT 92.535 113.625 92.725 114.985 ;
        RECT 92.895 114.645 93.170 114.785 ;
        RECT 92.895 114.475 93.175 114.645 ;
        RECT 92.895 113.625 93.170 114.475 ;
        RECT 93.375 114.185 93.545 114.985 ;
        RECT 93.715 114.195 93.885 115.325 ;
        RECT 94.055 114.695 94.225 115.665 ;
        RECT 94.735 114.865 95.070 115.835 ;
        RECT 98.635 115.665 100.665 115.835 ;
        RECT 94.055 114.365 94.250 114.695 ;
        RECT 94.475 114.365 94.730 114.695 ;
        RECT 94.475 114.195 94.645 114.365 ;
        RECT 94.900 114.195 95.070 114.865 ;
        RECT 97.545 115.245 98.060 115.655 ;
        RECT 97.545 114.435 97.885 115.245 ;
        RECT 98.635 115.000 98.805 115.665 ;
        RECT 99.200 115.325 100.325 115.495 ;
        RECT 98.055 114.810 98.805 115.000 ;
        RECT 98.975 114.985 99.985 115.155 ;
        RECT 97.545 114.265 98.775 114.435 ;
        RECT 93.715 114.025 94.645 114.195 ;
        RECT 93.715 113.990 93.890 114.025 ;
        RECT 93.360 113.625 93.890 113.990 ;
        RECT 94.815 113.625 95.070 114.195 ;
        RECT 97.820 113.660 98.065 114.265 ;
        RECT 98.975 113.625 99.165 114.985 ;
        RECT 99.335 114.645 99.610 114.785 ;
        RECT 99.335 114.475 99.615 114.645 ;
        RECT 99.335 113.625 99.610 114.475 ;
        RECT 99.815 114.185 99.985 114.985 ;
        RECT 100.155 114.195 100.325 115.325 ;
        RECT 100.495 114.695 100.665 115.665 ;
        RECT 101.175 114.865 101.510 115.835 ;
        RECT 112.435 115.665 114.465 115.835 ;
        RECT 100.495 114.365 100.690 114.695 ;
        RECT 100.915 114.365 101.170 114.695 ;
        RECT 100.915 114.195 101.085 114.365 ;
        RECT 101.340 114.195 101.510 114.865 ;
        RECT 111.345 115.245 111.860 115.655 ;
        RECT 111.345 114.435 111.685 115.245 ;
        RECT 112.435 115.000 112.605 115.665 ;
        RECT 113.000 115.325 114.125 115.495 ;
        RECT 111.855 114.810 112.605 115.000 ;
        RECT 112.775 114.985 113.785 115.155 ;
        RECT 111.345 114.265 112.575 114.435 ;
        RECT 100.155 114.025 101.085 114.195 ;
        RECT 100.155 113.990 100.330 114.025 ;
        RECT 99.800 113.625 100.330 113.990 ;
        RECT 101.255 113.625 101.510 114.195 ;
        RECT 111.620 113.660 111.865 114.265 ;
        RECT 112.775 113.625 112.965 114.985 ;
        RECT 113.135 114.645 113.410 114.785 ;
        RECT 113.135 114.475 113.415 114.645 ;
        RECT 113.135 113.625 113.410 114.475 ;
        RECT 113.615 114.185 113.785 114.985 ;
        RECT 113.955 114.195 114.125 115.325 ;
        RECT 114.295 114.695 114.465 115.665 ;
        RECT 114.975 114.865 115.310 115.835 ;
        RECT 117.330 115.335 117.585 115.835 ;
        RECT 117.330 115.165 118.080 115.335 ;
        RECT 114.295 114.365 114.490 114.695 ;
        RECT 114.715 114.365 114.970 114.695 ;
        RECT 114.715 114.195 114.885 114.365 ;
        RECT 115.140 114.195 115.310 114.865 ;
        RECT 117.330 114.345 117.680 114.995 ;
        RECT 113.955 114.025 114.885 114.195 ;
        RECT 113.955 113.990 114.130 114.025 ;
        RECT 113.600 113.625 114.130 113.990 ;
        RECT 115.055 113.625 115.310 114.195 ;
        RECT 117.850 114.175 118.080 115.165 ;
        RECT 117.330 114.005 118.080 114.175 ;
        RECT 117.330 113.715 117.585 114.005 ;
        RECT 118.255 113.715 118.425 115.835 ;
        RECT 118.595 115.035 118.920 115.820 ;
        RECT 119.510 115.505 119.760 115.835 ;
        RECT 119.975 115.505 120.655 115.835 ;
        RECT 119.510 115.375 119.680 115.505 ;
        RECT 119.285 115.205 119.680 115.375 ;
        RECT 118.655 113.985 119.115 115.035 ;
        RECT 119.285 113.845 119.455 115.205 ;
        RECT 119.850 114.945 120.315 115.335 ;
        RECT 119.625 114.135 119.975 114.755 ;
        RECT 120.145 114.355 120.315 114.945 ;
        RECT 120.485 114.725 120.655 115.505 ;
        RECT 120.825 115.405 120.995 115.745 ;
        RECT 121.730 115.405 121.900 115.745 ;
        RECT 120.825 115.235 121.900 115.405 ;
        RECT 122.735 115.375 122.905 115.835 ;
        RECT 123.140 115.495 124.010 115.835 ;
        RECT 122.345 115.205 122.905 115.375 ;
        RECT 122.345 115.065 122.515 115.205 ;
        RECT 121.015 114.895 122.515 115.065 ;
        RECT 123.210 115.035 123.670 115.325 ;
        RECT 120.485 114.555 122.175 114.725 ;
        RECT 120.145 114.135 120.500 114.355 ;
        RECT 120.670 113.845 120.840 114.555 ;
        RECT 121.045 114.135 121.835 114.385 ;
        RECT 122.005 114.375 122.175 114.555 ;
        RECT 122.345 114.205 122.515 114.895 ;
        RECT 119.285 113.675 119.780 113.845 ;
        RECT 119.985 113.675 120.840 113.845 ;
        RECT 122.255 113.815 122.515 114.205 ;
        RECT 122.705 115.025 123.670 115.035 ;
        RECT 123.840 115.115 124.010 115.495 ;
        RECT 124.600 115.455 124.770 115.745 ;
        RECT 124.600 115.285 125.400 115.455 ;
        RECT 122.705 114.865 123.380 115.025 ;
        RECT 123.840 114.945 125.060 115.115 ;
        RECT 122.705 114.075 122.915 114.865 ;
        RECT 123.840 114.855 124.010 114.945 ;
        RECT 123.085 114.075 123.435 114.695 ;
        RECT 123.605 114.685 124.010 114.855 ;
        RECT 123.605 113.905 123.775 114.685 ;
        RECT 123.945 114.235 124.165 114.515 ;
        RECT 124.345 114.405 124.885 114.775 ;
        RECT 125.230 114.695 125.400 115.285 ;
        RECT 126.095 114.815 126.350 115.695 ;
        RECT 125.230 114.665 125.970 114.695 ;
        RECT 123.945 114.065 124.475 114.235 ;
        RECT 122.255 113.645 122.605 113.815 ;
        RECT 122.825 113.625 123.775 113.905 ;
        RECT 124.305 113.835 124.475 114.065 ;
        RECT 124.645 114.005 124.885 114.405 ;
        RECT 125.055 114.365 125.970 114.665 ;
        RECT 125.055 114.190 125.380 114.365 ;
        RECT 125.055 113.835 125.375 114.190 ;
        RECT 126.140 114.165 126.350 114.815 ;
        RECT 124.305 113.665 125.375 113.835 ;
        RECT 126.095 113.635 126.350 114.165 ;
        RECT 17.420 112.945 17.675 113.105 ;
        RECT 17.335 112.775 17.675 112.945 ;
        RECT 17.420 112.575 17.675 112.775 ;
        RECT 17.420 111.715 17.600 112.575 ;
        RECT 18.320 112.375 18.570 113.025 ;
        RECT 17.770 112.045 18.570 112.375 ;
        RECT 17.420 111.045 17.675 111.715 ;
        RECT 18.320 111.455 18.570 112.045 ;
        RECT 18.770 112.690 19.090 113.020 ;
        RECT 20.130 112.895 20.980 113.065 ;
        RECT 18.770 111.795 18.960 112.690 ;
        RECT 19.280 112.365 19.940 112.635 ;
        RECT 19.610 112.305 19.940 112.365 ;
        RECT 19.130 112.135 19.460 112.195 ;
        RECT 20.130 112.135 20.300 112.895 ;
        RECT 22.060 112.645 22.310 113.075 ;
        RECT 20.470 112.475 21.720 112.645 ;
        RECT 20.470 112.355 20.800 112.475 ;
        RECT 19.130 111.965 21.030 112.135 ;
        RECT 18.770 111.625 20.690 111.795 ;
        RECT 18.770 111.605 19.090 111.625 ;
        RECT 18.320 110.945 18.650 111.455 ;
        RECT 18.920 110.995 19.090 111.605 ;
        RECT 20.860 111.455 21.030 111.965 ;
        RECT 21.200 111.895 21.380 112.305 ;
        RECT 21.550 111.715 21.720 112.475 ;
        RECT 19.820 111.285 21.030 111.455 ;
        RECT 21.200 111.405 21.720 111.715 ;
        RECT 21.890 112.305 22.310 112.645 ;
        RECT 23.180 112.905 24.195 113.105 ;
        RECT 22.600 112.305 23.010 112.635 ;
        RECT 21.890 111.535 22.080 112.305 ;
        RECT 23.180 112.175 23.350 112.905 ;
        RECT 24.495 112.735 24.665 113.065 ;
        RECT 23.520 112.355 23.870 112.725 ;
        RECT 23.180 112.135 23.600 112.175 ;
        RECT 22.250 111.965 23.600 112.135 ;
        RECT 22.250 111.805 22.500 111.965 ;
        RECT 23.010 111.535 23.260 111.795 ;
        RECT 21.890 111.285 23.260 111.535 ;
        RECT 19.820 110.995 20.060 111.285 ;
        RECT 20.860 111.205 21.030 111.285 ;
        RECT 20.860 110.955 21.490 111.205 ;
        RECT 22.460 110.995 22.630 111.285 ;
        RECT 23.430 111.120 23.600 111.965 ;
        RECT 24.050 111.795 24.270 112.665 ;
        RECT 24.495 112.545 25.190 112.735 ;
        RECT 23.770 111.415 24.270 111.795 ;
        RECT 24.440 111.745 24.850 112.365 ;
        RECT 25.020 111.575 25.190 112.545 ;
        RECT 24.495 111.405 25.190 111.575 ;
        RECT 23.430 110.950 24.260 111.120 ;
        RECT 24.495 110.905 24.665 111.405 ;
        RECT 25.380 110.905 25.605 113.025 ;
        RECT 26.275 112.735 26.445 113.025 ;
        RECT 25.780 112.565 26.445 112.735 ;
        RECT 26.710 112.735 26.965 113.025 ;
        RECT 26.710 112.565 27.460 112.735 ;
        RECT 25.780 111.575 26.010 112.565 ;
        RECT 26.180 111.745 26.530 112.395 ;
        RECT 26.710 111.745 27.060 112.395 ;
        RECT 27.230 111.575 27.460 112.565 ;
        RECT 25.780 111.405 26.445 111.575 ;
        RECT 26.275 110.905 26.445 111.405 ;
        RECT 26.710 111.405 27.460 111.575 ;
        RECT 26.710 110.905 26.965 111.405 ;
        RECT 27.635 110.905 27.805 113.025 ;
        RECT 28.665 112.895 29.160 113.065 ;
        RECT 29.365 112.895 30.220 113.065 ;
        RECT 28.035 111.705 28.495 112.755 ;
        RECT 27.975 110.920 28.300 111.705 ;
        RECT 28.665 111.535 28.835 112.895 ;
        RECT 29.005 111.985 29.355 112.605 ;
        RECT 29.525 112.385 29.880 112.605 ;
        RECT 29.525 111.795 29.695 112.385 ;
        RECT 30.050 112.185 30.220 112.895 ;
        RECT 31.635 112.925 31.985 113.095 ;
        RECT 30.425 112.355 31.215 112.605 ;
        RECT 31.635 112.535 31.895 112.925 ;
        RECT 32.205 112.835 33.155 113.115 ;
        RECT 31.385 112.185 31.555 112.365 ;
        RECT 28.665 111.365 29.060 111.535 ;
        RECT 29.230 111.405 29.695 111.795 ;
        RECT 29.865 112.015 31.555 112.185 ;
        RECT 28.890 111.235 29.060 111.365 ;
        RECT 29.865 111.235 30.035 112.015 ;
        RECT 31.725 111.845 31.895 112.535 ;
        RECT 30.395 111.675 31.895 111.845 ;
        RECT 32.085 111.875 32.295 112.665 ;
        RECT 32.465 112.045 32.815 112.665 ;
        RECT 32.985 112.055 33.155 112.835 ;
        RECT 33.685 112.905 34.755 113.075 ;
        RECT 33.685 112.675 33.855 112.905 ;
        RECT 33.325 112.505 33.855 112.675 ;
        RECT 33.325 112.225 33.545 112.505 ;
        RECT 34.025 112.335 34.265 112.735 ;
        RECT 32.985 111.885 33.390 112.055 ;
        RECT 33.725 111.965 34.265 112.335 ;
        RECT 34.435 112.550 34.755 112.905 ;
        RECT 35.475 112.575 35.730 113.105 ;
        RECT 34.435 112.375 34.760 112.550 ;
        RECT 34.435 112.075 35.350 112.375 ;
        RECT 34.610 112.045 35.350 112.075 ;
        RECT 32.085 111.715 32.760 111.875 ;
        RECT 33.220 111.795 33.390 111.885 ;
        RECT 32.085 111.705 33.050 111.715 ;
        RECT 31.725 111.535 31.895 111.675 ;
        RECT 28.890 110.905 29.140 111.235 ;
        RECT 29.355 110.905 30.035 111.235 ;
        RECT 30.205 111.335 31.280 111.505 ;
        RECT 31.725 111.365 32.285 111.535 ;
        RECT 32.590 111.415 33.050 111.705 ;
        RECT 33.220 111.625 34.440 111.795 ;
        RECT 30.205 110.995 30.375 111.335 ;
        RECT 31.110 110.995 31.280 111.335 ;
        RECT 32.115 110.905 32.285 111.365 ;
        RECT 33.220 111.245 33.390 111.625 ;
        RECT 34.610 111.455 34.780 112.045 ;
        RECT 35.520 111.925 35.730 112.575 ;
        RECT 32.520 110.905 33.390 111.245 ;
        RECT 33.980 111.285 34.780 111.455 ;
        RECT 33.980 110.995 34.150 111.285 ;
        RECT 35.475 111.045 35.730 111.925 ;
        RECT 35.905 112.610 36.165 113.115 ;
        RECT 36.855 112.735 37.025 113.115 ;
        RECT 35.905 111.810 36.075 112.610 ;
        RECT 36.360 112.565 37.025 112.735 ;
        RECT 36.360 112.310 36.530 112.565 ;
        RECT 36.245 111.980 36.530 112.310 ;
        RECT 36.765 112.015 37.095 112.385 ;
        RECT 37.745 112.045 38.060 112.605 ;
        RECT 38.230 112.295 38.480 113.105 ;
        RECT 39.090 112.295 39.340 113.105 ;
        RECT 39.940 112.635 40.200 113.090 ;
        RECT 40.800 112.635 41.060 113.090 ;
        RECT 41.660 112.635 41.920 113.090 ;
        RECT 42.505 112.635 42.780 113.090 ;
        RECT 43.365 112.635 43.625 113.090 ;
        RECT 44.225 112.635 44.485 113.090 ;
        RECT 45.085 112.635 45.345 113.090 ;
        RECT 45.955 112.635 46.215 113.090 ;
        RECT 39.940 112.465 46.685 112.635 ;
        RECT 79.585 112.485 79.915 113.115 ;
        RECT 38.230 112.045 45.350 112.295 ;
        RECT 36.360 111.835 36.530 111.980 ;
        RECT 35.905 110.905 36.175 111.810 ;
        RECT 36.360 111.665 37.025 111.835 ;
        RECT 36.855 110.905 37.025 111.665 ;
        RECT 38.230 110.905 38.475 112.045 ;
        RECT 39.090 110.910 39.340 112.045 ;
        RECT 45.520 111.875 46.685 112.465 ;
        RECT 79.165 112.045 79.495 112.295 ;
        RECT 79.665 111.885 79.915 112.485 ;
        RECT 39.940 111.650 46.685 111.875 ;
        RECT 39.940 111.635 45.345 111.650 ;
        RECT 39.940 110.910 40.200 111.635 ;
        RECT 40.800 110.910 41.060 111.635 ;
        RECT 41.660 110.910 41.920 111.635 ;
        RECT 42.520 110.910 42.780 111.635 ;
        RECT 43.365 110.910 43.625 111.635 ;
        RECT 44.225 110.910 44.485 111.635 ;
        RECT 45.085 110.910 45.345 111.635 ;
        RECT 45.955 110.910 46.245 111.650 ;
        RECT 79.585 110.905 79.915 111.885 ;
        RECT 81.175 112.635 81.345 113.115 ;
        RECT 82.015 112.635 82.185 113.115 ;
        RECT 82.855 112.635 83.025 113.115 ;
        RECT 81.175 112.465 82.185 112.635 ;
        RECT 82.390 112.465 83.025 112.635 ;
        RECT 93.845 112.485 94.175 113.115 ;
        RECT 106.285 112.610 106.545 113.115 ;
        RECT 107.235 112.735 107.405 113.115 ;
        RECT 81.175 111.925 81.670 112.465 ;
        RECT 82.390 112.295 82.560 112.465 ;
        RECT 82.060 112.125 82.560 112.295 ;
        RECT 81.175 111.755 82.185 111.925 ;
        RECT 81.175 110.905 81.345 111.755 ;
        RECT 82.015 110.905 82.185 111.755 ;
        RECT 82.390 111.885 82.560 112.125 ;
        RECT 82.730 112.055 83.110 112.295 ;
        RECT 93.845 111.885 94.095 112.485 ;
        RECT 94.265 112.045 94.595 112.295 ;
        RECT 82.390 111.715 83.105 111.885 ;
        RECT 82.775 110.905 83.105 111.715 ;
        RECT 93.845 110.905 94.175 111.885 ;
        RECT 106.285 111.810 106.455 112.610 ;
        RECT 106.740 112.565 107.405 112.735 ;
        RECT 115.585 112.635 115.845 113.090 ;
        RECT 116.455 112.635 116.715 113.090 ;
        RECT 117.315 112.635 117.575 113.090 ;
        RECT 118.175 112.635 118.435 113.090 ;
        RECT 119.020 112.635 119.295 113.090 ;
        RECT 119.880 112.635 120.140 113.090 ;
        RECT 120.740 112.635 121.000 113.090 ;
        RECT 121.600 112.635 121.860 113.090 ;
        RECT 106.740 112.310 106.910 112.565 ;
        RECT 115.115 112.465 121.860 112.635 ;
        RECT 106.625 111.980 106.910 112.310 ;
        RECT 107.145 112.015 107.475 112.385 ;
        RECT 106.740 111.835 106.910 111.980 ;
        RECT 115.115 111.875 116.280 112.465 ;
        RECT 122.460 112.295 122.710 113.105 ;
        RECT 123.320 112.295 123.570 113.105 ;
        RECT 124.315 112.735 124.485 113.115 ;
        RECT 116.450 112.045 123.570 112.295 ;
        RECT 123.740 112.045 124.055 112.605 ;
        RECT 124.315 112.565 124.980 112.735 ;
        RECT 125.175 112.610 125.435 113.115 ;
        RECT 106.285 110.905 106.555 111.810 ;
        RECT 106.740 111.665 107.405 111.835 ;
        RECT 107.235 110.905 107.405 111.665 ;
        RECT 115.115 111.650 121.860 111.875 ;
        RECT 115.555 110.910 115.845 111.650 ;
        RECT 116.455 111.635 121.860 111.650 ;
        RECT 116.455 110.910 116.715 111.635 ;
        RECT 117.315 110.910 117.575 111.635 ;
        RECT 118.175 110.910 118.435 111.635 ;
        RECT 119.020 110.910 119.280 111.635 ;
        RECT 119.880 110.910 120.140 111.635 ;
        RECT 120.740 110.910 121.000 111.635 ;
        RECT 121.600 110.910 121.860 111.635 ;
        RECT 122.460 110.910 122.710 112.045 ;
        RECT 123.325 110.905 123.570 112.045 ;
        RECT 124.245 112.015 124.575 112.385 ;
        RECT 124.810 112.310 124.980 112.565 ;
        RECT 124.810 111.980 125.095 112.310 ;
        RECT 124.810 111.835 124.980 111.980 ;
        RECT 124.315 111.665 124.980 111.835 ;
        RECT 125.265 111.810 125.435 112.610 ;
        RECT 124.315 110.905 124.485 111.665 ;
        RECT 125.165 110.905 125.435 111.810 ;
        RECT 23.465 109.415 23.795 110.395 ;
        RECT 26.335 109.635 26.505 110.395 ;
        RECT 26.335 109.465 27.000 109.635 ;
        RECT 27.185 109.490 27.455 110.395 ;
        RECT 23.045 109.005 23.375 109.255 ;
        RECT 23.545 108.815 23.795 109.415 ;
        RECT 26.830 109.320 27.000 109.465 ;
        RECT 26.265 108.915 26.595 109.285 ;
        RECT 26.830 108.990 27.115 109.320 ;
        RECT 23.465 108.185 23.795 108.815 ;
        RECT 26.830 108.735 27.000 108.990 ;
        RECT 26.335 108.565 27.000 108.735 ;
        RECT 27.285 108.690 27.455 109.490 ;
        RECT 27.715 109.635 27.885 110.395 ;
        RECT 27.715 109.465 28.380 109.635 ;
        RECT 28.565 109.490 28.835 110.395 ;
        RECT 28.210 109.320 28.380 109.465 ;
        RECT 27.645 108.915 27.975 109.285 ;
        RECT 28.210 108.990 28.495 109.320 ;
        RECT 28.210 108.735 28.380 108.990 ;
        RECT 26.335 108.185 26.505 108.565 ;
        RECT 27.195 108.185 27.455 108.690 ;
        RECT 27.715 108.565 28.380 108.735 ;
        RECT 28.665 108.690 28.835 109.490 ;
        RECT 29.490 109.255 29.735 110.395 ;
        RECT 30.350 109.255 30.600 110.390 ;
        RECT 31.200 109.665 31.460 110.390 ;
        RECT 32.060 109.665 32.320 110.390 ;
        RECT 32.920 109.665 33.180 110.390 ;
        RECT 33.780 109.665 34.040 110.390 ;
        RECT 34.625 109.665 34.885 110.390 ;
        RECT 35.485 109.665 35.745 110.390 ;
        RECT 36.345 109.665 36.605 110.390 ;
        RECT 31.200 109.650 36.605 109.665 ;
        RECT 37.215 109.650 37.505 110.390 ;
        RECT 38.210 109.895 38.465 110.395 ;
        RECT 38.210 109.725 38.960 109.895 ;
        RECT 31.200 109.425 37.945 109.650 ;
        RECT 29.005 108.695 29.320 109.255 ;
        RECT 29.490 109.005 36.610 109.255 ;
        RECT 27.715 108.185 27.885 108.565 ;
        RECT 28.575 108.185 28.835 108.690 ;
        RECT 29.490 108.195 29.740 109.005 ;
        RECT 30.350 108.195 30.600 109.005 ;
        RECT 36.780 108.835 37.945 109.425 ;
        RECT 38.210 108.905 38.560 109.555 ;
        RECT 31.200 108.665 37.945 108.835 ;
        RECT 38.730 108.735 38.960 109.725 ;
        RECT 31.200 108.210 31.460 108.665 ;
        RECT 32.060 108.210 32.320 108.665 ;
        RECT 32.920 108.210 33.180 108.665 ;
        RECT 33.765 108.210 34.040 108.665 ;
        RECT 34.625 108.210 34.885 108.665 ;
        RECT 35.485 108.210 35.745 108.665 ;
        RECT 36.345 108.210 36.605 108.665 ;
        RECT 37.215 108.210 37.475 108.665 ;
        RECT 38.210 108.565 38.960 108.735 ;
        RECT 38.210 108.275 38.465 108.565 ;
        RECT 39.135 108.275 39.305 110.395 ;
        RECT 39.475 109.595 39.800 110.380 ;
        RECT 40.390 110.065 40.640 110.395 ;
        RECT 40.855 110.065 41.535 110.395 ;
        RECT 40.390 109.935 40.560 110.065 ;
        RECT 40.165 109.765 40.560 109.935 ;
        RECT 39.535 108.545 39.995 109.595 ;
        RECT 40.165 108.405 40.335 109.765 ;
        RECT 40.730 109.505 41.195 109.895 ;
        RECT 40.505 108.695 40.855 109.315 ;
        RECT 41.025 108.915 41.195 109.505 ;
        RECT 41.365 109.285 41.535 110.065 ;
        RECT 41.705 109.965 41.875 110.305 ;
        RECT 42.610 109.965 42.780 110.305 ;
        RECT 41.705 109.795 42.780 109.965 ;
        RECT 43.615 109.935 43.785 110.395 ;
        RECT 44.020 110.055 44.890 110.395 ;
        RECT 43.225 109.765 43.785 109.935 ;
        RECT 43.225 109.625 43.395 109.765 ;
        RECT 41.895 109.455 43.395 109.625 ;
        RECT 44.090 109.595 44.550 109.885 ;
        RECT 41.365 109.115 43.055 109.285 ;
        RECT 41.025 108.695 41.380 108.915 ;
        RECT 41.550 108.405 41.720 109.115 ;
        RECT 41.925 108.695 42.715 108.945 ;
        RECT 42.885 108.935 43.055 109.115 ;
        RECT 43.225 108.765 43.395 109.455 ;
        RECT 40.165 108.235 40.660 108.405 ;
        RECT 40.865 108.235 41.720 108.405 ;
        RECT 43.135 108.375 43.395 108.765 ;
        RECT 43.585 109.585 44.550 109.595 ;
        RECT 44.720 109.675 44.890 110.055 ;
        RECT 45.480 110.015 45.650 110.305 ;
        RECT 45.480 109.845 46.280 110.015 ;
        RECT 43.585 109.425 44.260 109.585 ;
        RECT 44.720 109.505 45.940 109.675 ;
        RECT 43.585 108.635 43.795 109.425 ;
        RECT 44.720 109.415 44.890 109.505 ;
        RECT 43.965 108.635 44.315 109.255 ;
        RECT 44.485 109.245 44.890 109.415 ;
        RECT 44.485 108.465 44.655 109.245 ;
        RECT 44.825 108.795 45.045 109.075 ;
        RECT 45.225 108.965 45.765 109.335 ;
        RECT 46.110 109.255 46.280 109.845 ;
        RECT 46.975 109.375 47.230 110.255 ;
        RECT 47.495 109.635 47.665 110.395 ;
        RECT 47.495 109.465 48.160 109.635 ;
        RECT 48.345 109.490 48.615 110.395 ;
        RECT 46.110 109.225 46.850 109.255 ;
        RECT 44.825 108.625 45.355 108.795 ;
        RECT 43.135 108.205 43.485 108.375 ;
        RECT 43.705 108.185 44.655 108.465 ;
        RECT 45.185 108.395 45.355 108.625 ;
        RECT 45.525 108.565 45.765 108.965 ;
        RECT 45.935 108.925 46.850 109.225 ;
        RECT 45.935 108.750 46.260 108.925 ;
        RECT 45.935 108.395 46.255 108.750 ;
        RECT 47.020 108.725 47.230 109.375 ;
        RECT 47.990 109.320 48.160 109.465 ;
        RECT 47.425 108.915 47.755 109.285 ;
        RECT 47.990 108.990 48.275 109.320 ;
        RECT 47.990 108.735 48.160 108.990 ;
        RECT 45.185 108.225 46.255 108.395 ;
        RECT 46.975 108.195 47.230 108.725 ;
        RECT 47.495 108.565 48.160 108.735 ;
        RECT 48.445 108.690 48.615 109.490 ;
        RECT 51.175 109.635 51.345 110.395 ;
        RECT 51.175 109.465 51.840 109.635 ;
        RECT 52.025 109.490 52.295 110.395 ;
        RECT 51.670 109.320 51.840 109.465 ;
        RECT 51.105 108.915 51.435 109.285 ;
        RECT 51.670 108.990 51.955 109.320 ;
        RECT 51.670 108.735 51.840 108.990 ;
        RECT 47.495 108.185 47.665 108.565 ;
        RECT 48.355 108.185 48.615 108.690 ;
        RECT 51.175 108.565 51.840 108.735 ;
        RECT 52.125 108.690 52.295 109.490 ;
        RECT 57.155 109.635 57.325 110.395 ;
        RECT 57.155 109.465 57.820 109.635 ;
        RECT 58.005 109.490 58.275 110.395 ;
        RECT 57.650 109.320 57.820 109.465 ;
        RECT 57.085 108.915 57.415 109.285 ;
        RECT 57.650 108.990 57.935 109.320 ;
        RECT 57.650 108.735 57.820 108.990 ;
        RECT 51.175 108.185 51.345 108.565 ;
        RECT 52.035 108.185 52.295 108.690 ;
        RECT 57.155 108.565 57.820 108.735 ;
        RECT 58.105 108.690 58.275 109.490 ;
        RECT 60.295 109.585 60.625 110.395 ;
        RECT 60.295 109.415 61.010 109.585 ;
        RECT 60.290 109.005 60.670 109.245 ;
        RECT 60.840 109.175 61.010 109.415 ;
        RECT 61.215 109.545 61.385 110.395 ;
        RECT 62.055 109.545 62.225 110.395 ;
        RECT 61.215 109.375 62.225 109.545 ;
        RECT 63.595 109.635 63.765 110.395 ;
        RECT 63.595 109.465 64.260 109.635 ;
        RECT 64.445 109.490 64.715 110.395 ;
        RECT 65.415 109.650 65.705 110.390 ;
        RECT 66.315 109.665 66.575 110.390 ;
        RECT 67.175 109.665 67.435 110.390 ;
        RECT 68.035 109.665 68.295 110.390 ;
        RECT 68.880 109.665 69.140 110.390 ;
        RECT 69.740 109.665 70.000 110.390 ;
        RECT 70.600 109.665 70.860 110.390 ;
        RECT 71.460 109.665 71.720 110.390 ;
        RECT 66.315 109.650 71.720 109.665 ;
        RECT 60.840 109.005 61.340 109.175 ;
        RECT 60.840 108.835 61.010 109.005 ;
        RECT 61.730 108.865 62.225 109.375 ;
        RECT 64.090 109.320 64.260 109.465 ;
        RECT 63.525 108.915 63.855 109.285 ;
        RECT 64.090 108.990 64.375 109.320 ;
        RECT 61.725 108.835 62.225 108.865 ;
        RECT 57.155 108.185 57.325 108.565 ;
        RECT 58.015 108.185 58.275 108.690 ;
        RECT 60.375 108.665 61.010 108.835 ;
        RECT 61.215 108.665 62.225 108.835 ;
        RECT 64.090 108.735 64.260 108.990 ;
        RECT 60.375 108.185 60.545 108.665 ;
        RECT 61.215 108.185 61.385 108.665 ;
        RECT 62.055 108.185 62.225 108.665 ;
        RECT 63.595 108.565 64.260 108.735 ;
        RECT 64.545 108.690 64.715 109.490 ;
        RECT 63.595 108.185 63.765 108.565 ;
        RECT 64.455 108.185 64.715 108.690 ;
        RECT 64.975 109.425 71.720 109.650 ;
        RECT 64.975 108.835 66.140 109.425 ;
        RECT 72.320 109.255 72.570 110.390 ;
        RECT 73.185 109.255 73.430 110.395 ;
        RECT 74.985 109.415 75.315 110.395 ;
        RECT 77.375 109.650 77.665 110.390 ;
        RECT 78.275 109.665 78.535 110.390 ;
        RECT 79.135 109.665 79.395 110.390 ;
        RECT 79.995 109.665 80.255 110.390 ;
        RECT 80.840 109.665 81.100 110.390 ;
        RECT 81.700 109.665 81.960 110.390 ;
        RECT 82.560 109.665 82.820 110.390 ;
        RECT 83.420 109.665 83.680 110.390 ;
        RECT 78.275 109.650 83.680 109.665 ;
        RECT 76.935 109.425 83.680 109.650 ;
        RECT 66.310 109.005 73.430 109.255 ;
        RECT 64.975 108.665 71.720 108.835 ;
        RECT 65.445 108.210 65.705 108.665 ;
        RECT 66.315 108.210 66.575 108.665 ;
        RECT 67.175 108.210 67.435 108.665 ;
        RECT 68.035 108.210 68.295 108.665 ;
        RECT 68.880 108.210 69.155 108.665 ;
        RECT 69.740 108.210 70.000 108.665 ;
        RECT 70.600 108.210 70.860 108.665 ;
        RECT 71.460 108.210 71.720 108.665 ;
        RECT 72.320 108.195 72.570 109.005 ;
        RECT 73.180 108.195 73.430 109.005 ;
        RECT 73.600 108.695 73.915 109.255 ;
        RECT 74.985 108.815 75.235 109.415 ;
        RECT 75.405 109.005 75.735 109.255 ;
        RECT 76.935 108.835 78.100 109.425 ;
        RECT 84.280 109.255 84.530 110.390 ;
        RECT 85.145 109.255 85.390 110.395 ;
        RECT 86.485 109.415 86.815 110.395 ;
        RECT 87.515 109.635 87.685 110.395 ;
        RECT 87.515 109.465 88.180 109.635 ;
        RECT 88.365 109.490 88.635 110.395 ;
        RECT 89.335 109.650 89.625 110.390 ;
        RECT 90.235 109.665 90.495 110.390 ;
        RECT 91.095 109.665 91.355 110.390 ;
        RECT 91.955 109.665 92.215 110.390 ;
        RECT 92.800 109.665 93.060 110.390 ;
        RECT 93.660 109.665 93.920 110.390 ;
        RECT 94.520 109.665 94.780 110.390 ;
        RECT 95.380 109.665 95.640 110.390 ;
        RECT 90.235 109.650 95.640 109.665 ;
        RECT 78.270 109.005 85.390 109.255 ;
        RECT 74.985 108.185 75.315 108.815 ;
        RECT 76.935 108.665 83.680 108.835 ;
        RECT 77.405 108.210 77.665 108.665 ;
        RECT 78.275 108.210 78.535 108.665 ;
        RECT 79.135 108.210 79.395 108.665 ;
        RECT 79.995 108.210 80.255 108.665 ;
        RECT 80.840 108.210 81.115 108.665 ;
        RECT 81.700 108.210 81.960 108.665 ;
        RECT 82.560 108.210 82.820 108.665 ;
        RECT 83.420 108.210 83.680 108.665 ;
        RECT 84.280 108.195 84.530 109.005 ;
        RECT 85.140 108.195 85.390 109.005 ;
        RECT 85.560 108.695 85.875 109.255 ;
        RECT 86.065 109.005 86.395 109.255 ;
        RECT 86.565 108.815 86.815 109.415 ;
        RECT 88.010 109.320 88.180 109.465 ;
        RECT 87.445 108.915 87.775 109.285 ;
        RECT 88.010 108.990 88.295 109.320 ;
        RECT 86.485 108.185 86.815 108.815 ;
        RECT 88.010 108.735 88.180 108.990 ;
        RECT 87.515 108.565 88.180 108.735 ;
        RECT 88.465 108.690 88.635 109.490 ;
        RECT 87.515 108.185 87.685 108.565 ;
        RECT 88.375 108.185 88.635 108.690 ;
        RECT 88.895 109.425 95.640 109.650 ;
        RECT 88.895 108.835 90.060 109.425 ;
        RECT 96.240 109.255 96.490 110.390 ;
        RECT 97.105 109.255 97.350 110.395 ;
        RECT 99.365 109.415 99.695 110.395 ;
        RECT 100.395 109.635 100.565 110.395 ;
        RECT 100.395 109.465 101.060 109.635 ;
        RECT 101.245 109.490 101.515 110.395 ;
        RECT 102.675 109.650 102.965 110.390 ;
        RECT 103.575 109.665 103.835 110.390 ;
        RECT 104.435 109.665 104.695 110.390 ;
        RECT 105.295 109.665 105.555 110.390 ;
        RECT 106.140 109.665 106.400 110.390 ;
        RECT 107.000 109.665 107.260 110.390 ;
        RECT 107.860 109.665 108.120 110.390 ;
        RECT 108.720 109.665 108.980 110.390 ;
        RECT 103.575 109.650 108.980 109.665 ;
        RECT 90.230 109.005 97.350 109.255 ;
        RECT 88.895 108.665 95.640 108.835 ;
        RECT 89.365 108.210 89.625 108.665 ;
        RECT 90.235 108.210 90.495 108.665 ;
        RECT 91.095 108.210 91.355 108.665 ;
        RECT 91.955 108.210 92.215 108.665 ;
        RECT 92.800 108.210 93.075 108.665 ;
        RECT 93.660 108.210 93.920 108.665 ;
        RECT 94.520 108.210 94.780 108.665 ;
        RECT 95.380 108.210 95.640 108.665 ;
        RECT 96.240 108.195 96.490 109.005 ;
        RECT 97.100 108.195 97.350 109.005 ;
        RECT 97.520 108.695 97.835 109.255 ;
        RECT 98.945 109.005 99.275 109.255 ;
        RECT 99.445 108.815 99.695 109.415 ;
        RECT 100.890 109.320 101.060 109.465 ;
        RECT 100.325 108.915 100.655 109.285 ;
        RECT 100.890 108.990 101.175 109.320 ;
        RECT 99.365 108.185 99.695 108.815 ;
        RECT 100.890 108.735 101.060 108.990 ;
        RECT 100.395 108.565 101.060 108.735 ;
        RECT 101.345 108.690 101.515 109.490 ;
        RECT 100.395 108.185 100.565 108.565 ;
        RECT 101.255 108.185 101.515 108.690 ;
        RECT 102.235 109.425 108.980 109.650 ;
        RECT 102.235 108.835 103.400 109.425 ;
        RECT 109.580 109.255 109.830 110.390 ;
        RECT 110.445 109.255 110.690 110.395 ;
        RECT 111.435 109.635 111.605 110.395 ;
        RECT 111.435 109.465 112.100 109.635 ;
        RECT 112.285 109.490 112.555 110.395 ;
        RECT 111.930 109.320 112.100 109.465 ;
        RECT 103.570 109.005 110.690 109.255 ;
        RECT 102.235 108.665 108.980 108.835 ;
        RECT 102.705 108.210 102.965 108.665 ;
        RECT 103.575 108.210 103.835 108.665 ;
        RECT 104.435 108.210 104.695 108.665 ;
        RECT 105.295 108.210 105.555 108.665 ;
        RECT 106.140 108.210 106.415 108.665 ;
        RECT 107.000 108.210 107.260 108.665 ;
        RECT 107.860 108.210 108.120 108.665 ;
        RECT 108.720 108.210 108.980 108.665 ;
        RECT 109.580 108.195 109.830 109.005 ;
        RECT 110.440 108.195 110.690 109.005 ;
        RECT 110.860 108.695 111.175 109.255 ;
        RECT 111.365 108.915 111.695 109.285 ;
        RECT 111.930 108.990 112.215 109.320 ;
        RECT 111.930 108.735 112.100 108.990 ;
        RECT 111.435 108.565 112.100 108.735 ;
        RECT 112.385 108.690 112.555 109.490 ;
        RECT 112.815 109.635 112.985 110.395 ;
        RECT 112.815 109.465 113.480 109.635 ;
        RECT 113.665 109.490 113.935 110.395 ;
        RECT 113.310 109.320 113.480 109.465 ;
        RECT 112.745 108.915 113.075 109.285 ;
        RECT 113.310 108.990 113.595 109.320 ;
        RECT 113.310 108.735 113.480 108.990 ;
        RECT 111.435 108.185 111.605 108.565 ;
        RECT 112.295 108.185 112.555 108.690 ;
        RECT 112.815 108.565 113.480 108.735 ;
        RECT 113.765 108.690 113.935 109.490 ;
        RECT 114.655 109.635 114.825 110.395 ;
        RECT 114.655 109.465 115.320 109.635 ;
        RECT 115.505 109.490 115.775 110.395 ;
        RECT 115.150 109.320 115.320 109.465 ;
        RECT 114.585 108.915 114.915 109.285 ;
        RECT 115.150 108.990 115.435 109.320 ;
        RECT 115.150 108.735 115.320 108.990 ;
        RECT 112.815 108.185 112.985 108.565 ;
        RECT 113.675 108.185 113.935 108.690 ;
        RECT 114.655 108.565 115.320 108.735 ;
        RECT 115.605 108.690 115.775 109.490 ;
        RECT 116.385 109.415 116.715 110.395 ;
        RECT 115.965 109.005 116.295 109.255 ;
        RECT 116.465 108.815 116.715 109.415 ;
        RECT 114.655 108.185 114.825 108.565 ;
        RECT 115.515 108.185 115.775 108.690 ;
        RECT 116.385 108.185 116.715 108.815 ;
        RECT 117.330 109.375 117.585 110.255 ;
        RECT 118.910 110.015 119.080 110.305 ;
        RECT 118.280 109.845 119.080 110.015 ;
        RECT 119.670 110.055 120.540 110.395 ;
        RECT 117.330 108.725 117.540 109.375 ;
        RECT 118.280 109.255 118.450 109.845 ;
        RECT 119.670 109.675 119.840 110.055 ;
        RECT 120.775 109.935 120.945 110.395 ;
        RECT 121.780 109.965 121.950 110.305 ;
        RECT 122.685 109.965 122.855 110.305 ;
        RECT 118.620 109.505 119.840 109.675 ;
        RECT 120.010 109.595 120.470 109.885 ;
        RECT 120.775 109.765 121.335 109.935 ;
        RECT 121.780 109.795 122.855 109.965 ;
        RECT 123.025 110.065 123.705 110.395 ;
        RECT 123.920 110.065 124.170 110.395 ;
        RECT 121.165 109.625 121.335 109.765 ;
        RECT 120.010 109.585 120.975 109.595 ;
        RECT 119.670 109.415 119.840 109.505 ;
        RECT 120.300 109.425 120.975 109.585 ;
        RECT 117.710 109.225 118.450 109.255 ;
        RECT 117.710 108.925 118.625 109.225 ;
        RECT 118.300 108.750 118.625 108.925 ;
        RECT 117.330 108.195 117.585 108.725 ;
        RECT 118.305 108.395 118.625 108.750 ;
        RECT 118.795 108.965 119.335 109.335 ;
        RECT 119.670 109.245 120.075 109.415 ;
        RECT 118.795 108.565 119.035 108.965 ;
        RECT 119.515 108.795 119.735 109.075 ;
        RECT 119.205 108.625 119.735 108.795 ;
        RECT 119.205 108.395 119.375 108.625 ;
        RECT 118.305 108.225 119.375 108.395 ;
        RECT 119.905 108.465 120.075 109.245 ;
        RECT 120.245 108.635 120.595 109.255 ;
        RECT 120.765 108.635 120.975 109.425 ;
        RECT 121.165 109.455 122.665 109.625 ;
        RECT 121.165 108.765 121.335 109.455 ;
        RECT 123.025 109.285 123.195 110.065 ;
        RECT 124.000 109.935 124.170 110.065 ;
        RECT 121.505 109.115 123.195 109.285 ;
        RECT 123.365 109.505 123.830 109.895 ;
        RECT 124.000 109.765 124.395 109.935 ;
        RECT 121.505 108.935 121.675 109.115 ;
        RECT 119.905 108.185 120.855 108.465 ;
        RECT 121.165 108.375 121.425 108.765 ;
        RECT 121.845 108.695 122.635 108.945 ;
        RECT 121.075 108.205 121.425 108.375 ;
        RECT 122.840 108.405 123.010 109.115 ;
        RECT 123.365 108.915 123.535 109.505 ;
        RECT 123.180 108.695 123.535 108.915 ;
        RECT 123.705 108.695 124.055 109.315 ;
        RECT 124.225 108.405 124.395 109.765 ;
        RECT 124.760 109.595 125.085 110.380 ;
        RECT 124.565 108.545 125.025 109.595 ;
        RECT 122.840 108.235 123.695 108.405 ;
        RECT 123.900 108.235 124.395 108.405 ;
        RECT 125.255 108.275 125.425 110.395 ;
        RECT 126.095 109.895 126.350 110.395 ;
        RECT 125.600 109.725 126.350 109.895 ;
        RECT 125.600 108.735 125.830 109.725 ;
        RECT 126.000 108.905 126.350 109.555 ;
        RECT 125.600 108.565 126.350 108.735 ;
        RECT 126.095 108.275 126.350 108.565 ;
        RECT 17.945 107.045 18.275 107.675 ;
        RECT 18.890 107.135 19.145 107.665 ;
        RECT 19.865 107.465 20.935 107.635 ;
        RECT 17.945 106.445 18.195 107.045 ;
        RECT 18.365 106.605 18.695 106.855 ;
        RECT 18.890 106.485 19.100 107.135 ;
        RECT 19.865 107.110 20.185 107.465 ;
        RECT 19.860 106.935 20.185 107.110 ;
        RECT 19.270 106.635 20.185 106.935 ;
        RECT 20.355 106.895 20.595 107.295 ;
        RECT 20.765 107.235 20.935 107.465 ;
        RECT 21.465 107.395 22.415 107.675 ;
        RECT 22.635 107.485 22.985 107.655 ;
        RECT 20.765 107.065 21.295 107.235 ;
        RECT 19.270 106.605 20.010 106.635 ;
        RECT 17.945 105.465 18.275 106.445 ;
        RECT 18.890 105.605 19.145 106.485 ;
        RECT 19.840 106.015 20.010 106.605 ;
        RECT 20.355 106.525 20.895 106.895 ;
        RECT 21.075 106.785 21.295 107.065 ;
        RECT 21.465 106.615 21.635 107.395 ;
        RECT 21.230 106.445 21.635 106.615 ;
        RECT 21.805 106.605 22.155 107.225 ;
        RECT 21.230 106.355 21.400 106.445 ;
        RECT 22.325 106.435 22.535 107.225 ;
        RECT 20.180 106.185 21.400 106.355 ;
        RECT 21.860 106.275 22.535 106.435 ;
        RECT 19.840 105.845 20.640 106.015 ;
        RECT 20.470 105.555 20.640 105.845 ;
        RECT 21.230 105.805 21.400 106.185 ;
        RECT 21.570 106.265 22.535 106.275 ;
        RECT 22.725 107.095 22.985 107.485 ;
        RECT 24.400 107.455 25.255 107.625 ;
        RECT 25.460 107.455 25.955 107.625 ;
        RECT 22.725 106.405 22.895 107.095 ;
        RECT 23.065 106.745 23.235 106.925 ;
        RECT 23.405 106.915 24.195 107.165 ;
        RECT 24.400 106.745 24.570 107.455 ;
        RECT 24.740 106.945 25.095 107.165 ;
        RECT 23.065 106.575 24.755 106.745 ;
        RECT 21.570 105.975 22.030 106.265 ;
        RECT 22.725 106.235 24.225 106.405 ;
        RECT 22.725 106.095 22.895 106.235 ;
        RECT 22.335 105.925 22.895 106.095 ;
        RECT 21.230 105.465 22.100 105.805 ;
        RECT 22.335 105.465 22.505 105.925 ;
        RECT 23.340 105.895 24.415 106.065 ;
        RECT 23.340 105.555 23.510 105.895 ;
        RECT 24.245 105.555 24.415 105.895 ;
        RECT 24.585 105.795 24.755 106.575 ;
        RECT 24.925 106.355 25.095 106.945 ;
        RECT 25.265 106.545 25.615 107.165 ;
        RECT 24.925 105.965 25.390 106.355 ;
        RECT 25.785 106.095 25.955 107.455 ;
        RECT 26.125 106.265 26.585 107.315 ;
        RECT 25.560 105.925 25.955 106.095 ;
        RECT 25.560 105.795 25.730 105.925 ;
        RECT 24.585 105.465 25.265 105.795 ;
        RECT 25.480 105.465 25.730 105.795 ;
        RECT 26.320 105.480 26.645 106.265 ;
        RECT 26.815 105.465 26.985 107.585 ;
        RECT 27.655 107.295 27.910 107.585 ;
        RECT 27.160 107.125 27.910 107.295 ;
        RECT 28.090 107.135 28.345 107.665 ;
        RECT 29.065 107.465 30.135 107.635 ;
        RECT 27.160 106.135 27.390 107.125 ;
        RECT 27.560 106.305 27.910 106.955 ;
        RECT 28.090 106.485 28.300 107.135 ;
        RECT 29.065 107.110 29.385 107.465 ;
        RECT 29.060 106.935 29.385 107.110 ;
        RECT 28.470 106.635 29.385 106.935 ;
        RECT 29.555 106.895 29.795 107.295 ;
        RECT 29.965 107.235 30.135 107.465 ;
        RECT 30.665 107.395 31.615 107.675 ;
        RECT 31.835 107.485 32.185 107.655 ;
        RECT 29.965 107.065 30.495 107.235 ;
        RECT 28.470 106.605 29.210 106.635 ;
        RECT 27.160 105.965 27.910 106.135 ;
        RECT 27.655 105.465 27.910 105.965 ;
        RECT 28.090 105.605 28.345 106.485 ;
        RECT 29.040 106.015 29.210 106.605 ;
        RECT 29.555 106.525 30.095 106.895 ;
        RECT 30.275 106.785 30.495 107.065 ;
        RECT 30.665 106.615 30.835 107.395 ;
        RECT 30.430 106.445 30.835 106.615 ;
        RECT 31.005 106.605 31.355 107.225 ;
        RECT 30.430 106.355 30.600 106.445 ;
        RECT 31.525 106.435 31.735 107.225 ;
        RECT 29.380 106.185 30.600 106.355 ;
        RECT 31.060 106.275 31.735 106.435 ;
        RECT 29.040 105.845 29.840 106.015 ;
        RECT 29.670 105.555 29.840 105.845 ;
        RECT 30.430 105.805 30.600 106.185 ;
        RECT 30.770 106.265 31.735 106.275 ;
        RECT 31.925 107.095 32.185 107.485 ;
        RECT 33.600 107.455 34.455 107.625 ;
        RECT 34.660 107.455 35.155 107.625 ;
        RECT 31.925 106.405 32.095 107.095 ;
        RECT 32.265 106.745 32.435 106.925 ;
        RECT 32.605 106.915 33.395 107.165 ;
        RECT 33.600 106.745 33.770 107.455 ;
        RECT 33.940 106.945 34.295 107.165 ;
        RECT 32.265 106.575 33.955 106.745 ;
        RECT 30.770 105.975 31.230 106.265 ;
        RECT 31.925 106.235 33.425 106.405 ;
        RECT 31.925 106.095 32.095 106.235 ;
        RECT 31.535 105.925 32.095 106.095 ;
        RECT 30.430 105.465 31.300 105.805 ;
        RECT 31.535 105.465 31.705 105.925 ;
        RECT 32.540 105.895 33.615 106.065 ;
        RECT 32.540 105.555 32.710 105.895 ;
        RECT 33.445 105.555 33.615 105.895 ;
        RECT 33.785 105.795 33.955 106.575 ;
        RECT 34.125 106.355 34.295 106.945 ;
        RECT 34.465 106.545 34.815 107.165 ;
        RECT 34.125 105.965 34.590 106.355 ;
        RECT 34.985 106.095 35.155 107.455 ;
        RECT 35.325 106.265 35.785 107.315 ;
        RECT 34.760 105.925 35.155 106.095 ;
        RECT 34.760 105.795 34.930 105.925 ;
        RECT 33.785 105.465 34.465 105.795 ;
        RECT 34.680 105.465 34.930 105.795 ;
        RECT 35.520 105.480 35.845 106.265 ;
        RECT 36.015 105.465 36.185 107.585 ;
        RECT 36.855 107.295 37.110 107.585 ;
        RECT 36.360 107.125 37.110 107.295 ;
        RECT 36.360 106.135 36.590 107.125 ;
        RECT 38.185 107.045 38.515 107.675 ;
        RECT 39.685 107.195 39.945 107.650 ;
        RECT 40.555 107.195 40.815 107.650 ;
        RECT 41.415 107.195 41.675 107.650 ;
        RECT 42.275 107.195 42.535 107.650 ;
        RECT 43.120 107.195 43.395 107.650 ;
        RECT 43.980 107.195 44.240 107.650 ;
        RECT 44.840 107.195 45.100 107.650 ;
        RECT 45.700 107.195 45.960 107.650 ;
        RECT 36.760 106.305 37.110 106.955 ;
        RECT 37.765 106.605 38.095 106.855 ;
        RECT 38.265 106.445 38.515 107.045 ;
        RECT 36.360 105.965 37.110 106.135 ;
        RECT 36.855 105.465 37.110 105.965 ;
        RECT 38.185 105.465 38.515 106.445 ;
        RECT 39.215 107.025 45.960 107.195 ;
        RECT 39.215 106.435 40.380 107.025 ;
        RECT 46.560 106.855 46.810 107.665 ;
        RECT 47.420 106.855 47.670 107.665 ;
        RECT 40.550 106.605 47.670 106.855 ;
        RECT 47.840 106.605 48.155 107.165 ;
        RECT 48.330 107.135 48.585 107.665 ;
        RECT 49.305 107.465 50.375 107.635 ;
        RECT 39.215 106.210 45.960 106.435 ;
        RECT 39.655 105.470 39.945 106.210 ;
        RECT 40.555 106.195 45.960 106.210 ;
        RECT 40.555 105.470 40.815 106.195 ;
        RECT 41.415 105.470 41.675 106.195 ;
        RECT 42.275 105.470 42.535 106.195 ;
        RECT 43.120 105.470 43.380 106.195 ;
        RECT 43.980 105.470 44.240 106.195 ;
        RECT 44.840 105.470 45.100 106.195 ;
        RECT 45.700 105.470 45.960 106.195 ;
        RECT 46.560 105.470 46.810 106.605 ;
        RECT 47.425 105.465 47.670 106.605 ;
        RECT 48.330 106.485 48.540 107.135 ;
        RECT 49.305 107.110 49.625 107.465 ;
        RECT 49.300 106.935 49.625 107.110 ;
        RECT 48.710 106.635 49.625 106.935 ;
        RECT 49.795 106.895 50.035 107.295 ;
        RECT 50.205 107.235 50.375 107.465 ;
        RECT 50.905 107.395 51.855 107.675 ;
        RECT 52.075 107.485 52.425 107.655 ;
        RECT 50.205 107.065 50.735 107.235 ;
        RECT 48.710 106.605 49.450 106.635 ;
        RECT 48.330 105.605 48.585 106.485 ;
        RECT 49.280 106.015 49.450 106.605 ;
        RECT 49.795 106.525 50.335 106.895 ;
        RECT 50.515 106.785 50.735 107.065 ;
        RECT 50.905 106.615 51.075 107.395 ;
        RECT 50.670 106.445 51.075 106.615 ;
        RECT 51.245 106.605 51.595 107.225 ;
        RECT 50.670 106.355 50.840 106.445 ;
        RECT 51.765 106.435 51.975 107.225 ;
        RECT 49.620 106.185 50.840 106.355 ;
        RECT 51.300 106.275 51.975 106.435 ;
        RECT 49.280 105.845 50.080 106.015 ;
        RECT 49.910 105.555 50.080 105.845 ;
        RECT 50.670 105.805 50.840 106.185 ;
        RECT 51.010 106.265 51.975 106.275 ;
        RECT 52.165 107.095 52.425 107.485 ;
        RECT 53.840 107.455 54.695 107.625 ;
        RECT 54.900 107.455 55.395 107.625 ;
        RECT 52.165 106.405 52.335 107.095 ;
        RECT 52.505 106.745 52.675 106.925 ;
        RECT 52.845 106.915 53.635 107.165 ;
        RECT 53.840 106.745 54.010 107.455 ;
        RECT 54.180 106.945 54.535 107.165 ;
        RECT 52.505 106.575 54.195 106.745 ;
        RECT 51.010 105.975 51.470 106.265 ;
        RECT 52.165 106.235 53.665 106.405 ;
        RECT 52.165 106.095 52.335 106.235 ;
        RECT 51.775 105.925 52.335 106.095 ;
        RECT 50.670 105.465 51.540 105.805 ;
        RECT 51.775 105.465 51.945 105.925 ;
        RECT 52.780 105.895 53.855 106.065 ;
        RECT 52.780 105.555 52.950 105.895 ;
        RECT 53.685 105.555 53.855 105.895 ;
        RECT 54.025 105.795 54.195 106.575 ;
        RECT 54.365 106.355 54.535 106.945 ;
        RECT 54.705 106.545 55.055 107.165 ;
        RECT 54.365 105.965 54.830 106.355 ;
        RECT 55.225 106.095 55.395 107.455 ;
        RECT 55.565 106.265 56.025 107.315 ;
        RECT 55.000 105.925 55.395 106.095 ;
        RECT 55.000 105.795 55.170 105.925 ;
        RECT 54.025 105.465 54.705 105.795 ;
        RECT 54.920 105.465 55.170 105.795 ;
        RECT 55.760 105.480 56.085 106.265 ;
        RECT 56.255 105.465 56.425 107.585 ;
        RECT 57.095 107.295 57.350 107.585 ;
        RECT 56.600 107.125 57.350 107.295 ;
        RECT 56.600 106.135 56.830 107.125 ;
        RECT 57.965 107.045 58.295 107.675 ;
        RECT 60.725 107.045 61.055 107.675 ;
        RECT 61.755 107.295 61.925 107.675 ;
        RECT 61.755 107.125 62.420 107.295 ;
        RECT 62.615 107.170 62.875 107.675 ;
        RECT 57.000 106.305 57.350 106.955 ;
        RECT 57.965 106.445 58.215 107.045 ;
        RECT 58.385 106.605 58.715 106.855 ;
        RECT 60.305 106.605 60.635 106.855 ;
        RECT 60.805 106.445 61.055 107.045 ;
        RECT 61.685 106.575 62.015 106.945 ;
        RECT 62.250 106.870 62.420 107.125 ;
        RECT 56.600 105.965 57.350 106.135 ;
        RECT 57.095 105.465 57.350 105.965 ;
        RECT 57.965 105.465 58.295 106.445 ;
        RECT 60.725 105.465 61.055 106.445 ;
        RECT 62.250 106.540 62.535 106.870 ;
        RECT 62.250 106.395 62.420 106.540 ;
        RECT 61.755 106.225 62.420 106.395 ;
        RECT 62.705 106.370 62.875 107.170 ;
        RECT 63.945 107.045 64.275 107.675 ;
        RECT 63.525 106.605 63.855 106.855 ;
        RECT 64.025 106.445 64.275 107.045 ;
        RECT 61.755 105.465 61.925 106.225 ;
        RECT 62.605 105.465 62.875 106.370 ;
        RECT 63.945 105.465 64.275 106.445 ;
        RECT 64.890 107.135 65.145 107.665 ;
        RECT 65.865 107.465 66.935 107.635 ;
        RECT 64.890 106.485 65.100 107.135 ;
        RECT 65.865 107.110 66.185 107.465 ;
        RECT 65.860 106.935 66.185 107.110 ;
        RECT 65.270 106.635 66.185 106.935 ;
        RECT 66.355 106.895 66.595 107.295 ;
        RECT 66.765 107.235 66.935 107.465 ;
        RECT 67.465 107.395 68.415 107.675 ;
        RECT 68.635 107.485 68.985 107.655 ;
        RECT 66.765 107.065 67.295 107.235 ;
        RECT 65.270 106.605 66.010 106.635 ;
        RECT 64.890 105.605 65.145 106.485 ;
        RECT 65.840 106.015 66.010 106.605 ;
        RECT 66.355 106.525 66.895 106.895 ;
        RECT 67.075 106.785 67.295 107.065 ;
        RECT 67.465 106.615 67.635 107.395 ;
        RECT 67.230 106.445 67.635 106.615 ;
        RECT 67.805 106.605 68.155 107.225 ;
        RECT 67.230 106.355 67.400 106.445 ;
        RECT 68.325 106.435 68.535 107.225 ;
        RECT 66.180 106.185 67.400 106.355 ;
        RECT 67.860 106.275 68.535 106.435 ;
        RECT 65.840 105.845 66.640 106.015 ;
        RECT 66.470 105.555 66.640 105.845 ;
        RECT 67.230 105.805 67.400 106.185 ;
        RECT 67.570 106.265 68.535 106.275 ;
        RECT 68.725 107.095 68.985 107.485 ;
        RECT 70.400 107.455 71.255 107.625 ;
        RECT 71.460 107.455 71.955 107.625 ;
        RECT 68.725 106.405 68.895 107.095 ;
        RECT 69.065 106.745 69.235 106.925 ;
        RECT 69.405 106.915 70.195 107.165 ;
        RECT 70.400 106.745 70.570 107.455 ;
        RECT 70.740 106.945 71.095 107.165 ;
        RECT 69.065 106.575 70.755 106.745 ;
        RECT 67.570 105.975 68.030 106.265 ;
        RECT 68.725 106.235 70.225 106.405 ;
        RECT 68.725 106.095 68.895 106.235 ;
        RECT 68.335 105.925 68.895 106.095 ;
        RECT 67.230 105.465 68.100 105.805 ;
        RECT 68.335 105.465 68.505 105.925 ;
        RECT 69.340 105.895 70.415 106.065 ;
        RECT 69.340 105.555 69.510 105.895 ;
        RECT 70.245 105.555 70.415 105.895 ;
        RECT 70.585 105.795 70.755 106.575 ;
        RECT 70.925 106.355 71.095 106.945 ;
        RECT 71.265 106.545 71.615 107.165 ;
        RECT 70.925 105.965 71.390 106.355 ;
        RECT 71.785 106.095 71.955 107.455 ;
        RECT 72.125 106.265 72.585 107.315 ;
        RECT 71.560 105.925 71.955 106.095 ;
        RECT 71.560 105.795 71.730 105.925 ;
        RECT 70.585 105.465 71.265 105.795 ;
        RECT 71.480 105.465 71.730 105.795 ;
        RECT 72.320 105.480 72.645 106.265 ;
        RECT 72.815 105.465 72.985 107.585 ;
        RECT 73.655 107.295 73.910 107.585 ;
        RECT 73.160 107.125 73.910 107.295 ;
        RECT 73.160 106.135 73.390 107.125 ;
        RECT 75.445 107.045 75.775 107.675 ;
        RECT 76.475 107.295 76.645 107.675 ;
        RECT 76.475 107.125 77.140 107.295 ;
        RECT 77.335 107.170 77.595 107.675 ;
        RECT 73.560 106.305 73.910 106.955 ;
        RECT 75.445 106.445 75.695 107.045 ;
        RECT 75.865 106.605 76.195 106.855 ;
        RECT 76.405 106.575 76.735 106.945 ;
        RECT 76.970 106.870 77.140 107.125 ;
        RECT 76.970 106.540 77.255 106.870 ;
        RECT 73.160 105.965 73.910 106.135 ;
        RECT 73.655 105.465 73.910 105.965 ;
        RECT 75.445 105.465 75.775 106.445 ;
        RECT 76.970 106.395 77.140 106.540 ;
        RECT 76.475 106.225 77.140 106.395 ;
        RECT 77.425 106.370 77.595 107.170 ;
        RECT 76.475 105.465 76.645 106.225 ;
        RECT 77.325 105.465 77.595 106.370 ;
        RECT 77.770 107.135 78.025 107.665 ;
        RECT 78.745 107.465 79.815 107.635 ;
        RECT 77.770 106.485 77.980 107.135 ;
        RECT 78.745 107.110 79.065 107.465 ;
        RECT 78.740 106.935 79.065 107.110 ;
        RECT 78.150 106.635 79.065 106.935 ;
        RECT 79.235 106.895 79.475 107.295 ;
        RECT 79.645 107.235 79.815 107.465 ;
        RECT 80.345 107.395 81.295 107.675 ;
        RECT 81.515 107.485 81.865 107.655 ;
        RECT 79.645 107.065 80.175 107.235 ;
        RECT 78.150 106.605 78.890 106.635 ;
        RECT 77.770 105.605 78.025 106.485 ;
        RECT 78.720 106.015 78.890 106.605 ;
        RECT 79.235 106.525 79.775 106.895 ;
        RECT 79.955 106.785 80.175 107.065 ;
        RECT 80.345 106.615 80.515 107.395 ;
        RECT 80.110 106.445 80.515 106.615 ;
        RECT 80.685 106.605 81.035 107.225 ;
        RECT 80.110 106.355 80.280 106.445 ;
        RECT 81.205 106.435 81.415 107.225 ;
        RECT 79.060 106.185 80.280 106.355 ;
        RECT 80.740 106.275 81.415 106.435 ;
        RECT 78.720 105.845 79.520 106.015 ;
        RECT 79.350 105.555 79.520 105.845 ;
        RECT 80.110 105.805 80.280 106.185 ;
        RECT 80.450 106.265 81.415 106.275 ;
        RECT 81.605 107.095 81.865 107.485 ;
        RECT 83.280 107.455 84.135 107.625 ;
        RECT 84.340 107.455 84.835 107.625 ;
        RECT 81.605 106.405 81.775 107.095 ;
        RECT 81.945 106.745 82.115 106.925 ;
        RECT 82.285 106.915 83.075 107.165 ;
        RECT 83.280 106.745 83.450 107.455 ;
        RECT 83.620 106.945 83.975 107.165 ;
        RECT 81.945 106.575 83.635 106.745 ;
        RECT 80.450 105.975 80.910 106.265 ;
        RECT 81.605 106.235 83.105 106.405 ;
        RECT 81.605 106.095 81.775 106.235 ;
        RECT 81.215 105.925 81.775 106.095 ;
        RECT 80.110 105.465 80.980 105.805 ;
        RECT 81.215 105.465 81.385 105.925 ;
        RECT 82.220 105.895 83.295 106.065 ;
        RECT 82.220 105.555 82.390 105.895 ;
        RECT 83.125 105.555 83.295 105.895 ;
        RECT 83.465 105.795 83.635 106.575 ;
        RECT 83.805 106.355 83.975 106.945 ;
        RECT 84.145 106.545 84.495 107.165 ;
        RECT 83.805 105.965 84.270 106.355 ;
        RECT 84.665 106.095 84.835 107.455 ;
        RECT 85.005 106.265 85.465 107.315 ;
        RECT 84.440 105.925 84.835 106.095 ;
        RECT 84.440 105.795 84.610 105.925 ;
        RECT 83.465 105.465 84.145 105.795 ;
        RECT 84.360 105.465 84.610 105.795 ;
        RECT 85.200 105.480 85.525 106.265 ;
        RECT 85.695 105.465 85.865 107.585 ;
        RECT 86.535 107.295 86.790 107.585 ;
        RECT 86.040 107.125 86.790 107.295 ;
        RECT 86.965 107.170 87.225 107.675 ;
        RECT 87.915 107.295 88.085 107.675 ;
        RECT 86.040 106.135 86.270 107.125 ;
        RECT 86.440 106.305 86.790 106.955 ;
        RECT 86.965 106.370 87.135 107.170 ;
        RECT 87.420 107.125 88.085 107.295 ;
        RECT 90.190 107.135 90.445 107.665 ;
        RECT 91.165 107.465 92.235 107.635 ;
        RECT 87.420 106.870 87.590 107.125 ;
        RECT 87.305 106.540 87.590 106.870 ;
        RECT 87.825 106.575 88.155 106.945 ;
        RECT 87.420 106.395 87.590 106.540 ;
        RECT 90.190 106.485 90.400 107.135 ;
        RECT 91.165 107.110 91.485 107.465 ;
        RECT 91.160 106.935 91.485 107.110 ;
        RECT 90.570 106.635 91.485 106.935 ;
        RECT 91.655 106.895 91.895 107.295 ;
        RECT 92.065 107.235 92.235 107.465 ;
        RECT 92.765 107.395 93.715 107.675 ;
        RECT 93.935 107.485 94.285 107.655 ;
        RECT 92.065 107.065 92.595 107.235 ;
        RECT 90.570 106.605 91.310 106.635 ;
        RECT 86.040 105.965 86.790 106.135 ;
        RECT 86.535 105.465 86.790 105.965 ;
        RECT 86.965 105.465 87.235 106.370 ;
        RECT 87.420 106.225 88.085 106.395 ;
        RECT 87.915 105.465 88.085 106.225 ;
        RECT 90.190 105.605 90.445 106.485 ;
        RECT 91.140 106.015 91.310 106.605 ;
        RECT 91.655 106.525 92.195 106.895 ;
        RECT 92.375 106.785 92.595 107.065 ;
        RECT 92.765 106.615 92.935 107.395 ;
        RECT 92.530 106.445 92.935 106.615 ;
        RECT 93.105 106.605 93.455 107.225 ;
        RECT 92.530 106.355 92.700 106.445 ;
        RECT 93.625 106.435 93.835 107.225 ;
        RECT 91.480 106.185 92.700 106.355 ;
        RECT 93.160 106.275 93.835 106.435 ;
        RECT 91.140 105.845 91.940 106.015 ;
        RECT 91.770 105.555 91.940 105.845 ;
        RECT 92.530 105.805 92.700 106.185 ;
        RECT 92.870 106.265 93.835 106.275 ;
        RECT 94.025 107.095 94.285 107.485 ;
        RECT 95.700 107.455 96.555 107.625 ;
        RECT 96.760 107.455 97.255 107.625 ;
        RECT 94.025 106.405 94.195 107.095 ;
        RECT 94.365 106.745 94.535 106.925 ;
        RECT 94.705 106.915 95.495 107.165 ;
        RECT 95.700 106.745 95.870 107.455 ;
        RECT 96.040 106.945 96.395 107.165 ;
        RECT 94.365 106.575 96.055 106.745 ;
        RECT 92.870 105.975 93.330 106.265 ;
        RECT 94.025 106.235 95.525 106.405 ;
        RECT 94.025 106.095 94.195 106.235 ;
        RECT 93.635 105.925 94.195 106.095 ;
        RECT 92.530 105.465 93.400 105.805 ;
        RECT 93.635 105.465 93.805 105.925 ;
        RECT 94.640 105.895 95.715 106.065 ;
        RECT 94.640 105.555 94.810 105.895 ;
        RECT 95.545 105.555 95.715 105.895 ;
        RECT 95.885 105.795 96.055 106.575 ;
        RECT 96.225 106.355 96.395 106.945 ;
        RECT 96.565 106.545 96.915 107.165 ;
        RECT 96.225 105.965 96.690 106.355 ;
        RECT 97.085 106.095 97.255 107.455 ;
        RECT 97.425 106.265 97.885 107.315 ;
        RECT 96.860 105.925 97.255 106.095 ;
        RECT 96.860 105.795 97.030 105.925 ;
        RECT 95.885 105.465 96.565 105.795 ;
        RECT 96.780 105.465 97.030 105.795 ;
        RECT 97.620 105.480 97.945 106.265 ;
        RECT 98.115 105.465 98.285 107.585 ;
        RECT 98.955 107.295 99.210 107.585 ;
        RECT 98.460 107.125 99.210 107.295 ;
        RECT 99.390 107.135 99.645 107.665 ;
        RECT 100.365 107.465 101.435 107.635 ;
        RECT 98.460 106.135 98.690 107.125 ;
        RECT 98.860 106.305 99.210 106.955 ;
        RECT 99.390 106.485 99.600 107.135 ;
        RECT 100.365 107.110 100.685 107.465 ;
        RECT 100.360 106.935 100.685 107.110 ;
        RECT 99.770 106.635 100.685 106.935 ;
        RECT 100.855 106.895 101.095 107.295 ;
        RECT 101.265 107.235 101.435 107.465 ;
        RECT 101.965 107.395 102.915 107.675 ;
        RECT 103.135 107.485 103.485 107.655 ;
        RECT 101.265 107.065 101.795 107.235 ;
        RECT 99.770 106.605 100.510 106.635 ;
        RECT 98.460 105.965 99.210 106.135 ;
        RECT 98.955 105.465 99.210 105.965 ;
        RECT 99.390 105.605 99.645 106.485 ;
        RECT 100.340 106.015 100.510 106.605 ;
        RECT 100.855 106.525 101.395 106.895 ;
        RECT 101.575 106.785 101.795 107.065 ;
        RECT 101.965 106.615 102.135 107.395 ;
        RECT 101.730 106.445 102.135 106.615 ;
        RECT 102.305 106.605 102.655 107.225 ;
        RECT 101.730 106.355 101.900 106.445 ;
        RECT 102.825 106.435 103.035 107.225 ;
        RECT 100.680 106.185 101.900 106.355 ;
        RECT 102.360 106.275 103.035 106.435 ;
        RECT 100.340 105.845 101.140 106.015 ;
        RECT 100.970 105.555 101.140 105.845 ;
        RECT 101.730 105.805 101.900 106.185 ;
        RECT 102.070 106.265 103.035 106.275 ;
        RECT 103.225 107.095 103.485 107.485 ;
        RECT 104.900 107.455 105.755 107.625 ;
        RECT 105.960 107.455 106.455 107.625 ;
        RECT 103.225 106.405 103.395 107.095 ;
        RECT 103.565 106.745 103.735 106.925 ;
        RECT 103.905 106.915 104.695 107.165 ;
        RECT 104.900 106.745 105.070 107.455 ;
        RECT 105.240 106.945 105.595 107.165 ;
        RECT 103.565 106.575 105.255 106.745 ;
        RECT 102.070 105.975 102.530 106.265 ;
        RECT 103.225 106.235 104.725 106.405 ;
        RECT 103.225 106.095 103.395 106.235 ;
        RECT 102.835 105.925 103.395 106.095 ;
        RECT 101.730 105.465 102.600 105.805 ;
        RECT 102.835 105.465 103.005 105.925 ;
        RECT 103.840 105.895 104.915 106.065 ;
        RECT 103.840 105.555 104.010 105.895 ;
        RECT 104.745 105.555 104.915 105.895 ;
        RECT 105.085 105.795 105.255 106.575 ;
        RECT 105.425 106.355 105.595 106.945 ;
        RECT 105.765 106.545 106.115 107.165 ;
        RECT 105.425 105.965 105.890 106.355 ;
        RECT 106.285 106.095 106.455 107.455 ;
        RECT 106.625 106.265 107.085 107.315 ;
        RECT 106.060 105.925 106.455 106.095 ;
        RECT 106.060 105.795 106.230 105.925 ;
        RECT 105.085 105.465 105.765 105.795 ;
        RECT 105.980 105.465 106.230 105.795 ;
        RECT 106.820 105.480 107.145 106.265 ;
        RECT 107.315 105.465 107.485 107.585 ;
        RECT 108.155 107.295 108.410 107.585 ;
        RECT 107.660 107.125 108.410 107.295 ;
        RECT 107.660 106.135 107.890 107.125 ;
        RECT 109.025 107.045 109.355 107.675 ;
        RECT 110.405 107.045 110.735 107.675 ;
        RECT 113.625 107.045 113.955 107.675 ;
        RECT 108.060 106.305 108.410 106.955 ;
        RECT 109.025 106.445 109.275 107.045 ;
        RECT 109.445 106.605 109.775 106.855 ;
        RECT 109.985 106.605 110.315 106.855 ;
        RECT 110.485 106.445 110.735 107.045 ;
        RECT 113.205 106.605 113.535 106.855 ;
        RECT 113.705 106.445 113.955 107.045 ;
        RECT 107.660 105.965 108.410 106.135 ;
        RECT 108.155 105.465 108.410 105.965 ;
        RECT 109.025 105.465 109.355 106.445 ;
        RECT 110.405 105.465 110.735 106.445 ;
        RECT 113.625 105.465 113.955 106.445 ;
        RECT 115.030 107.135 115.285 107.665 ;
        RECT 116.005 107.465 117.075 107.635 ;
        RECT 115.030 106.485 115.240 107.135 ;
        RECT 116.005 107.110 116.325 107.465 ;
        RECT 116.000 106.935 116.325 107.110 ;
        RECT 115.410 106.635 116.325 106.935 ;
        RECT 116.495 106.895 116.735 107.295 ;
        RECT 116.905 107.235 117.075 107.465 ;
        RECT 117.605 107.395 118.555 107.675 ;
        RECT 118.775 107.485 119.125 107.655 ;
        RECT 116.905 107.065 117.435 107.235 ;
        RECT 115.410 106.605 116.150 106.635 ;
        RECT 115.030 105.605 115.285 106.485 ;
        RECT 115.980 106.015 116.150 106.605 ;
        RECT 116.495 106.525 117.035 106.895 ;
        RECT 117.215 106.785 117.435 107.065 ;
        RECT 117.605 106.615 117.775 107.395 ;
        RECT 117.370 106.445 117.775 106.615 ;
        RECT 117.945 106.605 118.295 107.225 ;
        RECT 117.370 106.355 117.540 106.445 ;
        RECT 118.465 106.435 118.675 107.225 ;
        RECT 116.320 106.185 117.540 106.355 ;
        RECT 118.000 106.275 118.675 106.435 ;
        RECT 115.980 105.845 116.780 106.015 ;
        RECT 116.610 105.555 116.780 105.845 ;
        RECT 117.370 105.805 117.540 106.185 ;
        RECT 117.710 106.265 118.675 106.275 ;
        RECT 118.865 107.095 119.125 107.485 ;
        RECT 120.540 107.455 121.395 107.625 ;
        RECT 121.600 107.455 122.095 107.625 ;
        RECT 118.865 106.405 119.035 107.095 ;
        RECT 119.205 106.745 119.375 106.925 ;
        RECT 119.545 106.915 120.335 107.165 ;
        RECT 120.540 106.745 120.710 107.455 ;
        RECT 120.880 106.945 121.235 107.165 ;
        RECT 119.205 106.575 120.895 106.745 ;
        RECT 117.710 105.975 118.170 106.265 ;
        RECT 118.865 106.235 120.365 106.405 ;
        RECT 118.865 106.095 119.035 106.235 ;
        RECT 118.475 105.925 119.035 106.095 ;
        RECT 117.370 105.465 118.240 105.805 ;
        RECT 118.475 105.465 118.645 105.925 ;
        RECT 119.480 105.895 120.555 106.065 ;
        RECT 119.480 105.555 119.650 105.895 ;
        RECT 120.385 105.555 120.555 105.895 ;
        RECT 120.725 105.795 120.895 106.575 ;
        RECT 121.065 106.355 121.235 106.945 ;
        RECT 121.405 106.545 121.755 107.165 ;
        RECT 121.065 105.965 121.530 106.355 ;
        RECT 121.925 106.095 122.095 107.455 ;
        RECT 122.265 106.265 122.725 107.315 ;
        RECT 121.700 105.925 122.095 106.095 ;
        RECT 121.700 105.795 121.870 105.925 ;
        RECT 120.725 105.465 121.405 105.795 ;
        RECT 121.620 105.465 121.870 105.795 ;
        RECT 122.460 105.480 122.785 106.265 ;
        RECT 122.955 105.465 123.125 107.585 ;
        RECT 123.795 107.295 124.050 107.585 ;
        RECT 123.300 107.125 124.050 107.295 ;
        RECT 123.300 106.135 123.530 107.125 ;
        RECT 124.665 107.045 124.995 107.675 ;
        RECT 123.700 106.305 124.050 106.955 ;
        RECT 124.245 106.605 124.575 106.855 ;
        RECT 124.745 106.445 124.995 107.045 ;
        RECT 123.300 105.965 124.050 106.135 ;
        RECT 123.795 105.465 124.050 105.965 ;
        RECT 124.665 105.465 124.995 106.445 ;
        RECT 26.685 103.975 27.015 104.955 ;
        RECT 28.065 103.975 28.395 104.955 ;
        RECT 26.685 103.375 26.935 103.975 ;
        RECT 27.105 103.565 27.435 103.815 ;
        RECT 27.645 103.565 27.975 103.815 ;
        RECT 28.145 103.375 28.395 103.975 ;
        RECT 26.685 102.745 27.015 103.375 ;
        RECT 28.065 102.745 28.395 103.375 ;
        RECT 29.005 104.050 29.275 104.955 ;
        RECT 29.955 104.195 30.125 104.955 ;
        RECT 29.005 103.250 29.175 104.050 ;
        RECT 29.460 104.025 30.125 104.195 ;
        RECT 30.475 104.195 30.645 104.955 ;
        RECT 30.475 104.025 31.140 104.195 ;
        RECT 31.325 104.050 31.595 104.955 ;
        RECT 29.460 103.880 29.630 104.025 ;
        RECT 29.345 103.550 29.630 103.880 ;
        RECT 30.970 103.880 31.140 104.025 ;
        RECT 29.460 103.295 29.630 103.550 ;
        RECT 29.865 103.475 30.195 103.845 ;
        RECT 30.405 103.475 30.735 103.845 ;
        RECT 30.970 103.550 31.255 103.880 ;
        RECT 30.970 103.295 31.140 103.550 ;
        RECT 29.005 102.745 29.265 103.250 ;
        RECT 29.460 103.125 30.125 103.295 ;
        RECT 29.955 102.745 30.125 103.125 ;
        RECT 30.475 103.125 31.140 103.295 ;
        RECT 31.425 103.250 31.595 104.050 ;
        RECT 30.475 102.745 30.645 103.125 ;
        RECT 31.335 102.745 31.595 103.250 ;
        RECT 31.770 103.935 32.025 104.815 ;
        RECT 33.350 104.575 33.520 104.865 ;
        RECT 32.720 104.405 33.520 104.575 ;
        RECT 34.110 104.615 34.980 104.955 ;
        RECT 31.770 103.285 31.980 103.935 ;
        RECT 32.720 103.815 32.890 104.405 ;
        RECT 34.110 104.235 34.280 104.615 ;
        RECT 35.215 104.495 35.385 104.955 ;
        RECT 36.220 104.525 36.390 104.865 ;
        RECT 37.125 104.525 37.295 104.865 ;
        RECT 33.060 104.065 34.280 104.235 ;
        RECT 34.450 104.155 34.910 104.445 ;
        RECT 35.215 104.325 35.775 104.495 ;
        RECT 36.220 104.355 37.295 104.525 ;
        RECT 37.465 104.625 38.145 104.955 ;
        RECT 38.360 104.625 38.610 104.955 ;
        RECT 35.605 104.185 35.775 104.325 ;
        RECT 34.450 104.145 35.415 104.155 ;
        RECT 34.110 103.975 34.280 104.065 ;
        RECT 34.740 103.985 35.415 104.145 ;
        RECT 32.150 103.785 32.890 103.815 ;
        RECT 32.150 103.485 33.065 103.785 ;
        RECT 32.740 103.310 33.065 103.485 ;
        RECT 31.770 102.755 32.025 103.285 ;
        RECT 32.745 102.955 33.065 103.310 ;
        RECT 33.235 103.525 33.775 103.895 ;
        RECT 34.110 103.805 34.515 103.975 ;
        RECT 33.235 103.125 33.475 103.525 ;
        RECT 33.955 103.355 34.175 103.635 ;
        RECT 33.645 103.185 34.175 103.355 ;
        RECT 33.645 102.955 33.815 103.185 ;
        RECT 32.745 102.785 33.815 102.955 ;
        RECT 34.345 103.025 34.515 103.805 ;
        RECT 34.685 103.195 35.035 103.815 ;
        RECT 35.205 103.195 35.415 103.985 ;
        RECT 35.605 104.015 37.105 104.185 ;
        RECT 35.605 103.325 35.775 104.015 ;
        RECT 37.465 103.845 37.635 104.625 ;
        RECT 38.440 104.495 38.610 104.625 ;
        RECT 35.945 103.675 37.635 103.845 ;
        RECT 37.805 104.065 38.270 104.455 ;
        RECT 38.440 104.325 38.835 104.495 ;
        RECT 35.945 103.495 36.115 103.675 ;
        RECT 34.345 102.745 35.295 103.025 ;
        RECT 35.605 102.935 35.865 103.325 ;
        RECT 36.285 103.255 37.075 103.505 ;
        RECT 35.515 102.765 35.865 102.935 ;
        RECT 37.280 102.965 37.450 103.675 ;
        RECT 37.805 103.475 37.975 104.065 ;
        RECT 37.620 103.255 37.975 103.475 ;
        RECT 38.145 103.255 38.495 103.875 ;
        RECT 38.665 102.965 38.835 104.325 ;
        RECT 39.200 104.155 39.525 104.940 ;
        RECT 39.005 103.105 39.465 104.155 ;
        RECT 37.280 102.795 38.135 102.965 ;
        RECT 38.340 102.795 38.835 102.965 ;
        RECT 39.695 102.835 39.865 104.955 ;
        RECT 40.535 104.455 40.790 104.955 ;
        RECT 40.040 104.285 40.790 104.455 ;
        RECT 40.040 103.295 40.270 104.285 ;
        RECT 40.440 103.465 40.790 104.115 ;
        RECT 40.970 103.935 41.225 104.815 ;
        RECT 42.550 104.575 42.720 104.865 ;
        RECT 41.920 104.405 42.720 104.575 ;
        RECT 43.310 104.615 44.180 104.955 ;
        RECT 40.040 103.125 40.790 103.295 ;
        RECT 40.535 102.835 40.790 103.125 ;
        RECT 40.970 103.285 41.180 103.935 ;
        RECT 41.920 103.815 42.090 104.405 ;
        RECT 43.310 104.235 43.480 104.615 ;
        RECT 44.415 104.495 44.585 104.955 ;
        RECT 45.420 104.525 45.590 104.865 ;
        RECT 46.325 104.525 46.495 104.865 ;
        RECT 42.260 104.065 43.480 104.235 ;
        RECT 43.650 104.155 44.110 104.445 ;
        RECT 44.415 104.325 44.975 104.495 ;
        RECT 45.420 104.355 46.495 104.525 ;
        RECT 46.665 104.625 47.345 104.955 ;
        RECT 47.560 104.625 47.810 104.955 ;
        RECT 44.805 104.185 44.975 104.325 ;
        RECT 43.650 104.145 44.615 104.155 ;
        RECT 43.310 103.975 43.480 104.065 ;
        RECT 43.940 103.985 44.615 104.145 ;
        RECT 41.350 103.785 42.090 103.815 ;
        RECT 41.350 103.485 42.265 103.785 ;
        RECT 41.940 103.310 42.265 103.485 ;
        RECT 40.970 102.755 41.225 103.285 ;
        RECT 41.945 102.955 42.265 103.310 ;
        RECT 42.435 103.525 42.975 103.895 ;
        RECT 43.310 103.805 43.715 103.975 ;
        RECT 42.435 103.125 42.675 103.525 ;
        RECT 43.155 103.355 43.375 103.635 ;
        RECT 42.845 103.185 43.375 103.355 ;
        RECT 42.845 102.955 43.015 103.185 ;
        RECT 41.945 102.785 43.015 102.955 ;
        RECT 43.545 103.025 43.715 103.805 ;
        RECT 43.885 103.195 44.235 103.815 ;
        RECT 44.405 103.195 44.615 103.985 ;
        RECT 44.805 104.015 46.305 104.185 ;
        RECT 44.805 103.325 44.975 104.015 ;
        RECT 46.665 103.845 46.835 104.625 ;
        RECT 47.640 104.495 47.810 104.625 ;
        RECT 45.145 103.675 46.835 103.845 ;
        RECT 47.005 104.065 47.470 104.455 ;
        RECT 47.640 104.325 48.035 104.495 ;
        RECT 45.145 103.495 45.315 103.675 ;
        RECT 43.545 102.745 44.495 103.025 ;
        RECT 44.805 102.935 45.065 103.325 ;
        RECT 45.485 103.255 46.275 103.505 ;
        RECT 44.715 102.765 45.065 102.935 ;
        RECT 46.480 102.965 46.650 103.675 ;
        RECT 47.005 103.475 47.175 104.065 ;
        RECT 46.820 103.255 47.175 103.475 ;
        RECT 47.345 103.255 47.695 103.875 ;
        RECT 47.865 102.965 48.035 104.325 ;
        RECT 48.400 104.155 48.725 104.940 ;
        RECT 48.205 103.105 48.665 104.155 ;
        RECT 46.480 102.795 47.335 102.965 ;
        RECT 47.540 102.795 48.035 102.965 ;
        RECT 48.895 102.835 49.065 104.955 ;
        RECT 49.735 104.455 49.990 104.955 ;
        RECT 49.240 104.285 49.990 104.455 ;
        RECT 49.240 103.295 49.470 104.285 ;
        RECT 49.640 103.465 49.990 104.115 ;
        RECT 51.985 103.975 52.315 104.955 ;
        RECT 51.985 103.375 52.235 103.975 ;
        RECT 54.310 103.935 54.565 104.815 ;
        RECT 55.890 104.575 56.060 104.865 ;
        RECT 55.260 104.405 56.060 104.575 ;
        RECT 56.650 104.615 57.520 104.955 ;
        RECT 52.405 103.565 52.735 103.815 ;
        RECT 49.240 103.125 49.990 103.295 ;
        RECT 49.735 102.835 49.990 103.125 ;
        RECT 51.985 102.745 52.315 103.375 ;
        RECT 54.310 103.285 54.520 103.935 ;
        RECT 55.260 103.815 55.430 104.405 ;
        RECT 56.650 104.235 56.820 104.615 ;
        RECT 57.755 104.495 57.925 104.955 ;
        RECT 58.760 104.525 58.930 104.865 ;
        RECT 59.665 104.525 59.835 104.865 ;
        RECT 55.600 104.065 56.820 104.235 ;
        RECT 56.990 104.155 57.450 104.445 ;
        RECT 57.755 104.325 58.315 104.495 ;
        RECT 58.760 104.355 59.835 104.525 ;
        RECT 60.005 104.625 60.685 104.955 ;
        RECT 60.900 104.625 61.150 104.955 ;
        RECT 58.145 104.185 58.315 104.325 ;
        RECT 56.990 104.145 57.955 104.155 ;
        RECT 56.650 103.975 56.820 104.065 ;
        RECT 57.280 103.985 57.955 104.145 ;
        RECT 54.690 103.785 55.430 103.815 ;
        RECT 54.690 103.485 55.605 103.785 ;
        RECT 55.280 103.310 55.605 103.485 ;
        RECT 54.310 102.755 54.565 103.285 ;
        RECT 55.285 102.955 55.605 103.310 ;
        RECT 55.775 103.525 56.315 103.895 ;
        RECT 56.650 103.805 57.055 103.975 ;
        RECT 55.775 103.125 56.015 103.525 ;
        RECT 56.495 103.355 56.715 103.635 ;
        RECT 56.185 103.185 56.715 103.355 ;
        RECT 56.185 102.955 56.355 103.185 ;
        RECT 55.285 102.785 56.355 102.955 ;
        RECT 56.885 103.025 57.055 103.805 ;
        RECT 57.225 103.195 57.575 103.815 ;
        RECT 57.745 103.195 57.955 103.985 ;
        RECT 58.145 104.015 59.645 104.185 ;
        RECT 58.145 103.325 58.315 104.015 ;
        RECT 60.005 103.845 60.175 104.625 ;
        RECT 60.980 104.495 61.150 104.625 ;
        RECT 58.485 103.675 60.175 103.845 ;
        RECT 60.345 104.065 60.810 104.455 ;
        RECT 60.980 104.325 61.375 104.495 ;
        RECT 58.485 103.495 58.655 103.675 ;
        RECT 56.885 102.745 57.835 103.025 ;
        RECT 58.145 102.935 58.405 103.325 ;
        RECT 58.825 103.255 59.615 103.505 ;
        RECT 58.055 102.765 58.405 102.935 ;
        RECT 59.820 102.965 59.990 103.675 ;
        RECT 60.345 103.475 60.515 104.065 ;
        RECT 60.160 103.255 60.515 103.475 ;
        RECT 60.685 103.255 61.035 103.875 ;
        RECT 61.205 102.965 61.375 104.325 ;
        RECT 61.740 104.155 62.065 104.940 ;
        RECT 61.545 103.105 62.005 104.155 ;
        RECT 59.820 102.795 60.675 102.965 ;
        RECT 60.880 102.795 61.375 102.965 ;
        RECT 62.235 102.835 62.405 104.955 ;
        RECT 63.075 104.455 63.330 104.955 ;
        RECT 62.580 104.285 63.330 104.455 ;
        RECT 62.580 103.295 62.810 104.285 ;
        RECT 62.980 103.465 63.330 104.115 ;
        RECT 63.510 103.935 63.765 104.815 ;
        RECT 65.090 104.575 65.260 104.865 ;
        RECT 64.460 104.405 65.260 104.575 ;
        RECT 65.850 104.615 66.720 104.955 ;
        RECT 62.580 103.125 63.330 103.295 ;
        RECT 63.075 102.835 63.330 103.125 ;
        RECT 63.510 103.285 63.720 103.935 ;
        RECT 64.460 103.815 64.630 104.405 ;
        RECT 65.850 104.235 66.020 104.615 ;
        RECT 66.955 104.495 67.125 104.955 ;
        RECT 67.960 104.525 68.130 104.865 ;
        RECT 68.865 104.525 69.035 104.865 ;
        RECT 64.800 104.065 66.020 104.235 ;
        RECT 66.190 104.155 66.650 104.445 ;
        RECT 66.955 104.325 67.515 104.495 ;
        RECT 67.960 104.355 69.035 104.525 ;
        RECT 69.205 104.625 69.885 104.955 ;
        RECT 70.100 104.625 70.350 104.955 ;
        RECT 67.345 104.185 67.515 104.325 ;
        RECT 66.190 104.145 67.155 104.155 ;
        RECT 65.850 103.975 66.020 104.065 ;
        RECT 66.480 103.985 67.155 104.145 ;
        RECT 63.890 103.785 64.630 103.815 ;
        RECT 63.890 103.485 64.805 103.785 ;
        RECT 64.480 103.310 64.805 103.485 ;
        RECT 63.510 102.755 63.765 103.285 ;
        RECT 64.485 102.955 64.805 103.310 ;
        RECT 64.975 103.525 65.515 103.895 ;
        RECT 65.850 103.805 66.255 103.975 ;
        RECT 64.975 103.125 65.215 103.525 ;
        RECT 65.695 103.355 65.915 103.635 ;
        RECT 65.385 103.185 65.915 103.355 ;
        RECT 65.385 102.955 65.555 103.185 ;
        RECT 64.485 102.785 65.555 102.955 ;
        RECT 66.085 103.025 66.255 103.805 ;
        RECT 66.425 103.195 66.775 103.815 ;
        RECT 66.945 103.195 67.155 103.985 ;
        RECT 67.345 104.015 68.845 104.185 ;
        RECT 67.345 103.325 67.515 104.015 ;
        RECT 69.205 103.845 69.375 104.625 ;
        RECT 70.180 104.495 70.350 104.625 ;
        RECT 67.685 103.675 69.375 103.845 ;
        RECT 69.545 104.065 70.010 104.455 ;
        RECT 70.180 104.325 70.575 104.495 ;
        RECT 67.685 103.495 67.855 103.675 ;
        RECT 66.085 102.745 67.035 103.025 ;
        RECT 67.345 102.935 67.605 103.325 ;
        RECT 68.025 103.255 68.815 103.505 ;
        RECT 67.255 102.765 67.605 102.935 ;
        RECT 69.020 102.965 69.190 103.675 ;
        RECT 69.545 103.475 69.715 104.065 ;
        RECT 69.360 103.255 69.715 103.475 ;
        RECT 69.885 103.255 70.235 103.875 ;
        RECT 70.405 102.965 70.575 104.325 ;
        RECT 70.940 104.155 71.265 104.940 ;
        RECT 70.745 103.105 71.205 104.155 ;
        RECT 69.020 102.795 69.875 102.965 ;
        RECT 70.080 102.795 70.575 102.965 ;
        RECT 71.435 102.835 71.605 104.955 ;
        RECT 72.275 104.455 72.530 104.955 ;
        RECT 71.780 104.285 72.530 104.455 ;
        RECT 71.780 103.295 72.010 104.285 ;
        RECT 72.180 103.465 72.530 104.115 ;
        RECT 76.390 103.935 76.645 104.815 ;
        RECT 77.970 104.575 78.140 104.865 ;
        RECT 77.340 104.405 78.140 104.575 ;
        RECT 78.730 104.615 79.600 104.955 ;
        RECT 71.780 103.125 72.530 103.295 ;
        RECT 72.275 102.835 72.530 103.125 ;
        RECT 76.390 103.285 76.600 103.935 ;
        RECT 77.340 103.815 77.510 104.405 ;
        RECT 78.730 104.235 78.900 104.615 ;
        RECT 79.835 104.495 80.005 104.955 ;
        RECT 80.840 104.525 81.010 104.865 ;
        RECT 81.745 104.525 81.915 104.865 ;
        RECT 77.680 104.065 78.900 104.235 ;
        RECT 79.070 104.155 79.530 104.445 ;
        RECT 79.835 104.325 80.395 104.495 ;
        RECT 80.840 104.355 81.915 104.525 ;
        RECT 82.085 104.625 82.765 104.955 ;
        RECT 82.980 104.625 83.230 104.955 ;
        RECT 80.225 104.185 80.395 104.325 ;
        RECT 79.070 104.145 80.035 104.155 ;
        RECT 78.730 103.975 78.900 104.065 ;
        RECT 79.360 103.985 80.035 104.145 ;
        RECT 76.770 103.785 77.510 103.815 ;
        RECT 76.770 103.485 77.685 103.785 ;
        RECT 77.360 103.310 77.685 103.485 ;
        RECT 76.390 102.755 76.645 103.285 ;
        RECT 77.365 102.955 77.685 103.310 ;
        RECT 77.855 103.525 78.395 103.895 ;
        RECT 78.730 103.805 79.135 103.975 ;
        RECT 77.855 103.125 78.095 103.525 ;
        RECT 78.575 103.355 78.795 103.635 ;
        RECT 78.265 103.185 78.795 103.355 ;
        RECT 78.265 102.955 78.435 103.185 ;
        RECT 77.365 102.785 78.435 102.955 ;
        RECT 78.965 103.025 79.135 103.805 ;
        RECT 79.305 103.195 79.655 103.815 ;
        RECT 79.825 103.195 80.035 103.985 ;
        RECT 80.225 104.015 81.725 104.185 ;
        RECT 80.225 103.325 80.395 104.015 ;
        RECT 82.085 103.845 82.255 104.625 ;
        RECT 83.060 104.495 83.230 104.625 ;
        RECT 80.565 103.675 82.255 103.845 ;
        RECT 82.425 104.065 82.890 104.455 ;
        RECT 83.060 104.325 83.455 104.495 ;
        RECT 80.565 103.495 80.735 103.675 ;
        RECT 78.965 102.745 79.915 103.025 ;
        RECT 80.225 102.935 80.485 103.325 ;
        RECT 80.905 103.255 81.695 103.505 ;
        RECT 80.135 102.765 80.485 102.935 ;
        RECT 81.900 102.965 82.070 103.675 ;
        RECT 82.425 103.475 82.595 104.065 ;
        RECT 82.240 103.255 82.595 103.475 ;
        RECT 82.765 103.255 83.115 103.875 ;
        RECT 83.285 102.965 83.455 104.325 ;
        RECT 83.820 104.155 84.145 104.940 ;
        RECT 83.625 103.105 84.085 104.155 ;
        RECT 81.900 102.795 82.755 102.965 ;
        RECT 82.960 102.795 83.455 102.965 ;
        RECT 84.315 102.835 84.485 104.955 ;
        RECT 85.155 104.455 85.410 104.955 ;
        RECT 84.660 104.285 85.410 104.455 ;
        RECT 84.660 103.295 84.890 104.285 ;
        RECT 85.060 103.465 85.410 104.115 ;
        RECT 85.590 103.935 85.845 104.815 ;
        RECT 87.170 104.575 87.340 104.865 ;
        RECT 86.540 104.405 87.340 104.575 ;
        RECT 87.930 104.615 88.800 104.955 ;
        RECT 84.660 103.125 85.410 103.295 ;
        RECT 85.155 102.835 85.410 103.125 ;
        RECT 85.590 103.285 85.800 103.935 ;
        RECT 86.540 103.815 86.710 104.405 ;
        RECT 87.930 104.235 88.100 104.615 ;
        RECT 89.035 104.495 89.205 104.955 ;
        RECT 90.040 104.525 90.210 104.865 ;
        RECT 90.945 104.525 91.115 104.865 ;
        RECT 86.880 104.065 88.100 104.235 ;
        RECT 88.270 104.155 88.730 104.445 ;
        RECT 89.035 104.325 89.595 104.495 ;
        RECT 90.040 104.355 91.115 104.525 ;
        RECT 91.285 104.625 91.965 104.955 ;
        RECT 92.180 104.625 92.430 104.955 ;
        RECT 89.425 104.185 89.595 104.325 ;
        RECT 88.270 104.145 89.235 104.155 ;
        RECT 87.930 103.975 88.100 104.065 ;
        RECT 88.560 103.985 89.235 104.145 ;
        RECT 85.970 103.785 86.710 103.815 ;
        RECT 85.970 103.485 86.885 103.785 ;
        RECT 86.560 103.310 86.885 103.485 ;
        RECT 85.590 102.755 85.845 103.285 ;
        RECT 86.565 102.955 86.885 103.310 ;
        RECT 87.055 103.525 87.595 103.895 ;
        RECT 87.930 103.805 88.335 103.975 ;
        RECT 87.055 103.125 87.295 103.525 ;
        RECT 87.775 103.355 87.995 103.635 ;
        RECT 87.465 103.185 87.995 103.355 ;
        RECT 87.465 102.955 87.635 103.185 ;
        RECT 86.565 102.785 87.635 102.955 ;
        RECT 88.165 103.025 88.335 103.805 ;
        RECT 88.505 103.195 88.855 103.815 ;
        RECT 89.025 103.195 89.235 103.985 ;
        RECT 89.425 104.015 90.925 104.185 ;
        RECT 89.425 103.325 89.595 104.015 ;
        RECT 91.285 103.845 91.455 104.625 ;
        RECT 92.260 104.495 92.430 104.625 ;
        RECT 89.765 103.675 91.455 103.845 ;
        RECT 91.625 104.065 92.090 104.455 ;
        RECT 92.260 104.325 92.655 104.495 ;
        RECT 89.765 103.495 89.935 103.675 ;
        RECT 88.165 102.745 89.115 103.025 ;
        RECT 89.425 102.935 89.685 103.325 ;
        RECT 90.105 103.255 90.895 103.505 ;
        RECT 89.335 102.765 89.685 102.935 ;
        RECT 91.100 102.965 91.270 103.675 ;
        RECT 91.625 103.475 91.795 104.065 ;
        RECT 91.440 103.255 91.795 103.475 ;
        RECT 91.965 103.255 92.315 103.875 ;
        RECT 92.485 102.965 92.655 104.325 ;
        RECT 93.020 104.155 93.345 104.940 ;
        RECT 92.825 103.105 93.285 104.155 ;
        RECT 91.100 102.795 91.955 102.965 ;
        RECT 92.160 102.795 92.655 102.965 ;
        RECT 93.515 102.835 93.685 104.955 ;
        RECT 94.355 104.455 94.610 104.955 ;
        RECT 93.860 104.285 94.610 104.455 ;
        RECT 93.860 103.295 94.090 104.285 ;
        RECT 94.875 104.195 95.045 104.955 ;
        RECT 94.260 103.465 94.610 104.115 ;
        RECT 94.875 104.025 95.540 104.195 ;
        RECT 95.725 104.050 95.995 104.955 ;
        RECT 102.150 104.455 102.405 104.955 ;
        RECT 102.150 104.285 102.900 104.455 ;
        RECT 95.370 103.880 95.540 104.025 ;
        RECT 94.805 103.475 95.135 103.845 ;
        RECT 95.370 103.550 95.655 103.880 ;
        RECT 95.370 103.295 95.540 103.550 ;
        RECT 93.860 103.125 94.610 103.295 ;
        RECT 94.355 102.835 94.610 103.125 ;
        RECT 94.875 103.125 95.540 103.295 ;
        RECT 95.825 103.250 95.995 104.050 ;
        RECT 102.150 103.465 102.500 104.115 ;
        RECT 102.670 103.295 102.900 104.285 ;
        RECT 94.875 102.745 95.045 103.125 ;
        RECT 95.735 102.745 95.995 103.250 ;
        RECT 102.150 103.125 102.900 103.295 ;
        RECT 102.150 102.835 102.405 103.125 ;
        RECT 103.075 102.835 103.245 104.955 ;
        RECT 103.415 104.155 103.740 104.940 ;
        RECT 104.330 104.625 104.580 104.955 ;
        RECT 104.795 104.625 105.475 104.955 ;
        RECT 104.330 104.495 104.500 104.625 ;
        RECT 104.105 104.325 104.500 104.495 ;
        RECT 103.475 103.105 103.935 104.155 ;
        RECT 104.105 102.965 104.275 104.325 ;
        RECT 104.670 104.065 105.135 104.455 ;
        RECT 104.445 103.255 104.795 103.875 ;
        RECT 104.965 103.475 105.135 104.065 ;
        RECT 105.305 103.845 105.475 104.625 ;
        RECT 105.645 104.525 105.815 104.865 ;
        RECT 106.550 104.525 106.720 104.865 ;
        RECT 105.645 104.355 106.720 104.525 ;
        RECT 107.555 104.495 107.725 104.955 ;
        RECT 107.960 104.615 108.830 104.955 ;
        RECT 107.165 104.325 107.725 104.495 ;
        RECT 107.165 104.185 107.335 104.325 ;
        RECT 105.835 104.015 107.335 104.185 ;
        RECT 108.030 104.155 108.490 104.445 ;
        RECT 105.305 103.675 106.995 103.845 ;
        RECT 104.965 103.255 105.320 103.475 ;
        RECT 105.490 102.965 105.660 103.675 ;
        RECT 105.865 103.255 106.655 103.505 ;
        RECT 106.825 103.495 106.995 103.675 ;
        RECT 107.165 103.325 107.335 104.015 ;
        RECT 104.105 102.795 104.600 102.965 ;
        RECT 104.805 102.795 105.660 102.965 ;
        RECT 107.075 102.935 107.335 103.325 ;
        RECT 107.525 104.145 108.490 104.155 ;
        RECT 108.660 104.235 108.830 104.615 ;
        RECT 109.420 104.575 109.590 104.865 ;
        RECT 109.420 104.405 110.220 104.575 ;
        RECT 107.525 103.985 108.200 104.145 ;
        RECT 108.660 104.065 109.880 104.235 ;
        RECT 107.525 103.195 107.735 103.985 ;
        RECT 108.660 103.975 108.830 104.065 ;
        RECT 107.905 103.195 108.255 103.815 ;
        RECT 108.425 103.805 108.830 103.975 ;
        RECT 108.425 103.025 108.595 103.805 ;
        RECT 108.765 103.355 108.985 103.635 ;
        RECT 109.165 103.525 109.705 103.895 ;
        RECT 110.050 103.815 110.220 104.405 ;
        RECT 110.915 103.935 111.170 104.815 ;
        RECT 110.050 103.785 110.790 103.815 ;
        RECT 108.765 103.185 109.295 103.355 ;
        RECT 107.075 102.765 107.425 102.935 ;
        RECT 107.645 102.745 108.595 103.025 ;
        RECT 109.125 102.955 109.295 103.185 ;
        RECT 109.465 103.125 109.705 103.525 ;
        RECT 109.875 103.485 110.790 103.785 ;
        RECT 109.875 103.310 110.200 103.485 ;
        RECT 109.875 102.955 110.195 103.310 ;
        RECT 110.960 103.285 111.170 103.935 ;
        RECT 109.125 102.785 110.195 102.955 ;
        RECT 110.915 102.755 111.170 103.285 ;
        RECT 111.350 103.935 111.605 104.815 ;
        RECT 112.930 104.575 113.100 104.865 ;
        RECT 112.300 104.405 113.100 104.575 ;
        RECT 113.690 104.615 114.560 104.955 ;
        RECT 111.350 103.285 111.560 103.935 ;
        RECT 112.300 103.815 112.470 104.405 ;
        RECT 113.690 104.235 113.860 104.615 ;
        RECT 114.795 104.495 114.965 104.955 ;
        RECT 115.800 104.525 115.970 104.865 ;
        RECT 116.705 104.525 116.875 104.865 ;
        RECT 112.640 104.065 113.860 104.235 ;
        RECT 114.030 104.155 114.490 104.445 ;
        RECT 114.795 104.325 115.355 104.495 ;
        RECT 115.800 104.355 116.875 104.525 ;
        RECT 117.045 104.625 117.725 104.955 ;
        RECT 117.940 104.625 118.190 104.955 ;
        RECT 115.185 104.185 115.355 104.325 ;
        RECT 114.030 104.145 114.995 104.155 ;
        RECT 113.690 103.975 113.860 104.065 ;
        RECT 114.320 103.985 114.995 104.145 ;
        RECT 111.730 103.785 112.470 103.815 ;
        RECT 111.730 103.485 112.645 103.785 ;
        RECT 112.320 103.310 112.645 103.485 ;
        RECT 111.350 102.755 111.605 103.285 ;
        RECT 112.325 102.955 112.645 103.310 ;
        RECT 112.815 103.525 113.355 103.895 ;
        RECT 113.690 103.805 114.095 103.975 ;
        RECT 112.815 103.125 113.055 103.525 ;
        RECT 113.535 103.355 113.755 103.635 ;
        RECT 113.225 103.185 113.755 103.355 ;
        RECT 113.225 102.955 113.395 103.185 ;
        RECT 112.325 102.785 113.395 102.955 ;
        RECT 113.925 103.025 114.095 103.805 ;
        RECT 114.265 103.195 114.615 103.815 ;
        RECT 114.785 103.195 114.995 103.985 ;
        RECT 115.185 104.015 116.685 104.185 ;
        RECT 115.185 103.325 115.355 104.015 ;
        RECT 117.045 103.845 117.215 104.625 ;
        RECT 118.020 104.495 118.190 104.625 ;
        RECT 115.525 103.675 117.215 103.845 ;
        RECT 117.385 104.065 117.850 104.455 ;
        RECT 118.020 104.325 118.415 104.495 ;
        RECT 115.525 103.495 115.695 103.675 ;
        RECT 113.925 102.745 114.875 103.025 ;
        RECT 115.185 102.935 115.445 103.325 ;
        RECT 115.865 103.255 116.655 103.505 ;
        RECT 115.095 102.765 115.445 102.935 ;
        RECT 116.860 102.965 117.030 103.675 ;
        RECT 117.385 103.475 117.555 104.065 ;
        RECT 117.200 103.255 117.555 103.475 ;
        RECT 117.725 103.255 118.075 103.875 ;
        RECT 118.245 102.965 118.415 104.325 ;
        RECT 118.780 104.155 119.105 104.940 ;
        RECT 118.585 103.105 119.045 104.155 ;
        RECT 116.860 102.795 117.715 102.965 ;
        RECT 117.920 102.795 118.415 102.965 ;
        RECT 119.275 102.835 119.445 104.955 ;
        RECT 120.115 104.455 120.370 104.955 ;
        RECT 119.620 104.285 120.370 104.455 ;
        RECT 119.620 103.295 119.850 104.285 ;
        RECT 120.020 103.465 120.370 104.115 ;
        RECT 125.145 104.050 125.415 104.955 ;
        RECT 126.095 104.195 126.275 104.955 ;
        RECT 119.620 103.125 120.370 103.295 ;
        RECT 120.115 102.835 120.370 103.125 ;
        RECT 125.145 103.250 125.325 104.050 ;
        RECT 125.600 104.025 126.275 104.195 ;
        RECT 125.600 103.880 125.770 104.025 ;
        RECT 125.495 103.550 125.770 103.880 ;
        RECT 125.600 103.295 125.770 103.550 ;
        RECT 125.145 102.745 125.405 103.250 ;
        RECT 125.600 103.125 126.265 103.295 ;
        RECT 126.095 102.745 126.265 103.125 ;
        RECT 28.645 101.755 28.905 102.210 ;
        RECT 29.515 101.755 29.775 102.210 ;
        RECT 30.375 101.755 30.635 102.210 ;
        RECT 31.235 101.755 31.495 102.210 ;
        RECT 32.080 101.755 32.355 102.210 ;
        RECT 32.940 101.755 33.200 102.210 ;
        RECT 33.800 101.755 34.060 102.210 ;
        RECT 34.660 101.755 34.920 102.210 ;
        RECT 28.175 101.585 34.920 101.755 ;
        RECT 28.175 100.995 29.340 101.585 ;
        RECT 35.520 101.415 35.770 102.225 ;
        RECT 36.380 101.415 36.630 102.225 ;
        RECT 29.510 101.165 36.630 101.415 ;
        RECT 36.800 101.165 37.115 101.725 ;
        RECT 38.645 101.605 38.975 102.235 ;
        RECT 39.585 101.730 39.845 102.235 ;
        RECT 40.535 101.855 40.705 102.235 ;
        RECT 28.175 100.770 34.920 100.995 ;
        RECT 28.615 100.030 28.905 100.770 ;
        RECT 29.515 100.755 34.920 100.770 ;
        RECT 29.515 100.030 29.775 100.755 ;
        RECT 30.375 100.030 30.635 100.755 ;
        RECT 31.235 100.030 31.495 100.755 ;
        RECT 32.080 100.030 32.340 100.755 ;
        RECT 32.940 100.030 33.200 100.755 ;
        RECT 33.800 100.030 34.060 100.755 ;
        RECT 34.660 100.030 34.920 100.755 ;
        RECT 35.520 100.030 35.770 101.165 ;
        RECT 36.385 100.025 36.630 101.165 ;
        RECT 38.645 101.005 38.895 101.605 ;
        RECT 39.065 101.165 39.395 101.415 ;
        RECT 38.645 100.025 38.975 101.005 ;
        RECT 39.585 100.930 39.755 101.730 ;
        RECT 40.040 101.685 40.705 101.855 ;
        RECT 41.525 101.755 41.785 102.210 ;
        RECT 42.395 101.755 42.655 102.210 ;
        RECT 43.255 101.755 43.515 102.210 ;
        RECT 44.115 101.755 44.375 102.210 ;
        RECT 44.960 101.755 45.235 102.210 ;
        RECT 45.820 101.755 46.080 102.210 ;
        RECT 46.680 101.755 46.940 102.210 ;
        RECT 47.540 101.755 47.800 102.210 ;
        RECT 40.040 101.430 40.210 101.685 ;
        RECT 41.055 101.585 47.800 101.755 ;
        RECT 39.925 101.100 40.210 101.430 ;
        RECT 40.445 101.135 40.775 101.505 ;
        RECT 40.040 100.955 40.210 101.100 ;
        RECT 41.055 100.995 42.220 101.585 ;
        RECT 48.400 101.415 48.650 102.225 ;
        RECT 49.260 101.415 49.510 102.225 ;
        RECT 53.485 101.755 53.745 102.210 ;
        RECT 54.355 101.755 54.615 102.210 ;
        RECT 55.215 101.755 55.475 102.210 ;
        RECT 56.075 101.755 56.335 102.210 ;
        RECT 56.920 101.755 57.195 102.210 ;
        RECT 57.780 101.755 58.040 102.210 ;
        RECT 58.640 101.755 58.900 102.210 ;
        RECT 59.500 101.755 59.760 102.210 ;
        RECT 42.390 101.165 49.510 101.415 ;
        RECT 49.680 101.165 49.995 101.725 ;
        RECT 53.015 101.585 59.760 101.755 ;
        RECT 39.585 100.025 39.855 100.930 ;
        RECT 40.040 100.785 40.705 100.955 ;
        RECT 40.535 100.025 40.705 100.785 ;
        RECT 41.055 100.770 47.800 100.995 ;
        RECT 41.495 100.030 41.785 100.770 ;
        RECT 42.395 100.755 47.800 100.770 ;
        RECT 42.395 100.030 42.655 100.755 ;
        RECT 43.255 100.030 43.515 100.755 ;
        RECT 44.115 100.030 44.375 100.755 ;
        RECT 44.960 100.030 45.220 100.755 ;
        RECT 45.820 100.030 46.080 100.755 ;
        RECT 46.680 100.030 46.940 100.755 ;
        RECT 47.540 100.030 47.800 100.755 ;
        RECT 48.400 100.030 48.650 101.165 ;
        RECT 49.265 100.025 49.510 101.165 ;
        RECT 53.015 100.995 54.180 101.585 ;
        RECT 60.360 101.415 60.610 102.225 ;
        RECT 61.220 101.415 61.470 102.225 ;
        RECT 54.350 101.165 61.470 101.415 ;
        RECT 61.640 101.165 61.955 101.725 ;
        RECT 63.505 101.165 63.820 101.725 ;
        RECT 63.990 101.415 64.240 102.225 ;
        RECT 64.850 101.415 65.100 102.225 ;
        RECT 65.700 101.755 65.960 102.210 ;
        RECT 66.560 101.755 66.820 102.210 ;
        RECT 67.420 101.755 67.680 102.210 ;
        RECT 68.265 101.755 68.540 102.210 ;
        RECT 69.125 101.755 69.385 102.210 ;
        RECT 69.985 101.755 70.245 102.210 ;
        RECT 70.845 101.755 71.105 102.210 ;
        RECT 71.715 101.755 71.975 102.210 ;
        RECT 65.700 101.585 72.445 101.755 ;
        RECT 63.990 101.165 71.110 101.415 ;
        RECT 53.015 100.770 59.760 100.995 ;
        RECT 53.455 100.030 53.745 100.770 ;
        RECT 54.355 100.755 59.760 100.770 ;
        RECT 54.355 100.030 54.615 100.755 ;
        RECT 55.215 100.030 55.475 100.755 ;
        RECT 56.075 100.030 56.335 100.755 ;
        RECT 56.920 100.030 57.180 100.755 ;
        RECT 57.780 100.030 58.040 100.755 ;
        RECT 58.640 100.030 58.900 100.755 ;
        RECT 59.500 100.030 59.760 100.755 ;
        RECT 60.360 100.030 60.610 101.165 ;
        RECT 61.225 100.025 61.470 101.165 ;
        RECT 63.990 100.025 64.235 101.165 ;
        RECT 64.850 100.030 65.100 101.165 ;
        RECT 71.280 100.995 72.445 101.585 ;
        RECT 76.385 101.165 76.700 101.725 ;
        RECT 76.870 101.415 77.120 102.225 ;
        RECT 77.730 101.415 77.980 102.225 ;
        RECT 78.580 101.755 78.840 102.210 ;
        RECT 79.440 101.755 79.700 102.210 ;
        RECT 80.300 101.755 80.560 102.210 ;
        RECT 81.145 101.755 81.420 102.210 ;
        RECT 82.005 101.755 82.265 102.210 ;
        RECT 82.865 101.755 83.125 102.210 ;
        RECT 83.725 101.755 83.985 102.210 ;
        RECT 84.595 101.755 84.855 102.210 ;
        RECT 78.580 101.585 85.325 101.755 ;
        RECT 76.870 101.165 83.990 101.415 ;
        RECT 65.700 100.770 72.445 100.995 ;
        RECT 65.700 100.755 71.105 100.770 ;
        RECT 65.700 100.030 65.960 100.755 ;
        RECT 66.560 100.030 66.820 100.755 ;
        RECT 67.420 100.030 67.680 100.755 ;
        RECT 68.280 100.030 68.540 100.755 ;
        RECT 69.125 100.030 69.385 100.755 ;
        RECT 69.985 100.030 70.245 100.755 ;
        RECT 70.845 100.030 71.105 100.755 ;
        RECT 71.715 100.030 72.005 100.770 ;
        RECT 76.870 100.025 77.115 101.165 ;
        RECT 77.730 100.030 77.980 101.165 ;
        RECT 84.160 100.995 85.325 101.585 ;
        RECT 89.265 101.165 89.580 101.725 ;
        RECT 89.750 101.415 90.000 102.225 ;
        RECT 90.610 101.415 90.860 102.225 ;
        RECT 91.460 101.755 91.720 102.210 ;
        RECT 92.320 101.755 92.580 102.210 ;
        RECT 93.180 101.755 93.440 102.210 ;
        RECT 94.025 101.755 94.300 102.210 ;
        RECT 94.885 101.755 95.145 102.210 ;
        RECT 95.745 101.755 96.005 102.210 ;
        RECT 96.605 101.755 96.865 102.210 ;
        RECT 97.475 101.755 97.735 102.210 ;
        RECT 102.705 101.755 102.965 102.210 ;
        RECT 103.575 101.755 103.835 102.210 ;
        RECT 104.435 101.755 104.695 102.210 ;
        RECT 105.295 101.755 105.555 102.210 ;
        RECT 106.140 101.755 106.415 102.210 ;
        RECT 107.000 101.755 107.260 102.210 ;
        RECT 107.860 101.755 108.120 102.210 ;
        RECT 108.720 101.755 108.980 102.210 ;
        RECT 91.460 101.585 98.205 101.755 ;
        RECT 89.750 101.165 96.870 101.415 ;
        RECT 78.580 100.770 85.325 100.995 ;
        RECT 78.580 100.755 83.985 100.770 ;
        RECT 78.580 100.030 78.840 100.755 ;
        RECT 79.440 100.030 79.700 100.755 ;
        RECT 80.300 100.030 80.560 100.755 ;
        RECT 81.160 100.030 81.420 100.755 ;
        RECT 82.005 100.030 82.265 100.755 ;
        RECT 82.865 100.030 83.125 100.755 ;
        RECT 83.725 100.030 83.985 100.755 ;
        RECT 84.595 100.030 84.885 100.770 ;
        RECT 89.750 100.025 89.995 101.165 ;
        RECT 90.610 100.030 90.860 101.165 ;
        RECT 97.040 100.995 98.205 101.585 ;
        RECT 91.460 100.770 98.205 100.995 ;
        RECT 102.235 101.585 108.980 101.755 ;
        RECT 102.235 100.995 103.400 101.585 ;
        RECT 109.580 101.415 109.830 102.225 ;
        RECT 110.440 101.415 110.690 102.225 ;
        RECT 103.570 101.165 110.690 101.415 ;
        RECT 110.860 101.165 111.175 101.725 ;
        RECT 115.025 101.165 115.340 101.725 ;
        RECT 115.510 101.415 115.760 102.225 ;
        RECT 116.370 101.415 116.620 102.225 ;
        RECT 117.220 101.755 117.480 102.210 ;
        RECT 118.080 101.755 118.340 102.210 ;
        RECT 118.940 101.755 119.200 102.210 ;
        RECT 119.785 101.755 120.060 102.210 ;
        RECT 120.645 101.755 120.905 102.210 ;
        RECT 121.505 101.755 121.765 102.210 ;
        RECT 122.365 101.755 122.625 102.210 ;
        RECT 123.235 101.755 123.495 102.210 ;
        RECT 117.220 101.585 123.965 101.755 ;
        RECT 115.510 101.165 122.630 101.415 ;
        RECT 102.235 100.770 108.980 100.995 ;
        RECT 91.460 100.755 96.865 100.770 ;
        RECT 91.460 100.030 91.720 100.755 ;
        RECT 92.320 100.030 92.580 100.755 ;
        RECT 93.180 100.030 93.440 100.755 ;
        RECT 94.040 100.030 94.300 100.755 ;
        RECT 94.885 100.030 95.145 100.755 ;
        RECT 95.745 100.030 96.005 100.755 ;
        RECT 96.605 100.030 96.865 100.755 ;
        RECT 97.475 100.030 97.765 100.770 ;
        RECT 102.675 100.030 102.965 100.770 ;
        RECT 103.575 100.755 108.980 100.770 ;
        RECT 103.575 100.030 103.835 100.755 ;
        RECT 104.435 100.030 104.695 100.755 ;
        RECT 105.295 100.030 105.555 100.755 ;
        RECT 106.140 100.030 106.400 100.755 ;
        RECT 107.000 100.030 107.260 100.755 ;
        RECT 107.860 100.030 108.120 100.755 ;
        RECT 108.720 100.030 108.980 100.755 ;
        RECT 109.580 100.030 109.830 101.165 ;
        RECT 110.445 100.025 110.690 101.165 ;
        RECT 115.510 100.025 115.755 101.165 ;
        RECT 116.370 100.030 116.620 101.165 ;
        RECT 122.800 100.995 123.965 101.585 ;
        RECT 117.220 100.770 123.965 100.995 ;
        RECT 117.220 100.755 122.625 100.770 ;
        RECT 117.220 100.030 117.480 100.755 ;
        RECT 118.080 100.030 118.340 100.755 ;
        RECT 118.940 100.030 119.200 100.755 ;
        RECT 119.800 100.030 120.060 100.755 ;
        RECT 120.645 100.030 120.905 100.755 ;
        RECT 121.505 100.030 121.765 100.755 ;
        RECT 122.365 100.030 122.625 100.755 ;
        RECT 123.235 100.030 123.525 100.770 ;
        RECT 26.525 55.300 26.695 65.340 ;
        RECT 27.665 55.300 27.835 65.340 ;
        RECT 28.955 55.300 29.125 65.340 ;
        RECT 37.725 55.310 37.895 65.350 ;
        RECT 38.865 55.310 39.035 65.350 ;
        RECT 40.155 55.310 40.325 65.350 ;
        RECT 48.945 55.280 49.115 65.320 ;
        RECT 50.085 55.280 50.255 65.320 ;
        RECT 51.375 55.280 51.545 65.320 ;
        RECT 60.195 55.260 60.365 65.300 ;
        RECT 61.335 55.260 61.505 65.300 ;
        RECT 62.625 55.260 62.795 65.300 ;
        RECT 71.415 55.250 71.585 65.290 ;
        RECT 72.555 55.250 72.725 65.290 ;
        RECT 73.845 55.250 74.015 65.290 ;
        RECT 82.655 55.240 82.825 65.280 ;
        RECT 83.795 55.240 83.965 65.280 ;
        RECT 85.085 55.240 85.255 65.280 ;
        RECT 93.905 55.250 94.075 65.290 ;
        RECT 95.045 55.250 95.215 65.290 ;
        RECT 96.335 55.250 96.505 65.290 ;
        RECT 105.185 55.240 105.355 65.280 ;
        RECT 106.325 55.240 106.495 65.280 ;
        RECT 107.615 55.240 107.785 65.280 ;
        RECT 116.455 55.240 116.625 65.280 ;
        RECT 117.595 55.240 117.765 65.280 ;
        RECT 118.885 55.240 119.055 65.280 ;
        RECT 127.705 55.240 127.875 65.280 ;
        RECT 128.845 55.240 129.015 65.280 ;
        RECT 130.135 55.240 130.305 65.280 ;
        RECT 21.635 52.350 22.135 52.520 ;
        RECT 25.715 52.270 26.215 52.440 ;
        RECT 27.645 52.270 28.145 52.440 ;
        RECT 32.835 52.360 33.335 52.530 ;
        RECT 36.915 52.280 37.415 52.450 ;
        RECT 38.845 52.280 39.345 52.450 ;
        RECT 44.055 52.330 44.555 52.500 ;
        RECT 48.135 52.250 48.635 52.420 ;
        RECT 50.065 52.250 50.565 52.420 ;
        RECT 55.305 52.310 55.805 52.480 ;
        RECT 59.385 52.230 59.885 52.400 ;
        RECT 61.315 52.230 61.815 52.400 ;
        RECT 66.525 52.300 67.025 52.470 ;
        RECT 70.605 52.220 71.105 52.390 ;
        RECT 72.535 52.220 73.035 52.390 ;
        RECT 77.765 52.290 78.265 52.460 ;
        RECT 81.845 52.210 82.345 52.380 ;
        RECT 83.775 52.210 84.275 52.380 ;
        RECT 89.015 52.300 89.515 52.470 ;
        RECT 93.095 52.220 93.595 52.390 ;
        RECT 95.025 52.220 95.525 52.390 ;
        RECT 100.295 52.290 100.795 52.460 ;
        RECT 104.375 52.210 104.875 52.380 ;
        RECT 106.305 52.210 106.805 52.380 ;
        RECT 111.565 52.290 112.065 52.460 ;
        RECT 115.645 52.210 116.145 52.380 ;
        RECT 117.575 52.210 118.075 52.380 ;
        RECT 122.815 52.290 123.315 52.460 ;
        RECT 126.895 52.210 127.395 52.380 ;
        RECT 128.825 52.210 129.325 52.380 ;
        RECT 22.195 50.095 22.365 52.135 ;
        RECT 21.635 49.710 22.135 49.880 ;
        RECT 21.485 47.530 21.985 47.700 ;
        RECT 22.045 46.320 22.215 47.360 ;
        RECT 26.275 47.015 26.445 52.055 ;
        RECT 27.415 47.015 27.585 52.055 ;
        RECT 33.395 50.105 33.565 52.145 ;
        RECT 32.835 49.720 33.335 49.890 ;
        RECT 32.685 47.540 33.185 47.710 ;
        RECT 25.715 46.630 26.215 46.800 ;
        RECT 27.645 46.630 28.145 46.800 ;
        RECT 33.245 46.330 33.415 47.370 ;
        RECT 37.475 47.025 37.645 52.065 ;
        RECT 38.615 47.025 38.785 52.065 ;
        RECT 44.615 50.075 44.785 52.115 ;
        RECT 44.055 49.690 44.555 49.860 ;
        RECT 43.905 47.510 44.405 47.680 ;
        RECT 36.915 46.640 37.415 46.810 ;
        RECT 38.845 46.640 39.345 46.810 ;
        RECT 44.465 46.300 44.635 47.340 ;
        RECT 48.695 46.995 48.865 52.035 ;
        RECT 49.835 46.995 50.005 52.035 ;
        RECT 55.865 50.055 56.035 52.095 ;
        RECT 55.305 49.670 55.805 49.840 ;
        RECT 55.155 47.490 55.655 47.660 ;
        RECT 48.135 46.610 48.635 46.780 ;
        RECT 50.065 46.610 50.565 46.780 ;
        RECT 55.715 46.280 55.885 47.320 ;
        RECT 59.945 46.975 60.115 52.015 ;
        RECT 61.085 46.975 61.255 52.015 ;
        RECT 67.085 50.045 67.255 52.085 ;
        RECT 66.525 49.660 67.025 49.830 ;
        RECT 66.375 47.480 66.875 47.650 ;
        RECT 59.385 46.590 59.885 46.760 ;
        RECT 61.315 46.590 61.815 46.760 ;
        RECT 66.935 46.270 67.105 47.310 ;
        RECT 71.165 46.965 71.335 52.005 ;
        RECT 72.305 46.965 72.475 52.005 ;
        RECT 78.325 50.035 78.495 52.075 ;
        RECT 77.765 49.650 78.265 49.820 ;
        RECT 77.615 47.470 78.115 47.640 ;
        RECT 70.605 46.580 71.105 46.750 ;
        RECT 72.535 46.580 73.035 46.750 ;
        RECT 78.175 46.260 78.345 47.300 ;
        RECT 82.405 46.955 82.575 51.995 ;
        RECT 83.545 46.955 83.715 51.995 ;
        RECT 89.575 50.045 89.745 52.085 ;
        RECT 89.015 49.660 89.515 49.830 ;
        RECT 88.865 47.480 89.365 47.650 ;
        RECT 81.845 46.570 82.345 46.740 ;
        RECT 83.775 46.570 84.275 46.740 ;
        RECT 89.425 46.270 89.595 47.310 ;
        RECT 93.655 46.965 93.825 52.005 ;
        RECT 94.795 46.965 94.965 52.005 ;
        RECT 100.855 50.035 101.025 52.075 ;
        RECT 100.295 49.650 100.795 49.820 ;
        RECT 100.145 47.470 100.645 47.640 ;
        RECT 93.095 46.580 93.595 46.750 ;
        RECT 95.025 46.580 95.525 46.750 ;
        RECT 100.705 46.260 100.875 47.300 ;
        RECT 104.935 46.955 105.105 51.995 ;
        RECT 106.075 46.955 106.245 51.995 ;
        RECT 112.125 50.035 112.295 52.075 ;
        RECT 111.565 49.650 112.065 49.820 ;
        RECT 111.415 47.470 111.915 47.640 ;
        RECT 104.375 46.570 104.875 46.740 ;
        RECT 106.305 46.570 106.805 46.740 ;
        RECT 111.975 46.260 112.145 47.300 ;
        RECT 116.205 46.955 116.375 51.995 ;
        RECT 117.345 46.955 117.515 51.995 ;
        RECT 123.375 50.035 123.545 52.075 ;
        RECT 122.815 49.650 123.315 49.820 ;
        RECT 122.665 47.470 123.165 47.640 ;
        RECT 115.645 46.570 116.145 46.740 ;
        RECT 117.575 46.570 118.075 46.740 ;
        RECT 123.225 46.260 123.395 47.300 ;
        RECT 127.455 46.955 127.625 51.995 ;
        RECT 128.595 46.955 128.765 51.995 ;
        RECT 126.895 46.570 127.395 46.740 ;
        RECT 128.825 46.570 129.325 46.740 ;
        RECT 21.485 45.980 21.985 46.150 ;
        RECT 32.685 45.990 33.185 46.160 ;
        RECT 43.905 45.960 44.405 46.130 ;
        RECT 55.155 45.940 55.655 46.110 ;
        RECT 66.375 45.930 66.875 46.100 ;
        RECT 77.615 45.920 78.115 46.090 ;
        RECT 88.865 45.930 89.365 46.100 ;
        RECT 100.145 45.920 100.645 46.090 ;
        RECT 111.415 45.920 111.915 46.090 ;
        RECT 122.665 45.920 123.165 46.090 ;
        RECT 26.755 39.260 27.255 39.430 ;
        RECT 38.035 39.260 38.535 39.430 ;
        RECT 49.325 39.240 49.825 39.410 ;
        RECT 60.545 39.240 61.045 39.410 ;
        RECT 71.745 39.240 72.245 39.410 ;
        RECT 83.035 39.230 83.535 39.400 ;
        RECT 94.275 39.250 94.775 39.420 ;
        RECT 105.485 39.270 105.985 39.440 ;
        RECT 116.685 39.310 117.185 39.480 ;
        RECT 127.895 39.330 128.395 39.500 ;
        RECT 20.595 38.610 21.095 38.780 ;
        RECT 22.525 38.610 23.025 38.780 ;
        RECT 21.155 33.355 21.325 38.395 ;
        RECT 22.295 33.355 22.465 38.395 ;
        RECT 26.525 38.050 26.695 39.090 ;
        RECT 31.875 38.610 32.375 38.780 ;
        RECT 33.805 38.610 34.305 38.780 ;
        RECT 26.755 37.710 27.255 37.880 ;
        RECT 26.605 35.530 27.105 35.700 ;
        RECT 26.375 33.275 26.545 35.315 ;
        RECT 32.435 33.355 32.605 38.395 ;
        RECT 33.575 33.355 33.745 38.395 ;
        RECT 37.805 38.050 37.975 39.090 ;
        RECT 43.165 38.590 43.665 38.760 ;
        RECT 45.095 38.590 45.595 38.760 ;
        RECT 38.035 37.710 38.535 37.880 ;
        RECT 37.885 35.530 38.385 35.700 ;
        RECT 37.655 33.275 37.825 35.315 ;
        RECT 43.725 33.335 43.895 38.375 ;
        RECT 44.865 33.335 45.035 38.375 ;
        RECT 49.095 38.030 49.265 39.070 ;
        RECT 54.385 38.590 54.885 38.760 ;
        RECT 56.315 38.590 56.815 38.760 ;
        RECT 49.325 37.690 49.825 37.860 ;
        RECT 49.175 35.510 49.675 35.680 ;
        RECT 48.945 33.255 49.115 35.295 ;
        RECT 54.945 33.335 55.115 38.375 ;
        RECT 56.085 33.335 56.255 38.375 ;
        RECT 60.315 38.030 60.485 39.070 ;
        RECT 65.585 38.590 66.085 38.760 ;
        RECT 67.515 38.590 68.015 38.760 ;
        RECT 60.545 37.690 61.045 37.860 ;
        RECT 60.395 35.510 60.895 35.680 ;
        RECT 60.165 33.255 60.335 35.295 ;
        RECT 66.145 33.335 66.315 38.375 ;
        RECT 67.285 33.335 67.455 38.375 ;
        RECT 71.515 38.030 71.685 39.070 ;
        RECT 76.875 38.580 77.375 38.750 ;
        RECT 78.805 38.580 79.305 38.750 ;
        RECT 71.745 37.690 72.245 37.860 ;
        RECT 71.595 35.510 72.095 35.680 ;
        RECT 71.365 33.255 71.535 35.295 ;
        RECT 77.435 33.325 77.605 38.365 ;
        RECT 78.575 33.325 78.745 38.365 ;
        RECT 82.805 38.020 82.975 39.060 ;
        RECT 88.115 38.600 88.615 38.770 ;
        RECT 90.045 38.600 90.545 38.770 ;
        RECT 83.035 37.680 83.535 37.850 ;
        RECT 82.885 35.500 83.385 35.670 ;
        RECT 82.655 33.245 82.825 35.285 ;
        RECT 88.675 33.345 88.845 38.385 ;
        RECT 89.815 33.345 89.985 38.385 ;
        RECT 94.045 38.040 94.215 39.080 ;
        RECT 99.325 38.620 99.825 38.790 ;
        RECT 101.255 38.620 101.755 38.790 ;
        RECT 94.275 37.700 94.775 37.870 ;
        RECT 94.125 35.520 94.625 35.690 ;
        RECT 93.895 33.265 94.065 35.305 ;
        RECT 99.885 33.365 100.055 38.405 ;
        RECT 101.025 33.365 101.195 38.405 ;
        RECT 105.255 38.060 105.425 39.100 ;
        RECT 110.525 38.660 111.025 38.830 ;
        RECT 112.455 38.660 112.955 38.830 ;
        RECT 105.485 37.720 105.985 37.890 ;
        RECT 105.335 35.540 105.835 35.710 ;
        RECT 105.105 33.285 105.275 35.325 ;
        RECT 111.085 33.405 111.255 38.445 ;
        RECT 112.225 33.405 112.395 38.445 ;
        RECT 116.455 38.100 116.625 39.140 ;
        RECT 121.735 38.680 122.235 38.850 ;
        RECT 123.665 38.680 124.165 38.850 ;
        RECT 116.685 37.760 117.185 37.930 ;
        RECT 116.535 35.580 117.035 35.750 ;
        RECT 116.305 33.325 116.475 35.365 ;
        RECT 122.295 33.425 122.465 38.465 ;
        RECT 123.435 33.425 123.605 38.465 ;
        RECT 127.665 38.120 127.835 39.160 ;
        RECT 127.895 37.780 128.395 37.950 ;
        RECT 127.745 35.600 128.245 35.770 ;
        RECT 127.515 33.345 127.685 35.385 ;
        RECT 20.595 32.970 21.095 33.140 ;
        RECT 22.525 32.970 23.025 33.140 ;
        RECT 26.605 32.890 27.105 33.060 ;
        RECT 31.875 32.970 32.375 33.140 ;
        RECT 33.805 32.970 34.305 33.140 ;
        RECT 37.885 32.890 38.385 33.060 ;
        RECT 43.165 32.950 43.665 33.120 ;
        RECT 45.095 32.950 45.595 33.120 ;
        RECT 49.175 32.870 49.675 33.040 ;
        RECT 54.385 32.950 54.885 33.120 ;
        RECT 56.315 32.950 56.815 33.120 ;
        RECT 60.395 32.870 60.895 33.040 ;
        RECT 65.585 32.950 66.085 33.120 ;
        RECT 67.515 32.950 68.015 33.120 ;
        RECT 71.595 32.870 72.095 33.040 ;
        RECT 76.875 32.940 77.375 33.110 ;
        RECT 78.805 32.940 79.305 33.110 ;
        RECT 82.885 32.860 83.385 33.030 ;
        RECT 88.115 32.960 88.615 33.130 ;
        RECT 90.045 32.960 90.545 33.130 ;
        RECT 94.125 32.880 94.625 33.050 ;
        RECT 99.325 32.980 99.825 33.150 ;
        RECT 101.255 32.980 101.755 33.150 ;
        RECT 105.335 32.900 105.835 33.070 ;
        RECT 110.525 33.020 111.025 33.190 ;
        RECT 112.455 33.020 112.955 33.190 ;
        RECT 116.535 32.940 117.035 33.110 ;
        RECT 121.735 33.040 122.235 33.210 ;
        RECT 123.665 33.040 124.165 33.210 ;
        RECT 127.745 32.960 128.245 33.130 ;
        RECT 19.615 20.070 19.785 30.110 ;
        RECT 20.905 20.070 21.075 30.110 ;
        RECT 22.045 20.070 22.215 30.110 ;
        RECT 30.895 20.070 31.065 30.110 ;
        RECT 32.185 20.070 32.355 30.110 ;
        RECT 33.325 20.070 33.495 30.110 ;
        RECT 42.185 20.050 42.355 30.090 ;
        RECT 43.475 20.050 43.645 30.090 ;
        RECT 44.615 20.050 44.785 30.090 ;
        RECT 53.405 20.050 53.575 30.090 ;
        RECT 54.695 20.050 54.865 30.090 ;
        RECT 55.835 20.050 56.005 30.090 ;
        RECT 64.605 20.050 64.775 30.090 ;
        RECT 65.895 20.050 66.065 30.090 ;
        RECT 67.035 20.050 67.205 30.090 ;
        RECT 75.895 20.040 76.065 30.080 ;
        RECT 77.185 20.040 77.355 30.080 ;
        RECT 78.325 20.040 78.495 30.080 ;
        RECT 87.135 20.060 87.305 30.100 ;
        RECT 88.425 20.060 88.595 30.100 ;
        RECT 89.565 20.060 89.735 30.100 ;
        RECT 98.345 20.080 98.515 30.120 ;
        RECT 99.635 20.080 99.805 30.120 ;
        RECT 100.775 20.080 100.945 30.120 ;
        RECT 109.545 20.120 109.715 30.160 ;
        RECT 110.835 20.120 111.005 30.160 ;
        RECT 111.975 20.120 112.145 30.160 ;
        RECT 120.755 20.140 120.925 30.180 ;
        RECT 122.045 20.140 122.215 30.180 ;
        RECT 123.185 20.140 123.355 30.180 ;
      LAYER met1 ;
        RECT 80.065 207.450 80.355 207.495 ;
        RECT 80.970 207.450 81.290 207.510 ;
        RECT 80.065 207.310 81.290 207.450 ;
        RECT 80.065 207.265 80.355 207.310 ;
        RECT 80.970 207.250 81.290 207.310 ;
        RECT 71.310 207.110 71.630 207.170 ;
        RECT 74.545 207.110 74.835 207.155 ;
        RECT 71.310 206.970 74.835 207.110 ;
        RECT 71.310 206.910 71.630 206.970 ;
        RECT 74.545 206.925 74.835 206.970 ;
        RECT 75.450 207.110 75.770 207.170 ;
        RECT 79.605 207.110 79.895 207.155 ;
        RECT 75.450 206.970 79.895 207.110 ;
        RECT 75.450 206.910 75.770 206.970 ;
        RECT 79.605 206.925 79.895 206.970 ;
        RECT 74.990 206.230 75.310 206.490 ;
        RECT 75.910 206.430 76.230 206.490 ;
        RECT 77.765 206.430 78.055 206.475 ;
        RECT 75.910 206.290 78.055 206.430 ;
        RECT 75.910 206.230 76.230 206.290 ;
        RECT 77.765 206.245 78.055 206.290 ;
        RECT 71.310 205.410 71.630 205.470 ;
        RECT 69.100 205.270 71.630 205.410 ;
        RECT 66.265 204.730 66.555 204.775 ;
        RECT 67.185 204.730 67.475 204.775 ;
        RECT 69.100 204.730 69.240 205.270 ;
        RECT 71.310 205.210 71.630 205.270 ;
        RECT 74.990 205.410 75.310 205.470 ;
        RECT 74.990 205.270 76.600 205.410 ;
        RECT 74.990 205.210 75.310 205.270 ;
        RECT 70.045 205.070 70.335 205.115 ;
        RECT 73.285 205.070 73.935 205.115 ;
        RECT 70.045 204.930 73.935 205.070 ;
        RECT 70.045 204.885 70.635 204.930 ;
        RECT 73.285 204.885 73.935 204.930 ;
        RECT 66.265 204.590 69.240 204.730 ;
        RECT 66.265 204.545 66.555 204.590 ;
        RECT 67.185 204.545 67.475 204.590 ;
        RECT 70.345 204.570 70.635 204.885 ;
        RECT 75.910 204.870 76.230 205.130 ;
        RECT 76.460 205.070 76.600 205.270 ;
        RECT 79.245 205.070 79.535 205.115 ;
        RECT 82.485 205.070 83.135 205.115 ;
        RECT 76.460 204.930 83.135 205.070 ;
        RECT 79.245 204.885 79.835 204.930 ;
        RECT 82.485 204.885 83.135 204.930 ;
        RECT 71.425 204.730 71.715 204.775 ;
        RECT 75.005 204.730 75.295 204.775 ;
        RECT 76.840 204.730 77.130 204.775 ;
        RECT 71.425 204.590 77.130 204.730 ;
        RECT 67.645 204.390 67.935 204.435 ;
        RECT 70.480 204.390 70.620 204.570 ;
        RECT 71.425 204.545 71.715 204.590 ;
        RECT 75.005 204.545 75.295 204.590 ;
        RECT 76.840 204.545 77.130 204.590 ;
        RECT 79.545 204.570 79.835 204.885 ;
        RECT 80.625 204.730 80.915 204.775 ;
        RECT 84.205 204.730 84.495 204.775 ;
        RECT 86.040 204.730 86.330 204.775 ;
        RECT 80.625 204.590 86.330 204.730 ;
        RECT 80.625 204.545 80.915 204.590 ;
        RECT 84.205 204.545 84.495 204.590 ;
        RECT 86.040 204.545 86.330 204.590 ;
        RECT 67.645 204.250 70.620 204.390 ;
        RECT 77.305 204.390 77.595 204.435 ;
        RECT 86.505 204.390 86.795 204.435 ;
        RECT 88.330 204.390 88.650 204.450 ;
        RECT 77.305 204.250 88.650 204.390 ;
        RECT 67.645 204.205 67.935 204.250 ;
        RECT 77.305 204.205 77.595 204.250 ;
        RECT 86.505 204.205 86.795 204.250 ;
        RECT 88.330 204.190 88.650 204.250 ;
        RECT 71.425 204.050 71.715 204.095 ;
        RECT 74.545 204.050 74.835 204.095 ;
        RECT 76.435 204.050 76.725 204.095 ;
        RECT 71.425 203.910 76.725 204.050 ;
        RECT 71.425 203.865 71.715 203.910 ;
        RECT 74.545 203.865 74.835 203.910 ;
        RECT 76.435 203.865 76.725 203.910 ;
        RECT 80.625 204.050 80.915 204.095 ;
        RECT 83.745 204.050 84.035 204.095 ;
        RECT 85.635 204.050 85.925 204.095 ;
        RECT 80.625 203.910 85.925 204.050 ;
        RECT 80.625 203.865 80.915 203.910 ;
        RECT 83.745 203.865 84.035 203.910 ;
        RECT 85.635 203.865 85.925 203.910 ;
        RECT 65.330 203.710 65.650 203.770 ;
        RECT 65.805 203.710 66.095 203.755 ;
        RECT 65.330 203.570 66.095 203.710 ;
        RECT 65.330 203.510 65.650 203.570 ;
        RECT 65.805 203.525 66.095 203.570 ;
        RECT 68.565 203.710 68.855 203.755 ;
        RECT 69.010 203.710 69.330 203.770 ;
        RECT 68.565 203.570 69.330 203.710 ;
        RECT 68.565 203.525 68.855 203.570 ;
        RECT 69.010 203.510 69.330 203.570 ;
        RECT 77.750 203.510 78.070 203.770 ;
        RECT 79.130 203.710 79.450 203.770 ;
        RECT 85.190 203.710 85.480 203.755 ;
        RECT 79.130 203.570 85.480 203.710 ;
        RECT 79.130 203.510 79.450 203.570 ;
        RECT 85.190 203.525 85.480 203.570 ;
        RECT 73.625 202.690 73.915 202.735 ;
        RECT 75.450 202.690 75.770 202.750 ;
        RECT 73.625 202.550 75.770 202.690 ;
        RECT 73.625 202.505 73.915 202.550 ;
        RECT 75.450 202.490 75.770 202.550 ;
        RECT 79.130 202.490 79.450 202.750 ;
        RECT 61.155 202.350 61.445 202.395 ;
        RECT 63.045 202.350 63.335 202.395 ;
        RECT 66.165 202.350 66.455 202.395 ;
        RECT 61.155 202.210 66.455 202.350 ;
        RECT 61.155 202.165 61.445 202.210 ;
        RECT 63.045 202.165 63.335 202.210 ;
        RECT 66.165 202.165 66.455 202.210 ;
        RECT 82.465 202.350 82.755 202.395 ;
        RECT 85.585 202.350 85.875 202.395 ;
        RECT 87.475 202.350 87.765 202.395 ;
        RECT 82.465 202.210 87.765 202.350 ;
        RECT 82.465 202.165 82.755 202.210 ;
        RECT 85.585 202.165 85.875 202.210 ;
        RECT 87.475 202.165 87.765 202.210 ;
        RECT 61.650 201.810 61.970 202.070 ;
        RECT 72.230 202.010 72.550 202.070 ;
        RECT 77.750 202.010 78.070 202.070 ;
        RECT 71.400 201.870 78.070 202.010 ;
        RECT 60.270 201.470 60.590 201.730 ;
        RECT 71.400 201.715 71.540 201.870 ;
        RECT 72.230 201.810 72.550 201.870 ;
        RECT 77.750 201.810 78.070 201.870 ;
        RECT 84.650 202.010 84.970 202.070 ;
        RECT 86.965 202.010 87.255 202.055 ;
        RECT 84.650 201.870 87.255 202.010 ;
        RECT 84.650 201.810 84.970 201.870 ;
        RECT 86.965 201.825 87.255 201.870 ;
        RECT 88.330 201.810 88.650 202.070 ;
        RECT 60.750 201.670 61.040 201.715 ;
        RECT 62.585 201.670 62.875 201.715 ;
        RECT 66.165 201.670 66.455 201.715 ;
        RECT 60.750 201.530 66.455 201.670 ;
        RECT 60.750 201.485 61.040 201.530 ;
        RECT 62.585 201.485 62.875 201.530 ;
        RECT 66.165 201.485 66.455 201.530 ;
        RECT 63.945 201.330 64.595 201.375 ;
        RECT 65.330 201.330 65.650 201.390 ;
        RECT 67.245 201.375 67.535 201.690 ;
        RECT 71.325 201.485 71.615 201.715 ;
        RECT 72.705 201.670 72.995 201.715 ;
        RECT 71.860 201.530 72.995 201.670 ;
        RECT 67.245 201.330 67.835 201.375 ;
        RECT 63.945 201.190 67.835 201.330 ;
        RECT 63.945 201.145 64.595 201.190 ;
        RECT 65.330 201.130 65.650 201.190 ;
        RECT 67.545 201.145 67.835 201.190 ;
        RECT 70.390 201.130 70.710 201.390 ;
        RECT 71.860 201.330 72.000 201.530 ;
        RECT 72.705 201.485 72.995 201.530 ;
        RECT 78.210 201.470 78.530 201.730 ;
        RECT 71.170 201.190 72.000 201.330 ;
        RECT 72.245 201.330 72.535 201.375 ;
        RECT 73.610 201.330 73.930 201.390 ;
        RECT 72.245 201.190 73.930 201.330 ;
        RECT 69.010 200.990 69.330 201.050 ;
        RECT 71.170 200.990 71.310 201.190 ;
        RECT 72.245 201.145 72.535 201.190 ;
        RECT 73.610 201.130 73.930 201.190 ;
        RECT 76.830 201.130 77.150 201.390 ;
        RECT 81.385 201.375 81.675 201.690 ;
        RECT 82.465 201.670 82.755 201.715 ;
        RECT 86.045 201.670 86.335 201.715 ;
        RECT 87.880 201.670 88.170 201.715 ;
        RECT 82.465 201.530 88.170 201.670 ;
        RECT 82.465 201.485 82.755 201.530 ;
        RECT 86.045 201.485 86.335 201.530 ;
        RECT 87.880 201.485 88.170 201.530 ;
        RECT 81.085 201.330 81.675 201.375 ;
        RECT 83.270 201.330 83.590 201.390 ;
        RECT 84.325 201.330 84.975 201.375 ;
        RECT 81.085 201.190 84.975 201.330 ;
        RECT 81.085 201.145 81.375 201.190 ;
        RECT 83.270 201.130 83.590 201.190 ;
        RECT 84.325 201.145 84.975 201.190 ;
        RECT 69.010 200.850 71.310 200.990 ;
        RECT 69.010 200.790 69.330 200.850 ;
        RECT 77.290 200.790 77.610 201.050 ;
        RECT 78.670 200.990 78.990 201.050 ;
        RECT 79.605 200.990 79.895 201.035 ;
        RECT 78.670 200.850 79.895 200.990 ;
        RECT 78.670 200.790 78.990 200.850 ;
        RECT 79.605 200.805 79.895 200.850 ;
        RECT 61.650 199.970 61.970 200.030 ;
        RECT 65.805 199.970 66.095 200.015 ;
        RECT 61.650 199.830 66.095 199.970 ;
        RECT 61.650 199.770 61.970 199.830 ;
        RECT 65.805 199.785 66.095 199.830 ;
        RECT 69.010 199.770 69.330 200.030 ;
        RECT 72.230 199.770 72.550 200.030 ;
        RECT 75.465 199.970 75.755 200.015 ;
        RECT 76.830 199.970 77.150 200.030 ;
        RECT 75.465 199.830 77.150 199.970 ;
        RECT 75.465 199.785 75.755 199.830 ;
        RECT 76.830 199.770 77.150 199.830 ;
        RECT 78.210 199.970 78.530 200.030 ;
        RECT 79.145 199.970 79.435 200.015 ;
        RECT 78.210 199.830 79.435 199.970 ;
        RECT 78.210 199.770 78.530 199.830 ;
        RECT 79.145 199.785 79.435 199.830 ;
        RECT 83.270 199.770 83.590 200.030 ;
        RECT 84.650 199.770 84.970 200.030 ;
        RECT 68.565 199.630 68.855 199.675 ;
        RECT 74.070 199.630 74.390 199.690 ;
        RECT 74.545 199.630 74.835 199.675 ;
        RECT 68.565 199.490 71.310 199.630 ;
        RECT 68.565 199.445 68.855 199.490 ;
        RECT 66.710 199.090 67.030 199.350 ;
        RECT 70.390 199.090 70.710 199.350 ;
        RECT 71.170 199.290 71.310 199.490 ;
        RECT 74.070 199.490 74.835 199.630 ;
        RECT 74.070 199.430 74.390 199.490 ;
        RECT 74.545 199.445 74.835 199.490 ;
        RECT 75.910 199.630 76.230 199.690 ;
        RECT 79.905 199.630 80.195 199.675 ;
        RECT 75.910 199.490 80.195 199.630 ;
        RECT 75.910 199.430 76.230 199.490 ;
        RECT 79.905 199.445 80.195 199.490 ;
        RECT 80.970 199.630 81.290 199.690 ;
        RECT 81.905 199.630 82.195 199.675 ;
        RECT 80.970 199.490 82.195 199.630 ;
        RECT 80.970 199.430 81.290 199.490 ;
        RECT 81.905 199.445 82.195 199.490 ;
        RECT 71.785 199.290 72.075 199.335 ;
        RECT 78.670 199.290 78.990 199.350 ;
        RECT 71.170 199.150 78.990 199.290 ;
        RECT 71.785 199.105 72.075 199.150 ;
        RECT 78.670 199.090 78.990 199.150 ;
        RECT 81.445 199.105 81.735 199.335 ;
        RECT 82.365 199.105 82.655 199.335 ;
        RECT 67.980 198.950 68.270 198.995 ;
        RECT 72.230 198.950 72.550 199.010 ;
        RECT 67.980 198.810 72.550 198.950 ;
        RECT 67.980 198.765 68.270 198.810 ;
        RECT 72.230 198.750 72.550 198.810 ;
        RECT 77.750 198.950 78.070 199.010 ;
        RECT 81.520 198.950 81.660 199.105 ;
        RECT 77.750 198.810 81.660 198.950 ;
        RECT 82.440 198.950 82.580 199.105 ;
        RECT 83.730 199.090 84.050 199.350 ;
        RECT 84.205 199.105 84.495 199.335 ;
        RECT 84.280 198.950 84.420 199.105 ;
        RECT 82.440 198.810 84.420 198.950 ;
        RECT 77.750 198.750 78.070 198.810 ;
        RECT 70.390 198.610 70.710 198.670 ;
        RECT 74.070 198.610 74.390 198.670 ;
        RECT 70.390 198.470 74.390 198.610 ;
        RECT 70.390 198.410 70.710 198.470 ;
        RECT 74.070 198.410 74.390 198.470 ;
        RECT 74.545 198.610 74.835 198.655 ;
        RECT 75.450 198.610 75.770 198.670 ;
        RECT 74.545 198.470 75.770 198.610 ;
        RECT 74.545 198.425 74.835 198.470 ;
        RECT 75.450 198.410 75.770 198.470 ;
        RECT 77.290 198.610 77.610 198.670 ;
        RECT 82.440 198.610 82.580 198.810 ;
        RECT 77.290 198.470 82.580 198.610 ;
        RECT 77.290 198.410 77.610 198.470 ;
        RECT 67.185 198.270 67.475 198.315 ;
        RECT 67.630 198.270 67.950 198.330 ;
        RECT 67.185 198.130 67.950 198.270 ;
        RECT 67.185 198.085 67.475 198.130 ;
        RECT 67.630 198.070 67.950 198.130 ;
        RECT 70.850 198.070 71.170 198.330 ;
        RECT 80.050 198.070 80.370 198.330 ;
        RECT 66.710 197.250 67.030 197.310 ;
        RECT 69.485 197.250 69.775 197.295 ;
        RECT 66.710 197.110 69.775 197.250 ;
        RECT 66.710 197.050 67.030 197.110 ;
        RECT 69.485 197.065 69.775 197.110 ;
        RECT 70.390 197.050 70.710 197.310 ;
        RECT 79.145 197.250 79.435 197.295 ;
        RECT 80.050 197.250 80.370 197.310 ;
        RECT 79.145 197.110 80.370 197.250 ;
        RECT 79.145 197.065 79.435 197.110 ;
        RECT 80.050 197.050 80.370 197.110 ;
        RECT 76.370 196.910 76.690 196.970 ;
        RECT 77.750 196.910 78.070 196.970 ;
        RECT 73.700 196.770 78.070 196.910 ;
        RECT 73.700 196.630 73.840 196.770 ;
        RECT 76.370 196.710 76.690 196.770 ;
        RECT 77.750 196.710 78.070 196.770 ;
        RECT 111.905 196.910 112.195 196.955 ;
        RECT 115.025 196.910 115.315 196.955 ;
        RECT 116.915 196.910 117.205 196.955 ;
        RECT 111.905 196.770 117.205 196.910 ;
        RECT 111.905 196.725 112.195 196.770 ;
        RECT 115.025 196.725 115.315 196.770 ;
        RECT 116.915 196.725 117.205 196.770 ;
        RECT 73.150 196.370 73.470 196.630 ;
        RECT 73.610 196.370 73.930 196.630 ;
        RECT 74.070 196.370 74.390 196.630 ;
        RECT 53.385 196.230 53.675 196.275 ;
        RECT 55.210 196.230 55.530 196.290 ;
        RECT 56.605 196.230 56.895 196.275 ;
        RECT 53.385 196.090 56.895 196.230 ;
        RECT 53.385 196.045 53.675 196.090 ;
        RECT 55.210 196.030 55.530 196.090 ;
        RECT 56.605 196.045 56.895 196.090 ;
        RECT 72.705 196.230 72.995 196.275 ;
        RECT 75.450 196.230 75.770 196.290 ;
        RECT 72.705 196.090 75.770 196.230 ;
        RECT 72.705 196.045 72.995 196.090 ;
        RECT 75.450 196.030 75.770 196.090 ;
        RECT 77.750 196.230 78.070 196.290 ;
        RECT 78.225 196.230 78.515 196.275 ;
        RECT 77.750 196.090 78.515 196.230 ;
        RECT 77.750 196.030 78.070 196.090 ;
        RECT 78.225 196.045 78.515 196.090 ;
        RECT 107.650 196.030 107.970 196.290 ;
        RECT 71.325 195.890 71.615 195.935 ;
        RECT 75.910 195.890 76.230 195.950 ;
        RECT 71.325 195.750 76.230 195.890 ;
        RECT 71.325 195.705 71.615 195.750 ;
        RECT 75.910 195.690 76.230 195.750 ;
        RECT 77.290 195.690 77.610 195.950 ;
        RECT 110.825 195.935 111.115 196.250 ;
        RECT 111.905 196.230 112.195 196.275 ;
        RECT 115.485 196.230 115.775 196.275 ;
        RECT 117.320 196.230 117.610 196.275 ;
        RECT 111.905 196.090 117.610 196.230 ;
        RECT 111.905 196.045 112.195 196.090 ;
        RECT 115.485 196.045 115.775 196.090 ;
        RECT 117.320 196.045 117.610 196.090 ;
        RECT 117.785 196.230 118.075 196.275 ;
        RECT 120.990 196.230 121.310 196.290 ;
        RECT 117.785 196.090 121.310 196.230 ;
        RECT 117.785 196.045 118.075 196.090 ;
        RECT 120.990 196.030 121.310 196.090 ;
        RECT 108.125 195.890 108.415 195.935 ;
        RECT 110.525 195.890 111.115 195.935 ;
        RECT 113.765 195.890 114.415 195.935 ;
        RECT 108.125 195.750 114.415 195.890 ;
        RECT 108.125 195.705 108.415 195.750 ;
        RECT 110.525 195.705 110.815 195.750 ;
        RECT 113.765 195.705 114.415 195.750 ;
        RECT 116.390 195.690 116.710 195.950 ;
        RECT 51.990 195.550 52.310 195.610 ;
        RECT 52.925 195.550 53.215 195.595 ;
        RECT 51.990 195.410 53.215 195.550 ;
        RECT 51.990 195.350 52.310 195.410 ;
        RECT 52.925 195.365 53.215 195.410 ;
        RECT 56.145 195.550 56.435 195.595 ;
        RECT 56.590 195.550 56.910 195.610 ;
        RECT 56.145 195.410 56.910 195.550 ;
        RECT 56.145 195.365 56.435 195.410 ;
        RECT 56.590 195.350 56.910 195.410 ;
        RECT 70.325 195.550 70.615 195.595 ;
        RECT 71.785 195.550 72.075 195.595 ;
        RECT 70.325 195.410 72.075 195.550 ;
        RECT 70.325 195.365 70.615 195.410 ;
        RECT 71.785 195.365 72.075 195.410 ;
        RECT 73.150 195.550 73.470 195.610 ;
        RECT 74.530 195.550 74.850 195.610 ;
        RECT 77.380 195.550 77.520 195.690 ;
        RECT 73.150 195.410 77.520 195.550 ;
        RECT 73.150 195.350 73.470 195.410 ;
        RECT 74.530 195.350 74.850 195.410 ;
        RECT 109.030 195.350 109.350 195.610 ;
        RECT 75.465 194.530 75.755 194.575 ;
        RECT 75.910 194.530 76.230 194.590 ;
        RECT 75.465 194.390 76.230 194.530 ;
        RECT 75.465 194.345 75.755 194.390 ;
        RECT 75.910 194.330 76.230 194.390 ;
        RECT 83.730 194.530 84.050 194.590 ;
        RECT 83.730 194.390 107.880 194.530 ;
        RECT 83.730 194.330 84.050 194.390 ;
        RECT 47.385 194.190 48.035 194.235 ;
        RECT 50.985 194.190 51.275 194.235 ;
        RECT 51.990 194.190 52.310 194.250 ;
        RECT 47.385 194.050 52.310 194.190 ;
        RECT 47.385 194.005 48.035 194.050 ;
        RECT 50.685 194.005 51.275 194.050 ;
        RECT 44.190 193.850 44.480 193.895 ;
        RECT 46.025 193.850 46.315 193.895 ;
        RECT 49.605 193.850 49.895 193.895 ;
        RECT 44.190 193.710 49.895 193.850 ;
        RECT 44.190 193.665 44.480 193.710 ;
        RECT 46.025 193.665 46.315 193.710 ;
        RECT 49.605 193.665 49.895 193.710 ;
        RECT 50.685 193.690 50.975 194.005 ;
        RECT 51.990 193.990 52.310 194.050 ;
        RECT 54.405 194.190 54.695 194.235 ;
        RECT 56.590 194.190 56.910 194.250 ;
        RECT 57.645 194.190 58.295 194.235 ;
        RECT 54.405 194.050 58.295 194.190 ;
        RECT 54.405 194.005 54.995 194.050 ;
        RECT 54.705 193.690 54.995 194.005 ;
        RECT 56.590 193.990 56.910 194.050 ;
        RECT 57.645 194.005 58.295 194.050 ;
        RECT 58.890 194.190 59.210 194.250 ;
        RECT 60.285 194.190 60.575 194.235 ;
        RECT 71.310 194.190 71.630 194.250 ;
        RECT 83.820 194.190 83.960 194.330 ;
        RECT 58.890 194.050 60.575 194.190 ;
        RECT 58.890 193.990 59.210 194.050 ;
        RECT 60.285 194.005 60.575 194.050 ;
        RECT 71.170 194.050 83.960 194.190 ;
        RECT 71.170 193.990 71.630 194.050 ;
        RECT 55.785 193.850 56.075 193.895 ;
        RECT 59.365 193.850 59.655 193.895 ;
        RECT 61.200 193.850 61.490 193.895 ;
        RECT 55.785 193.710 61.490 193.850 ;
        RECT 55.785 193.665 56.075 193.710 ;
        RECT 59.365 193.665 59.655 193.710 ;
        RECT 61.200 193.665 61.490 193.710 ;
        RECT 66.710 193.850 67.030 193.910 ;
        RECT 71.170 193.850 71.310 193.990 ;
        RECT 66.710 193.710 71.310 193.850 ;
        RECT 66.710 193.650 67.030 193.710 ;
        RECT 72.245 193.665 72.535 193.895 ;
        RECT 37.730 193.510 38.050 193.570 ;
        RECT 43.725 193.510 44.015 193.555 ;
        RECT 37.730 193.370 44.015 193.510 ;
        RECT 37.730 193.310 38.050 193.370 ;
        RECT 43.725 193.325 44.015 193.370 ;
        RECT 45.090 193.310 45.410 193.570 ;
        RECT 60.270 193.510 60.590 193.570 ;
        RECT 61.665 193.510 61.955 193.555 ;
        RECT 63.950 193.510 64.270 193.570 ;
        RECT 60.270 193.370 64.270 193.510 ;
        RECT 72.320 193.510 72.460 193.665 ;
        RECT 73.610 193.650 73.930 193.910 ;
        RECT 74.070 193.850 74.390 193.910 ;
        RECT 77.290 193.850 77.610 193.910 ;
        RECT 78.225 193.850 78.515 193.895 ;
        RECT 74.070 193.710 78.515 193.850 ;
        RECT 74.070 193.650 74.390 193.710 ;
        RECT 77.290 193.650 77.610 193.710 ;
        RECT 78.225 193.665 78.515 193.710 ;
        RECT 84.650 193.850 84.970 193.910 ;
        RECT 86.045 193.850 86.335 193.895 ;
        RECT 84.650 193.710 86.335 193.850 ;
        RECT 84.650 193.650 84.970 193.710 ;
        RECT 86.045 193.665 86.335 193.710 ;
        RECT 86.490 193.650 86.810 193.910 ;
        RECT 90.170 193.850 90.490 193.910 ;
        RECT 96.240 193.895 96.380 194.390 ;
        RECT 107.740 194.250 107.880 194.390 ;
        RECT 96.625 194.190 96.915 194.235 ;
        RECT 99.025 194.190 99.315 194.235 ;
        RECT 102.265 194.190 102.915 194.235 ;
        RECT 96.625 194.050 102.915 194.190 ;
        RECT 96.625 194.005 96.915 194.050 ;
        RECT 99.025 194.005 99.615 194.050 ;
        RECT 102.265 194.005 102.915 194.050 ;
        RECT 107.650 194.190 107.970 194.250 ;
        RECT 107.650 194.050 116.160 194.190 ;
        RECT 90.645 193.850 90.935 193.895 ;
        RECT 90.170 193.710 90.935 193.850 ;
        RECT 90.170 193.650 90.490 193.710 ;
        RECT 90.645 193.665 90.935 193.710 ;
        RECT 91.565 193.665 91.855 193.895 ;
        RECT 96.165 193.665 96.455 193.895 ;
        RECT 99.325 193.690 99.615 194.005 ;
        RECT 107.650 193.990 107.970 194.050 ;
        RECT 116.020 193.910 116.160 194.050 ;
        RECT 100.405 193.850 100.695 193.895 ;
        RECT 103.985 193.850 104.275 193.895 ;
        RECT 105.820 193.850 106.110 193.895 ;
        RECT 100.405 193.710 106.110 193.850 ;
        RECT 100.405 193.665 100.695 193.710 ;
        RECT 103.985 193.665 104.275 193.710 ;
        RECT 105.820 193.665 106.110 193.710 ;
        RECT 112.265 193.665 112.555 193.895 ;
        RECT 74.530 193.510 74.850 193.570 ;
        RECT 75.910 193.510 76.230 193.570 ;
        RECT 72.320 193.370 76.230 193.510 ;
        RECT 60.270 193.310 60.590 193.370 ;
        RECT 61.665 193.325 61.955 193.370 ;
        RECT 63.950 193.310 64.270 193.370 ;
        RECT 74.530 193.310 74.850 193.370 ;
        RECT 75.910 193.310 76.230 193.370 ;
        RECT 76.845 193.325 77.135 193.555 ;
        RECT 44.595 193.170 44.885 193.215 ;
        RECT 46.485 193.170 46.775 193.215 ;
        RECT 49.605 193.170 49.895 193.215 ;
        RECT 44.595 193.030 49.895 193.170 ;
        RECT 44.595 192.985 44.885 193.030 ;
        RECT 46.485 192.985 46.775 193.030 ;
        RECT 49.605 192.985 49.895 193.030 ;
        RECT 55.785 193.170 56.075 193.215 ;
        RECT 58.905 193.170 59.195 193.215 ;
        RECT 60.795 193.170 61.085 193.215 ;
        RECT 55.785 193.030 61.085 193.170 ;
        RECT 55.785 192.985 56.075 193.030 ;
        RECT 58.905 192.985 59.195 193.030 ;
        RECT 60.795 192.985 61.085 193.030 ;
        RECT 75.005 193.170 75.295 193.215 ;
        RECT 76.920 193.170 77.060 193.325 ;
        RECT 85.110 193.310 85.430 193.570 ;
        RECT 91.640 193.510 91.780 193.665 ;
        RECT 88.420 193.370 91.780 193.510 ;
        RECT 88.420 193.215 88.560 193.370 ;
        RECT 104.890 193.310 105.210 193.570 ;
        RECT 106.285 193.510 106.575 193.555 ;
        RECT 107.190 193.510 107.510 193.570 ;
        RECT 106.285 193.370 107.510 193.510 ;
        RECT 106.285 193.325 106.575 193.370 ;
        RECT 107.190 193.310 107.510 193.370 ;
        RECT 109.030 193.510 109.350 193.570 ;
        RECT 109.965 193.510 110.255 193.555 ;
        RECT 110.870 193.510 111.190 193.570 ;
        RECT 109.030 193.370 111.190 193.510 ;
        RECT 109.030 193.310 109.350 193.370 ;
        RECT 109.965 193.325 110.255 193.370 ;
        RECT 110.870 193.310 111.190 193.370 ;
        RECT 111.345 193.325 111.635 193.555 ;
        RECT 75.005 193.030 77.060 193.170 ;
        RECT 75.005 192.985 75.295 193.030 ;
        RECT 88.345 192.985 88.635 193.215 ;
        RECT 100.405 193.170 100.695 193.215 ;
        RECT 103.525 193.170 103.815 193.215 ;
        RECT 105.415 193.170 105.705 193.215 ;
        RECT 111.420 193.170 111.560 193.325 ;
        RECT 111.790 193.310 112.110 193.570 ;
        RECT 100.405 193.030 105.705 193.170 ;
        RECT 100.405 192.985 100.695 193.030 ;
        RECT 103.525 192.985 103.815 193.030 ;
        RECT 105.415 192.985 105.705 193.030 ;
        RECT 105.900 193.030 111.560 193.170 ;
        RECT 105.900 192.890 106.040 193.030 ;
        RECT 50.610 192.830 50.930 192.890 ;
        RECT 52.465 192.830 52.755 192.875 ;
        RECT 50.610 192.690 52.755 192.830 ;
        RECT 50.610 192.630 50.930 192.690 ;
        RECT 52.465 192.645 52.755 192.690 ;
        RECT 52.910 192.630 53.230 192.890 ;
        RECT 66.250 192.630 66.570 192.890 ;
        RECT 69.010 192.830 69.330 192.890 ;
        RECT 72.705 192.830 72.995 192.875 ;
        RECT 69.010 192.690 72.995 192.830 ;
        RECT 69.010 192.630 69.330 192.690 ;
        RECT 72.705 192.645 72.995 192.690 ;
        RECT 75.450 192.830 75.770 192.890 ;
        RECT 76.385 192.830 76.675 192.875 ;
        RECT 75.450 192.690 76.675 192.830 ;
        RECT 75.450 192.630 75.770 192.690 ;
        RECT 76.385 192.645 76.675 192.690 ;
        RECT 90.185 192.830 90.475 192.875 ;
        RECT 90.630 192.830 90.950 192.890 ;
        RECT 90.185 192.690 90.950 192.830 ;
        RECT 90.185 192.645 90.475 192.690 ;
        RECT 90.630 192.630 90.950 192.690 ;
        RECT 92.485 192.830 92.775 192.875 ;
        RECT 93.850 192.830 94.170 192.890 ;
        RECT 92.485 192.690 94.170 192.830 ;
        RECT 92.485 192.645 92.775 192.690 ;
        RECT 93.850 192.630 94.170 192.690 ;
        RECT 97.530 192.630 97.850 192.890 ;
        RECT 105.810 192.630 106.130 192.890 ;
        RECT 106.745 192.830 107.035 192.875 ;
        RECT 107.650 192.830 107.970 192.890 ;
        RECT 112.340 192.830 112.480 193.665 ;
        RECT 115.930 193.650 116.250 193.910 ;
        RECT 106.745 192.690 112.480 192.830 ;
        RECT 106.745 192.645 107.035 192.690 ;
        RECT 107.650 192.630 107.970 192.690 ;
        RECT 114.090 192.630 114.410 192.890 ;
        RECT 115.470 192.630 115.790 192.890 ;
        RECT 45.090 191.810 45.410 191.870 ;
        RECT 51.545 191.810 51.835 191.855 ;
        RECT 45.090 191.670 51.835 191.810 ;
        RECT 45.090 191.610 45.410 191.670 ;
        RECT 51.545 191.625 51.835 191.670 ;
        RECT 58.890 191.610 59.210 191.870 ;
        RECT 103.525 191.810 103.815 191.855 ;
        RECT 104.890 191.810 105.210 191.870 ;
        RECT 103.525 191.670 105.210 191.810 ;
        RECT 103.525 191.625 103.815 191.670 ;
        RECT 104.890 191.610 105.210 191.670 ;
        RECT 40.605 191.470 40.895 191.515 ;
        RECT 43.725 191.470 44.015 191.515 ;
        RECT 45.615 191.470 45.905 191.515 ;
        RECT 40.605 191.330 45.905 191.470 ;
        RECT 40.605 191.285 40.895 191.330 ;
        RECT 43.725 191.285 44.015 191.330 ;
        RECT 45.615 191.285 45.905 191.330 ;
        RECT 56.605 191.285 56.895 191.515 ;
        RECT 62.995 191.470 63.285 191.515 ;
        RECT 64.885 191.470 65.175 191.515 ;
        RECT 68.005 191.470 68.295 191.515 ;
        RECT 62.995 191.330 68.295 191.470 ;
        RECT 62.995 191.285 63.285 191.330 ;
        RECT 64.885 191.285 65.175 191.330 ;
        RECT 68.005 191.285 68.295 191.330 ;
        RECT 69.010 191.470 69.330 191.530 ;
        RECT 70.865 191.470 71.155 191.515 ;
        RECT 69.010 191.330 71.155 191.470 ;
        RECT 42.790 191.130 43.110 191.190 ;
        RECT 45.105 191.130 45.395 191.175 ;
        RECT 42.790 190.990 45.395 191.130 ;
        RECT 42.790 190.930 43.110 190.990 ;
        RECT 45.105 190.945 45.395 190.990 ;
        RECT 47.850 191.130 48.170 191.190 ;
        RECT 53.385 191.130 53.675 191.175 ;
        RECT 47.850 190.990 53.675 191.130 ;
        RECT 47.850 190.930 48.170 190.990 ;
        RECT 53.385 190.945 53.675 190.990 ;
        RECT 38.190 190.450 38.510 190.510 ;
        RECT 39.525 190.495 39.815 190.810 ;
        RECT 40.605 190.790 40.895 190.835 ;
        RECT 44.185 190.790 44.475 190.835 ;
        RECT 46.020 190.790 46.310 190.835 ;
        RECT 40.605 190.650 46.310 190.790 ;
        RECT 40.605 190.605 40.895 190.650 ;
        RECT 44.185 190.605 44.475 190.650 ;
        RECT 46.020 190.605 46.310 190.650 ;
        RECT 46.485 190.605 46.775 190.835 ;
        RECT 39.225 190.450 39.815 190.495 ;
        RECT 42.465 190.450 43.115 190.495 ;
        RECT 38.190 190.310 43.115 190.450 ;
        RECT 46.560 190.450 46.700 190.605 ;
        RECT 52.450 190.590 52.770 190.850 ;
        RECT 56.680 190.790 56.820 191.285 ;
        RECT 69.010 191.270 69.330 191.330 ;
        RECT 70.865 191.285 71.155 191.330 ;
        RECT 71.325 191.285 71.615 191.515 ;
        RECT 76.845 191.470 77.135 191.515 ;
        RECT 73.700 191.330 77.135 191.470 ;
        RECT 63.505 191.130 63.795 191.175 ;
        RECT 71.400 191.130 71.540 191.285 ;
        RECT 73.700 191.175 73.840 191.330 ;
        RECT 76.845 191.285 77.135 191.330 ;
        RECT 90.140 191.470 90.430 191.515 ;
        RECT 92.920 191.470 93.210 191.515 ;
        RECT 94.780 191.470 95.070 191.515 ;
        RECT 90.140 191.330 95.070 191.470 ;
        RECT 90.140 191.285 90.430 191.330 ;
        RECT 92.920 191.285 93.210 191.330 ;
        RECT 94.780 191.285 95.070 191.330 ;
        RECT 113.285 191.470 113.575 191.515 ;
        RECT 116.405 191.470 116.695 191.515 ;
        RECT 118.295 191.470 118.585 191.515 ;
        RECT 113.285 191.330 118.585 191.470 ;
        RECT 113.285 191.285 113.575 191.330 ;
        RECT 116.405 191.285 116.695 191.330 ;
        RECT 118.295 191.285 118.585 191.330 ;
        RECT 73.625 191.130 73.915 191.175 ;
        RECT 63.505 190.990 71.540 191.130 ;
        RECT 72.780 190.990 73.915 191.130 ;
        RECT 63.505 190.945 63.795 190.990 ;
        RECT 57.985 190.790 58.275 190.835 ;
        RECT 56.680 190.650 58.275 190.790 ;
        RECT 57.985 190.605 58.275 190.650 ;
        RECT 62.125 190.605 62.415 190.835 ;
        RECT 62.590 190.790 62.880 190.835 ;
        RECT 64.425 190.790 64.715 190.835 ;
        RECT 68.005 190.790 68.295 190.835 ;
        RECT 62.590 190.650 68.295 190.790 ;
        RECT 62.590 190.605 62.880 190.650 ;
        RECT 64.425 190.605 64.715 190.650 ;
        RECT 68.005 190.605 68.295 190.650 ;
        RECT 62.200 190.450 62.340 190.605 ;
        RECT 63.950 190.450 64.270 190.510 ;
        RECT 66.250 190.495 66.570 190.510 ;
        RECT 46.560 190.310 64.270 190.450 ;
        RECT 38.190 190.250 38.510 190.310 ;
        RECT 39.225 190.265 39.515 190.310 ;
        RECT 42.465 190.265 43.115 190.310 ;
        RECT 63.950 190.250 64.270 190.310 ;
        RECT 65.785 190.450 66.570 190.495 ;
        RECT 69.085 190.495 69.375 190.810 ;
        RECT 70.390 190.790 70.710 190.850 ;
        RECT 72.780 190.790 72.920 190.990 ;
        RECT 73.625 190.945 73.915 190.990 ;
        RECT 76.370 190.930 76.690 191.190 ;
        RECT 77.290 191.130 77.610 191.190 ;
        RECT 87.410 191.130 87.730 191.190 ;
        RECT 93.405 191.130 93.695 191.175 ;
        RECT 93.850 191.130 94.170 191.190 ;
        RECT 77.290 190.990 78.440 191.130 ;
        RECT 77.290 190.930 77.610 190.990 ;
        RECT 70.390 190.650 72.920 190.790 ;
        RECT 70.390 190.590 70.710 190.650 ;
        RECT 73.150 190.590 73.470 190.850 ;
        RECT 75.450 190.790 75.770 190.850 ;
        RECT 78.300 190.835 78.440 190.990 ;
        RECT 87.410 190.990 93.160 191.130 ;
        RECT 87.410 190.930 87.730 190.990 ;
        RECT 77.765 190.790 78.055 190.835 ;
        RECT 75.450 190.650 78.055 190.790 ;
        RECT 75.450 190.590 75.770 190.650 ;
        RECT 77.765 190.605 78.055 190.650 ;
        RECT 78.225 190.605 78.515 190.835 ;
        RECT 90.140 190.790 90.430 190.835 ;
        RECT 93.020 190.790 93.160 190.990 ;
        RECT 93.405 190.990 94.170 191.130 ;
        RECT 93.405 190.945 93.695 190.990 ;
        RECT 93.850 190.930 94.170 190.990 ;
        RECT 98.450 190.930 98.770 191.190 ;
        RECT 98.925 191.130 99.215 191.175 ;
        RECT 105.810 191.130 106.130 191.190 ;
        RECT 106.745 191.130 107.035 191.175 ;
        RECT 98.925 190.990 103.280 191.130 ;
        RECT 98.925 190.945 99.215 190.990 ;
        RECT 95.245 190.790 95.535 190.835 ;
        RECT 90.140 190.650 92.675 190.790 ;
        RECT 93.020 190.650 95.535 190.790 ;
        RECT 90.140 190.605 90.430 190.650 ;
        RECT 69.085 190.450 69.675 190.495 ;
        RECT 65.785 190.310 69.675 190.450 ;
        RECT 65.785 190.265 66.570 190.310 ;
        RECT 69.385 190.265 69.675 190.310 ;
        RECT 88.280 190.450 88.570 190.495 ;
        RECT 90.630 190.450 90.950 190.510 ;
        RECT 92.460 190.495 92.675 190.650 ;
        RECT 95.245 190.605 95.535 190.650 ;
        RECT 97.990 190.790 98.310 190.850 ;
        RECT 99.000 190.790 99.140 190.945 ;
        RECT 102.605 190.790 102.895 190.835 ;
        RECT 97.990 190.650 99.140 190.790 ;
        RECT 101.300 190.650 102.895 190.790 ;
        RECT 103.140 190.790 103.280 190.990 ;
        RECT 105.810 190.990 107.035 191.130 ;
        RECT 105.810 190.930 106.130 190.990 ;
        RECT 106.745 190.945 107.035 190.990 ;
        RECT 107.650 190.930 107.970 191.190 ;
        RECT 108.125 190.790 108.415 190.835 ;
        RECT 103.140 190.650 108.415 190.790 ;
        RECT 97.990 190.590 98.310 190.650 ;
        RECT 91.540 190.450 91.830 190.495 ;
        RECT 88.280 190.310 91.830 190.450 ;
        RECT 88.280 190.265 88.570 190.310 ;
        RECT 66.250 190.250 66.570 190.265 ;
        RECT 90.630 190.250 90.950 190.310 ;
        RECT 91.540 190.265 91.830 190.310 ;
        RECT 92.460 190.450 92.750 190.495 ;
        RECT 94.320 190.450 94.610 190.495 ;
        RECT 92.460 190.310 94.610 190.450 ;
        RECT 92.460 190.265 92.750 190.310 ;
        RECT 94.320 190.265 94.610 190.310 ;
        RECT 37.745 190.110 38.035 190.155 ;
        RECT 40.030 190.110 40.350 190.170 ;
        RECT 37.745 189.970 40.350 190.110 ;
        RECT 37.745 189.925 38.035 189.970 ;
        RECT 40.030 189.910 40.350 189.970 ;
        RECT 54.290 189.910 54.610 190.170 ;
        RECT 54.750 189.910 55.070 190.170 ;
        RECT 75.910 190.110 76.230 190.170 ;
        RECT 77.305 190.110 77.595 190.155 ;
        RECT 75.910 189.970 77.595 190.110 ;
        RECT 75.910 189.910 76.230 189.970 ;
        RECT 77.305 189.925 77.595 189.970 ;
        RECT 78.210 190.110 78.530 190.170 ;
        RECT 84.650 190.110 84.970 190.170 ;
        RECT 101.300 190.155 101.440 190.650 ;
        RECT 102.605 190.605 102.895 190.650 ;
        RECT 108.125 190.605 108.415 190.650 ;
        RECT 112.205 190.495 112.495 190.810 ;
        RECT 113.285 190.790 113.575 190.835 ;
        RECT 116.865 190.790 117.155 190.835 ;
        RECT 118.700 190.790 118.990 190.835 ;
        RECT 113.285 190.650 118.990 190.790 ;
        RECT 113.285 190.605 113.575 190.650 ;
        RECT 116.865 190.605 117.155 190.650 ;
        RECT 118.700 190.605 118.990 190.650 ;
        RECT 119.165 190.790 119.455 190.835 ;
        RECT 120.990 190.790 121.310 190.850 ;
        RECT 119.165 190.650 121.310 190.790 ;
        RECT 119.165 190.605 119.455 190.650 ;
        RECT 120.990 190.590 121.310 190.650 ;
        RECT 115.470 190.495 115.790 190.510 ;
        RECT 111.905 190.450 112.495 190.495 ;
        RECT 115.145 190.450 115.795 190.495 ;
        RECT 111.905 190.310 115.795 190.450 ;
        RECT 111.905 190.265 112.195 190.310 ;
        RECT 115.145 190.265 115.795 190.310 ;
        RECT 115.470 190.250 115.790 190.265 ;
        RECT 117.770 190.250 118.090 190.510 ;
        RECT 86.275 190.110 86.565 190.155 ;
        RECT 99.385 190.110 99.675 190.155 ;
        RECT 78.210 189.970 99.675 190.110 ;
        RECT 78.210 189.910 78.530 189.970 ;
        RECT 84.650 189.910 84.970 189.970 ;
        RECT 86.275 189.925 86.565 189.970 ;
        RECT 99.385 189.925 99.675 189.970 ;
        RECT 101.225 189.925 101.515 190.155 ;
        RECT 109.950 189.910 110.270 190.170 ;
        RECT 110.410 189.910 110.730 190.170 ;
        RECT 36.825 189.090 37.115 189.135 ;
        RECT 51.085 189.090 51.375 189.135 ;
        RECT 52.450 189.090 52.770 189.150 ;
        RECT 36.825 188.950 38.420 189.090 ;
        RECT 36.825 188.905 37.115 188.950 ;
        RECT 29.925 188.410 30.215 188.455 ;
        RECT 34.510 188.410 34.830 188.470 ;
        RECT 29.925 188.270 34.830 188.410 ;
        RECT 29.925 188.225 30.215 188.270 ;
        RECT 34.510 188.210 34.830 188.270 ;
        RECT 35.890 188.210 36.210 188.470 ;
        RECT 37.730 188.210 38.050 188.470 ;
        RECT 38.280 188.410 38.420 188.950 ;
        RECT 51.085 188.950 52.770 189.090 ;
        RECT 51.085 188.905 51.375 188.950 ;
        RECT 52.450 188.890 52.770 188.950 ;
        RECT 71.785 189.090 72.075 189.135 ;
        RECT 73.150 189.090 73.470 189.150 ;
        RECT 89.725 189.090 90.015 189.135 ;
        RECT 71.785 188.950 73.470 189.090 ;
        RECT 71.785 188.905 72.075 188.950 ;
        RECT 73.150 188.890 73.470 188.950 ;
        RECT 85.200 188.950 90.015 189.090 ;
        RECT 38.670 188.750 38.960 188.795 ;
        RECT 40.530 188.750 40.820 188.795 ;
        RECT 38.670 188.610 40.820 188.750 ;
        RECT 38.670 188.565 38.960 188.610 ;
        RECT 40.530 188.565 40.820 188.610 ;
        RECT 41.450 188.750 41.740 188.795 ;
        RECT 44.710 188.750 45.000 188.795 ;
        RECT 41.450 188.610 45.000 188.750 ;
        RECT 41.450 188.565 41.740 188.610 ;
        RECT 39.585 188.410 39.875 188.455 ;
        RECT 38.280 188.270 39.875 188.410 ;
        RECT 40.605 188.410 40.820 188.565 ;
        RECT 42.850 188.410 43.140 188.455 ;
        RECT 40.605 188.270 43.140 188.410 ;
        RECT 39.585 188.225 39.875 188.270 ;
        RECT 42.850 188.225 43.140 188.270 ;
        RECT 29.465 188.070 29.755 188.115 ;
        RECT 30.370 188.070 30.690 188.130 ;
        RECT 29.465 187.930 30.690 188.070 ;
        RECT 29.465 187.885 29.755 187.930 ;
        RECT 30.370 187.870 30.690 187.930 ;
        RECT 34.985 188.070 35.275 188.115 ;
        RECT 43.340 188.070 43.480 188.610 ;
        RECT 44.710 188.565 45.000 188.610 ;
        RECT 48.785 188.750 49.075 188.795 ;
        RECT 54.750 188.750 55.070 188.810 ;
        RECT 48.785 188.610 55.070 188.750 ;
        RECT 48.785 188.565 49.075 188.610 ;
        RECT 54.750 188.550 55.070 188.610 ;
        RECT 81.380 188.750 81.670 188.795 ;
        RECT 84.640 188.750 84.930 188.795 ;
        RECT 85.200 188.750 85.340 188.950 ;
        RECT 89.725 188.905 90.015 188.950 ;
        RECT 90.645 188.905 90.935 189.135 ;
        RECT 81.380 188.610 85.340 188.750 ;
        RECT 85.560 188.750 85.850 188.795 ;
        RECT 87.420 188.750 87.710 188.795 ;
        RECT 90.720 188.750 90.860 188.905 ;
        RECT 97.990 188.890 98.310 189.150 ;
        RECT 114.105 189.090 114.395 189.135 ;
        RECT 116.390 189.090 116.710 189.150 ;
        RECT 114.105 188.950 116.710 189.090 ;
        RECT 114.105 188.905 114.395 188.950 ;
        RECT 116.390 188.890 116.710 188.950 ;
        RECT 116.865 189.090 117.155 189.135 ;
        RECT 117.770 189.090 118.090 189.150 ;
        RECT 116.865 188.950 118.090 189.090 ;
        RECT 116.865 188.905 117.155 188.950 ;
        RECT 117.770 188.890 118.090 188.950 ;
        RECT 85.560 188.610 87.710 188.750 ;
        RECT 81.380 188.565 81.670 188.610 ;
        RECT 84.640 188.565 84.930 188.610 ;
        RECT 85.560 188.565 85.850 188.610 ;
        RECT 87.420 188.565 87.710 188.610 ;
        RECT 88.420 188.610 90.860 188.750 ;
        RECT 99.945 188.750 100.235 188.795 ;
        RECT 102.590 188.750 102.910 188.810 ;
        RECT 103.185 188.750 103.835 188.795 ;
        RECT 99.945 188.610 103.835 188.750 ;
        RECT 49.245 188.225 49.535 188.455 ;
        RECT 83.240 188.410 83.530 188.455 ;
        RECT 85.560 188.410 85.775 188.565 ;
        RECT 83.240 188.270 85.775 188.410 ;
        RECT 86.505 188.410 86.795 188.455 ;
        RECT 88.420 188.410 88.560 188.610 ;
        RECT 99.945 188.565 100.535 188.610 ;
        RECT 86.505 188.270 88.560 188.410 ;
        RECT 83.240 188.225 83.530 188.270 ;
        RECT 86.505 188.225 86.795 188.270 ;
        RECT 34.985 187.930 43.480 188.070 ;
        RECT 34.985 187.885 35.275 187.930 ;
        RECT 47.850 187.870 48.170 188.130 ;
        RECT 38.210 187.730 38.500 187.775 ;
        RECT 40.070 187.730 40.360 187.775 ;
        RECT 42.850 187.730 43.140 187.775 ;
        RECT 38.210 187.590 43.140 187.730 ;
        RECT 38.210 187.545 38.500 187.590 ;
        RECT 40.070 187.545 40.360 187.590 ;
        RECT 42.850 187.545 43.140 187.590 ;
        RECT 41.410 187.390 41.730 187.450 ;
        RECT 46.715 187.390 47.005 187.435 ;
        RECT 49.320 187.390 49.460 188.225 ;
        RECT 90.170 188.210 90.490 188.470 ;
        RECT 91.090 188.410 91.410 188.470 ;
        RECT 91.565 188.410 91.855 188.455 ;
        RECT 91.090 188.270 91.855 188.410 ;
        RECT 91.090 188.210 91.410 188.270 ;
        RECT 91.565 188.225 91.855 188.270 ;
        RECT 100.245 188.250 100.535 188.565 ;
        RECT 102.590 188.550 102.910 188.610 ;
        RECT 103.185 188.565 103.835 188.610 ;
        RECT 101.325 188.410 101.615 188.455 ;
        RECT 104.905 188.410 105.195 188.455 ;
        RECT 106.740 188.410 107.030 188.455 ;
        RECT 101.325 188.270 107.030 188.410 ;
        RECT 101.325 188.225 101.615 188.270 ;
        RECT 104.905 188.225 105.195 188.270 ;
        RECT 106.740 188.225 107.030 188.270 ;
        RECT 109.950 188.410 110.270 188.470 ;
        RECT 113.185 188.410 113.475 188.455 ;
        RECT 109.950 188.270 113.475 188.410 ;
        RECT 109.950 188.210 110.270 188.270 ;
        RECT 113.185 188.225 113.475 188.270 ;
        RECT 114.090 188.410 114.410 188.470 ;
        RECT 115.945 188.410 116.235 188.455 ;
        RECT 114.090 188.270 116.235 188.410 ;
        RECT 114.090 188.210 114.410 188.270 ;
        RECT 115.945 188.225 116.235 188.270 ;
        RECT 50.610 188.070 50.930 188.130 ;
        RECT 51.545 188.070 51.835 188.115 ;
        RECT 50.610 187.930 51.835 188.070 ;
        RECT 50.610 187.870 50.930 187.930 ;
        RECT 51.545 187.885 51.835 187.930 ;
        RECT 69.010 187.870 69.330 188.130 ;
        RECT 79.375 188.070 79.665 188.115 ;
        RECT 85.570 188.070 85.890 188.130 ;
        RECT 79.375 187.930 85.890 188.070 ;
        RECT 79.375 187.885 79.665 187.930 ;
        RECT 85.570 187.870 85.890 187.930 ;
        RECT 87.410 188.070 87.730 188.130 ;
        RECT 88.345 188.070 88.635 188.115 ;
        RECT 87.410 187.930 88.635 188.070 ;
        RECT 87.410 187.870 87.730 187.930 ;
        RECT 88.345 187.885 88.635 187.930 ;
        RECT 95.245 188.070 95.535 188.115 ;
        RECT 97.530 188.070 97.850 188.130 ;
        RECT 107.190 188.070 107.510 188.130 ;
        RECT 120.990 188.070 121.310 188.130 ;
        RECT 95.245 187.930 106.960 188.070 ;
        RECT 95.245 187.885 95.535 187.930 ;
        RECT 97.530 187.870 97.850 187.930 ;
        RECT 83.240 187.730 83.530 187.775 ;
        RECT 86.020 187.730 86.310 187.775 ;
        RECT 87.880 187.730 88.170 187.775 ;
        RECT 83.240 187.590 88.170 187.730 ;
        RECT 83.240 187.545 83.530 187.590 ;
        RECT 86.020 187.545 86.310 187.590 ;
        RECT 87.880 187.545 88.170 187.590 ;
        RECT 101.325 187.730 101.615 187.775 ;
        RECT 104.445 187.730 104.735 187.775 ;
        RECT 106.335 187.730 106.625 187.775 ;
        RECT 101.325 187.590 106.625 187.730 ;
        RECT 106.820 187.730 106.960 187.930 ;
        RECT 107.190 187.930 121.310 188.070 ;
        RECT 107.190 187.870 107.510 187.930 ;
        RECT 120.990 187.870 121.310 187.930 ;
        RECT 107.650 187.730 107.970 187.790 ;
        RECT 106.820 187.590 107.970 187.730 ;
        RECT 101.325 187.545 101.615 187.590 ;
        RECT 104.445 187.545 104.735 187.590 ;
        RECT 106.335 187.545 106.625 187.590 ;
        RECT 107.650 187.530 107.970 187.590 ;
        RECT 41.410 187.250 49.460 187.390 ;
        RECT 96.610 187.390 96.930 187.450 ;
        RECT 98.465 187.390 98.755 187.435 ;
        RECT 96.610 187.250 98.755 187.390 ;
        RECT 41.410 187.190 41.730 187.250 ;
        RECT 46.715 187.205 47.005 187.250 ;
        RECT 96.610 187.190 96.930 187.250 ;
        RECT 98.465 187.205 98.755 187.250 ;
        RECT 102.130 187.390 102.450 187.450 ;
        RECT 105.890 187.390 106.180 187.435 ;
        RECT 102.130 187.250 106.180 187.390 ;
        RECT 102.130 187.190 102.450 187.250 ;
        RECT 105.890 187.205 106.180 187.250 ;
        RECT 38.190 186.170 38.510 186.430 ;
        RECT 98.450 186.370 98.770 186.430 ;
        RECT 85.660 186.230 98.770 186.370 ;
        RECT 26.655 186.030 26.945 186.075 ;
        RECT 28.545 186.030 28.835 186.075 ;
        RECT 31.665 186.030 31.955 186.075 ;
        RECT 26.655 185.890 31.955 186.030 ;
        RECT 26.655 185.845 26.945 185.890 ;
        RECT 28.545 185.845 28.835 185.890 ;
        RECT 31.665 185.845 31.955 185.890 ;
        RECT 35.890 186.030 36.210 186.090 ;
        RECT 39.125 186.030 39.415 186.075 ;
        RECT 35.890 185.890 39.415 186.030 ;
        RECT 35.890 185.830 36.210 185.890 ;
        RECT 39.125 185.845 39.415 185.890 ;
        RECT 43.250 186.030 43.570 186.090 ;
        RECT 50.625 186.030 50.915 186.075 ;
        RECT 43.250 185.890 50.915 186.030 ;
        RECT 43.250 185.830 43.570 185.890 ;
        RECT 50.625 185.845 50.915 185.890 ;
        RECT 53.485 186.030 53.775 186.075 ;
        RECT 56.605 186.030 56.895 186.075 ;
        RECT 58.495 186.030 58.785 186.075 ;
        RECT 53.485 185.890 58.785 186.030 ;
        RECT 53.485 185.845 53.775 185.890 ;
        RECT 56.605 185.845 56.895 185.890 ;
        RECT 58.495 185.845 58.785 185.890 ;
        RECT 85.660 185.750 85.800 186.230 ;
        RECT 88.805 186.030 89.095 186.075 ;
        RECT 91.090 186.030 91.410 186.090 ;
        RECT 88.805 185.890 91.410 186.030 ;
        RECT 88.805 185.845 89.095 185.890 ;
        RECT 91.090 185.830 91.410 185.890 ;
        RECT 35.430 185.690 35.750 185.750 ;
        RECT 41.885 185.690 42.175 185.735 ;
        RECT 46.945 185.690 47.235 185.735 ;
        RECT 47.850 185.690 48.170 185.750 ;
        RECT 55.210 185.690 55.530 185.750 ;
        RECT 35.430 185.550 48.170 185.690 ;
        RECT 35.430 185.490 35.750 185.550 ;
        RECT 41.885 185.505 42.175 185.550 ;
        RECT 46.945 185.505 47.235 185.550 ;
        RECT 47.850 185.490 48.170 185.550 ;
        RECT 49.780 185.550 55.530 185.690 ;
        RECT 25.770 185.150 26.090 185.410 ;
        RECT 26.250 185.350 26.540 185.395 ;
        RECT 28.085 185.350 28.375 185.395 ;
        RECT 31.665 185.350 31.955 185.395 ;
        RECT 26.250 185.210 31.955 185.350 ;
        RECT 26.250 185.165 26.540 185.210 ;
        RECT 28.085 185.165 28.375 185.210 ;
        RECT 31.665 185.165 31.955 185.210 ;
        RECT 27.150 184.810 27.470 185.070 ;
        RECT 29.445 185.010 30.095 185.055 ;
        RECT 30.370 185.010 30.690 185.070 ;
        RECT 32.745 185.055 33.035 185.370 ;
        RECT 34.510 185.350 34.830 185.410 ;
        RECT 49.780 185.395 49.920 185.550 ;
        RECT 55.210 185.490 55.530 185.550 ;
        RECT 85.570 185.490 85.890 185.750 ;
        RECT 86.490 185.490 86.810 185.750 ;
        RECT 92.945 185.690 93.235 185.735 ;
        RECT 96.610 185.690 96.930 185.750 ;
        RECT 97.160 185.735 97.300 186.230 ;
        RECT 98.450 186.170 98.770 186.230 ;
        RECT 101.225 186.370 101.515 186.415 ;
        RECT 102.130 186.370 102.450 186.430 ;
        RECT 101.225 186.230 102.450 186.370 ;
        RECT 101.225 186.185 101.515 186.230 ;
        RECT 102.130 186.170 102.450 186.230 ;
        RECT 102.590 186.170 102.910 186.430 ;
        RECT 110.885 186.370 111.175 186.415 ;
        RECT 111.790 186.370 112.110 186.430 ;
        RECT 110.885 186.230 112.110 186.370 ;
        RECT 110.885 186.185 111.175 186.230 ;
        RECT 111.790 186.170 112.110 186.230 ;
        RECT 98.540 186.030 98.680 186.170 ;
        RECT 105.810 186.030 106.130 186.090 ;
        RECT 98.540 185.890 106.130 186.030 ;
        RECT 105.810 185.830 106.130 185.890 ;
        RECT 92.945 185.550 96.930 185.690 ;
        RECT 92.945 185.505 93.235 185.550 ;
        RECT 96.610 185.490 96.930 185.550 ;
        RECT 97.085 185.505 97.375 185.735 ;
        RECT 37.745 185.350 38.035 185.395 ;
        RECT 34.140 185.210 38.035 185.350 ;
        RECT 32.745 185.010 33.335 185.055 ;
        RECT 29.445 184.870 33.335 185.010 ;
        RECT 29.445 184.825 30.095 184.870 ;
        RECT 30.370 184.810 30.690 184.870 ;
        RECT 33.045 184.825 33.335 184.870 ;
        RECT 31.290 184.670 31.610 184.730 ;
        RECT 34.140 184.670 34.280 185.210 ;
        RECT 34.510 185.150 34.830 185.210 ;
        RECT 37.745 185.165 38.035 185.210 ;
        RECT 49.705 185.165 49.995 185.395 ;
        RECT 39.570 185.010 39.890 185.070 ;
        RECT 52.405 185.055 52.695 185.370 ;
        RECT 53.485 185.350 53.775 185.395 ;
        RECT 57.065 185.350 57.355 185.395 ;
        RECT 58.900 185.350 59.190 185.395 ;
        RECT 53.485 185.210 59.190 185.350 ;
        RECT 53.485 185.165 53.775 185.210 ;
        RECT 57.065 185.165 57.355 185.210 ;
        RECT 58.900 185.165 59.190 185.210 ;
        RECT 59.365 185.350 59.655 185.395 ;
        RECT 63.950 185.350 64.270 185.410 ;
        RECT 59.365 185.210 64.270 185.350 ;
        RECT 59.365 185.165 59.655 185.210 ;
        RECT 63.950 185.150 64.270 185.210 ;
        RECT 79.590 185.150 79.910 185.410 ;
        RECT 90.170 185.150 90.490 185.410 ;
        RECT 95.705 185.350 95.995 185.395 ;
        RECT 97.160 185.350 97.760 185.360 ;
        RECT 99.370 185.350 99.690 185.410 ;
        RECT 100.305 185.350 100.595 185.395 ;
        RECT 95.705 185.220 98.220 185.350 ;
        RECT 95.705 185.210 97.300 185.220 ;
        RECT 97.620 185.210 98.220 185.220 ;
        RECT 95.705 185.165 95.995 185.210 ;
        RECT 46.485 185.010 46.775 185.055 ;
        RECT 39.570 184.870 46.775 185.010 ;
        RECT 39.570 184.810 39.890 184.870 ;
        RECT 46.485 184.825 46.775 184.870 ;
        RECT 49.245 185.010 49.535 185.055 ;
        RECT 52.105 185.010 52.695 185.055 ;
        RECT 55.345 185.010 55.995 185.055 ;
        RECT 49.245 184.870 55.995 185.010 ;
        RECT 49.245 184.825 49.535 184.870 ;
        RECT 52.105 184.825 52.395 184.870 ;
        RECT 55.345 184.825 55.995 184.870 ;
        RECT 57.985 185.010 58.275 185.055 ;
        RECT 61.650 185.010 61.970 185.070 ;
        RECT 86.965 185.010 87.255 185.055 ;
        RECT 57.985 184.870 61.970 185.010 ;
        RECT 57.985 184.825 58.275 184.870 ;
        RECT 61.650 184.810 61.970 184.870 ;
        RECT 82.900 184.870 87.255 185.010 ;
        RECT 31.290 184.530 34.280 184.670 ;
        RECT 34.525 184.670 34.815 184.715 ;
        RECT 36.350 184.670 36.670 184.730 ;
        RECT 34.525 184.530 36.670 184.670 ;
        RECT 31.290 184.470 31.610 184.530 ;
        RECT 34.525 184.485 34.815 184.530 ;
        RECT 36.350 184.470 36.670 184.530 ;
        RECT 40.950 184.470 41.270 184.730 ;
        RECT 41.410 184.470 41.730 184.730 ;
        RECT 41.870 184.670 42.190 184.730 ;
        RECT 44.185 184.670 44.475 184.715 ;
        RECT 41.870 184.530 44.475 184.670 ;
        RECT 41.870 184.470 42.190 184.530 ;
        RECT 44.185 184.485 44.475 184.530 ;
        RECT 46.010 184.470 46.330 184.730 ;
        RECT 80.970 184.670 81.290 184.730 ;
        RECT 82.900 184.715 83.040 184.870 ;
        RECT 86.965 184.825 87.255 184.870 ;
        RECT 82.825 184.670 83.115 184.715 ;
        RECT 80.970 184.530 83.115 184.670 ;
        RECT 80.970 184.470 81.290 184.530 ;
        RECT 82.825 184.485 83.115 184.530 ;
        RECT 84.650 184.670 84.970 184.730 ;
        RECT 89.725 184.670 90.015 184.715 ;
        RECT 84.650 184.530 90.015 184.670 ;
        RECT 90.260 184.670 90.400 185.150 ;
        RECT 91.550 185.010 91.870 185.070 ;
        RECT 98.080 185.055 98.220 185.210 ;
        RECT 99.370 185.210 100.595 185.350 ;
        RECT 99.370 185.150 99.690 185.210 ;
        RECT 100.305 185.165 100.595 185.210 ;
        RECT 103.065 185.165 103.355 185.395 ;
        RECT 108.125 185.350 108.415 185.395 ;
        RECT 110.410 185.350 110.730 185.410 ;
        RECT 108.125 185.210 110.730 185.350 ;
        RECT 108.125 185.165 108.415 185.210 ;
        RECT 97.545 185.010 97.835 185.055 ;
        RECT 91.550 184.870 97.835 185.010 ;
        RECT 91.550 184.810 91.870 184.870 ;
        RECT 97.545 184.825 97.835 184.870 ;
        RECT 98.005 184.825 98.295 185.055 ;
        RECT 103.140 185.010 103.280 185.165 ;
        RECT 110.410 185.150 110.730 185.210 ;
        RECT 98.540 184.870 103.280 185.010 ;
        RECT 97.070 184.670 97.390 184.730 ;
        RECT 98.540 184.670 98.680 184.870 ;
        RECT 90.260 184.530 98.680 184.670 ;
        RECT 98.910 184.670 99.230 184.730 ;
        RECT 99.845 184.670 100.135 184.715 ;
        RECT 98.910 184.530 100.135 184.670 ;
        RECT 84.650 184.470 84.970 184.530 ;
        RECT 89.725 184.485 90.015 184.530 ;
        RECT 97.070 184.470 97.390 184.530 ;
        RECT 98.910 184.470 99.230 184.530 ;
        RECT 99.845 184.485 100.135 184.530 ;
        RECT 23.025 183.650 23.315 183.695 ;
        RECT 27.150 183.650 27.470 183.710 ;
        RECT 23.025 183.510 27.470 183.650 ;
        RECT 23.025 183.465 23.315 183.510 ;
        RECT 27.150 183.450 27.470 183.510 ;
        RECT 42.790 183.450 43.110 183.710 ;
        RECT 46.010 183.650 46.330 183.710 ;
        RECT 46.485 183.650 46.775 183.695 ;
        RECT 46.010 183.510 46.775 183.650 ;
        RECT 46.010 183.450 46.330 183.510 ;
        RECT 46.485 183.465 46.775 183.510 ;
        RECT 61.650 183.450 61.970 183.710 ;
        RECT 76.370 183.650 76.690 183.710 ;
        RECT 90.185 183.650 90.475 183.695 ;
        RECT 74.160 183.510 76.690 183.650 ;
        RECT 30.385 183.310 30.675 183.355 ;
        RECT 32.685 183.310 32.975 183.355 ;
        RECT 34.050 183.310 34.370 183.370 ;
        RECT 30.385 183.170 34.370 183.310 ;
        RECT 30.385 183.125 30.675 183.170 ;
        RECT 32.685 183.125 32.975 183.170 ;
        RECT 34.050 183.110 34.370 183.170 ;
        RECT 50.165 183.310 50.455 183.355 ;
        RECT 50.165 183.170 62.800 183.310 ;
        RECT 50.165 183.125 50.455 183.170 ;
        RECT 22.105 182.970 22.395 183.015 ;
        RECT 23.485 182.970 23.775 183.015 ;
        RECT 22.105 182.830 23.775 182.970 ;
        RECT 22.105 182.785 22.395 182.830 ;
        RECT 23.485 182.785 23.775 182.830 ;
        RECT 27.625 182.970 27.915 183.015 ;
        RECT 34.510 182.970 34.830 183.030 ;
        RECT 27.625 182.830 34.830 182.970 ;
        RECT 27.625 182.785 27.915 182.830 ;
        RECT 34.510 182.770 34.830 182.830 ;
        RECT 41.870 182.770 42.190 183.030 ;
        RECT 49.690 182.970 50.010 183.030 ;
        RECT 52.465 182.970 52.755 183.015 ;
        RECT 43.340 182.830 48.080 182.970 ;
        RECT 43.340 182.690 43.480 182.830 ;
        RECT 26.705 182.445 26.995 182.675 ;
        RECT 33.145 182.445 33.435 182.675 ;
        RECT 34.065 182.630 34.355 182.675 ;
        RECT 35.430 182.630 35.750 182.690 ;
        RECT 34.065 182.490 35.750 182.630 ;
        RECT 34.065 182.445 34.355 182.490 ;
        RECT 26.780 182.290 26.920 182.445 ;
        RECT 30.845 182.290 31.135 182.335 ;
        RECT 26.780 182.150 31.135 182.290 ;
        RECT 33.220 182.290 33.360 182.445 ;
        RECT 35.430 182.430 35.750 182.490 ;
        RECT 38.205 182.630 38.495 182.675 ;
        RECT 40.030 182.630 40.350 182.690 ;
        RECT 38.205 182.490 40.350 182.630 ;
        RECT 38.205 182.445 38.495 182.490 ;
        RECT 40.030 182.430 40.350 182.490 ;
        RECT 43.250 182.430 43.570 182.690 ;
        RECT 47.405 182.445 47.695 182.675 ;
        RECT 47.940 182.630 48.080 182.830 ;
        RECT 49.690 182.830 52.755 182.970 ;
        RECT 49.690 182.770 50.010 182.830 ;
        RECT 52.465 182.785 52.755 182.830 ;
        RECT 55.210 182.970 55.530 183.030 ;
        RECT 56.590 182.970 56.910 183.030 ;
        RECT 62.660 183.015 62.800 183.170 ;
        RECT 55.210 182.830 56.910 182.970 ;
        RECT 55.210 182.770 55.530 182.830 ;
        RECT 56.590 182.770 56.910 182.830 ;
        RECT 59.825 182.970 60.115 183.015 ;
        RECT 60.285 182.970 60.575 183.015 ;
        RECT 59.825 182.830 60.575 182.970 ;
        RECT 59.825 182.785 60.115 182.830 ;
        RECT 60.285 182.785 60.575 182.830 ;
        RECT 62.585 182.785 62.875 183.015 ;
        RECT 73.610 182.770 73.930 183.030 ;
        RECT 74.160 183.015 74.300 183.510 ;
        RECT 76.370 183.450 76.690 183.510 ;
        RECT 87.040 183.510 90.475 183.650 ;
        RECT 75.450 183.310 75.770 183.370 ;
        RECT 84.650 183.355 84.970 183.370 ;
        RECT 87.040 183.355 87.180 183.510 ;
        RECT 90.185 183.465 90.475 183.510 ;
        RECT 90.630 183.650 90.950 183.710 ;
        RECT 91.550 183.650 91.870 183.710 ;
        RECT 92.485 183.650 92.775 183.695 ;
        RECT 90.630 183.510 92.775 183.650 ;
        RECT 90.630 183.450 90.950 183.510 ;
        RECT 91.550 183.450 91.870 183.510 ;
        RECT 92.485 183.465 92.775 183.510 ;
        RECT 96.610 183.650 96.930 183.710 ;
        RECT 101.210 183.650 101.530 183.710 ;
        RECT 104.905 183.650 105.195 183.695 ;
        RECT 96.610 183.510 105.195 183.650 ;
        RECT 96.610 183.450 96.930 183.510 ;
        RECT 101.210 183.450 101.530 183.510 ;
        RECT 104.905 183.465 105.195 183.510 ;
        RECT 109.490 183.650 109.810 183.710 ;
        RECT 111.805 183.650 112.095 183.695 ;
        RECT 109.490 183.510 112.095 183.650 ;
        RECT 109.490 183.450 109.810 183.510 ;
        RECT 111.805 183.465 112.095 183.510 ;
        RECT 81.085 183.310 81.375 183.355 ;
        RECT 84.325 183.310 84.975 183.355 ;
        RECT 75.450 183.170 77.520 183.310 ;
        RECT 75.450 183.110 75.770 183.170 ;
        RECT 74.085 182.785 74.375 183.015 ;
        RECT 74.545 182.970 74.835 183.015 ;
        RECT 74.990 182.970 75.310 183.030 ;
        RECT 74.545 182.830 75.310 182.970 ;
        RECT 74.545 182.785 74.835 182.830 ;
        RECT 52.925 182.630 53.215 182.675 ;
        RECT 47.940 182.490 53.215 182.630 ;
        RECT 52.925 182.445 53.215 182.490 ;
        RECT 53.385 182.445 53.675 182.675 ;
        RECT 36.350 182.290 36.670 182.350 ;
        RECT 33.220 182.150 36.670 182.290 ;
        RECT 30.845 182.105 31.135 182.150 ;
        RECT 36.350 182.090 36.670 182.150 ;
        RECT 41.870 182.290 42.190 182.350 ;
        RECT 43.340 182.290 43.480 182.430 ;
        RECT 41.870 182.150 43.480 182.290 ;
        RECT 47.480 182.290 47.620 182.445 ;
        RECT 50.625 182.290 50.915 182.335 ;
        RECT 53.460 182.290 53.600 182.445 ;
        RECT 57.050 182.430 57.370 182.690 ;
        RECT 65.790 182.630 66.110 182.690 ;
        RECT 69.010 182.630 69.330 182.690 ;
        RECT 73.165 182.630 73.455 182.675 ;
        RECT 65.790 182.490 73.455 182.630 ;
        RECT 65.790 182.430 66.110 182.490 ;
        RECT 69.010 182.430 69.330 182.490 ;
        RECT 73.165 182.445 73.455 182.490 ;
        RECT 56.130 182.290 56.450 182.350 ;
        RECT 47.480 182.150 50.915 182.290 ;
        RECT 41.870 182.090 42.190 182.150 ;
        RECT 50.625 182.105 50.915 182.150 ;
        RECT 53.000 182.150 56.450 182.290 ;
        RECT 39.570 181.950 39.890 182.010 ;
        RECT 40.965 181.950 41.255 181.995 ;
        RECT 39.570 181.810 41.255 181.950 ;
        RECT 39.570 181.750 39.890 181.810 ;
        RECT 40.965 181.765 41.255 181.810 ;
        RECT 47.850 181.950 48.170 182.010 ;
        RECT 53.000 181.950 53.140 182.150 ;
        RECT 56.130 182.090 56.450 182.150 ;
        RECT 69.470 182.290 69.790 182.350 ;
        RECT 71.310 182.290 71.630 182.350 ;
        RECT 74.620 182.290 74.760 182.785 ;
        RECT 74.990 182.770 75.310 182.830 ;
        RECT 75.925 182.970 76.215 183.015 ;
        RECT 76.370 182.970 76.690 183.030 ;
        RECT 77.380 183.015 77.520 183.170 ;
        RECT 81.085 183.170 84.975 183.310 ;
        RECT 81.085 183.125 81.675 183.170 ;
        RECT 84.325 183.125 84.975 183.170 ;
        RECT 86.965 183.125 87.255 183.355 ;
        RECT 87.410 183.310 87.730 183.370 ;
        RECT 93.965 183.310 94.255 183.355 ;
        RECT 96.150 183.310 96.470 183.370 ;
        RECT 97.205 183.310 97.855 183.355 ;
        RECT 87.410 183.170 88.560 183.310 ;
        RECT 75.925 182.830 76.690 182.970 ;
        RECT 75.925 182.785 76.215 182.830 ;
        RECT 76.370 182.770 76.690 182.830 ;
        RECT 76.845 182.785 77.135 183.015 ;
        RECT 77.305 182.785 77.595 183.015 ;
        RECT 76.920 182.630 77.060 182.785 ;
        RECT 77.750 182.770 78.070 183.030 ;
        RECT 81.385 182.810 81.675 183.125 ;
        RECT 84.650 183.110 84.970 183.125 ;
        RECT 87.410 183.110 87.730 183.170 ;
        RECT 88.420 183.015 88.560 183.170 ;
        RECT 93.965 183.170 97.855 183.310 ;
        RECT 93.965 183.125 94.555 183.170 ;
        RECT 82.465 182.970 82.755 183.015 ;
        RECT 86.045 182.970 86.335 183.015 ;
        RECT 87.880 182.970 88.170 183.015 ;
        RECT 82.465 182.830 88.170 182.970 ;
        RECT 82.465 182.785 82.755 182.830 ;
        RECT 86.045 182.785 86.335 182.830 ;
        RECT 87.880 182.785 88.170 182.830 ;
        RECT 88.345 182.785 88.635 183.015 ;
        RECT 79.590 182.630 79.910 182.690 ;
        RECT 76.920 182.490 79.910 182.630 ;
        RECT 88.420 182.630 88.560 182.785 ;
        RECT 91.090 182.770 91.410 183.030 ;
        RECT 94.265 182.810 94.555 183.125 ;
        RECT 96.150 183.110 96.470 183.170 ;
        RECT 97.205 183.125 97.855 183.170 ;
        RECT 99.830 183.110 100.150 183.370 ;
        RECT 116.965 183.310 117.255 183.355 ;
        RECT 120.205 183.310 120.855 183.355 ;
        RECT 116.965 183.170 120.855 183.310 ;
        RECT 116.965 183.125 117.555 183.170 ;
        RECT 120.205 183.125 120.855 183.170 ;
        RECT 122.845 183.310 123.135 183.355 ;
        RECT 124.210 183.310 124.530 183.370 ;
        RECT 122.845 183.170 124.530 183.310 ;
        RECT 122.845 183.125 123.135 183.170 ;
        RECT 117.265 183.030 117.555 183.125 ;
        RECT 124.210 183.110 124.530 183.170 ;
        RECT 95.345 182.970 95.635 183.015 ;
        RECT 98.925 182.970 99.215 183.015 ;
        RECT 100.760 182.970 101.050 183.015 ;
        RECT 95.345 182.830 101.050 182.970 ;
        RECT 95.345 182.785 95.635 182.830 ;
        RECT 98.925 182.785 99.215 182.830 ;
        RECT 100.760 182.785 101.050 182.830 ;
        RECT 104.445 182.785 104.735 183.015 ;
        RECT 111.790 182.970 112.110 183.030 ;
        RECT 112.265 182.970 112.555 183.015 ;
        RECT 111.790 182.830 112.555 182.970 ;
        RECT 101.225 182.630 101.515 182.675 ;
        RECT 88.420 182.490 101.515 182.630 ;
        RECT 79.590 182.430 79.910 182.490 ;
        RECT 101.225 182.445 101.515 182.490 ;
        RECT 77.290 182.290 77.610 182.350 ;
        RECT 69.470 182.150 77.610 182.290 ;
        RECT 69.470 182.090 69.790 182.150 ;
        RECT 71.310 182.090 71.630 182.150 ;
        RECT 73.240 182.010 73.380 182.150 ;
        RECT 77.290 182.090 77.610 182.150 ;
        RECT 82.465 182.290 82.755 182.335 ;
        RECT 85.585 182.290 85.875 182.335 ;
        RECT 87.475 182.290 87.765 182.335 ;
        RECT 82.465 182.150 87.765 182.290 ;
        RECT 82.465 182.105 82.755 182.150 ;
        RECT 85.585 182.105 85.875 182.150 ;
        RECT 87.475 182.105 87.765 182.150 ;
        RECT 95.345 182.290 95.635 182.335 ;
        RECT 98.465 182.290 98.755 182.335 ;
        RECT 100.355 182.290 100.645 182.335 ;
        RECT 95.345 182.150 100.645 182.290 ;
        RECT 95.345 182.105 95.635 182.150 ;
        RECT 98.465 182.105 98.755 182.150 ;
        RECT 100.355 182.105 100.645 182.150 ;
        RECT 47.850 181.810 53.140 181.950 ;
        RECT 47.850 181.750 48.170 181.810 ;
        RECT 55.670 181.750 55.990 182.010 ;
        RECT 61.190 181.750 61.510 182.010 ;
        RECT 72.245 181.950 72.535 181.995 ;
        RECT 72.690 181.950 73.010 182.010 ;
        RECT 72.245 181.810 73.010 181.950 ;
        RECT 72.245 181.765 72.535 181.810 ;
        RECT 72.690 181.750 73.010 181.810 ;
        RECT 73.150 181.750 73.470 182.010 ;
        RECT 79.130 181.750 79.450 182.010 ;
        RECT 83.270 181.950 83.590 182.010 ;
        RECT 91.090 181.950 91.410 182.010 ;
        RECT 83.270 181.810 91.410 181.950 ;
        RECT 83.270 181.750 83.590 181.810 ;
        RECT 91.090 181.750 91.410 181.810 ;
        RECT 94.770 181.950 95.090 182.010 ;
        RECT 102.605 181.950 102.895 181.995 ;
        RECT 94.770 181.810 102.895 181.950 ;
        RECT 104.520 181.950 104.660 182.785 ;
        RECT 111.790 182.770 112.110 182.830 ;
        RECT 112.265 182.785 112.555 182.830 ;
        RECT 117.265 182.810 117.630 183.030 ;
        RECT 117.310 182.770 117.630 182.810 ;
        RECT 118.345 182.970 118.635 183.015 ;
        RECT 121.925 182.970 122.215 183.015 ;
        RECT 123.760 182.970 124.050 183.015 ;
        RECT 118.345 182.830 124.050 182.970 ;
        RECT 118.345 182.785 118.635 182.830 ;
        RECT 121.925 182.785 122.215 182.830 ;
        RECT 123.760 182.785 124.050 182.830 ;
        RECT 105.810 182.430 106.130 182.690 ;
        RECT 109.950 182.430 110.270 182.690 ;
        RECT 110.885 182.445 111.175 182.675 ;
        RECT 120.990 182.630 121.310 182.690 ;
        RECT 124.225 182.630 124.515 182.675 ;
        RECT 124.670 182.630 124.990 182.690 ;
        RECT 120.990 182.490 124.990 182.630 ;
        RECT 105.900 182.290 106.040 182.430 ;
        RECT 110.960 182.290 111.100 182.445 ;
        RECT 120.990 182.430 121.310 182.490 ;
        RECT 124.225 182.445 124.515 182.490 ;
        RECT 124.670 182.430 124.990 182.490 ;
        RECT 105.900 182.150 111.100 182.290 ;
        RECT 112.710 182.290 113.030 182.350 ;
        RECT 115.485 182.290 115.775 182.335 ;
        RECT 112.710 182.150 115.775 182.290 ;
        RECT 112.710 182.090 113.030 182.150 ;
        RECT 115.485 182.105 115.775 182.150 ;
        RECT 118.345 182.290 118.635 182.335 ;
        RECT 121.465 182.290 121.755 182.335 ;
        RECT 123.355 182.290 123.645 182.335 ;
        RECT 118.345 182.150 123.645 182.290 ;
        RECT 118.345 182.105 118.635 182.150 ;
        RECT 121.465 182.105 121.755 182.150 ;
        RECT 123.355 182.105 123.645 182.150 ;
        RECT 106.745 181.950 107.035 181.995 ;
        RECT 109.030 181.950 109.350 182.010 ;
        RECT 104.520 181.810 109.350 181.950 ;
        RECT 94.770 181.750 95.090 181.810 ;
        RECT 102.605 181.765 102.895 181.810 ;
        RECT 106.745 181.765 107.035 181.810 ;
        RECT 109.030 181.750 109.350 181.810 ;
        RECT 114.105 181.950 114.395 181.995 ;
        RECT 119.150 181.950 119.470 182.010 ;
        RECT 114.105 181.810 119.470 181.950 ;
        RECT 114.105 181.765 114.395 181.810 ;
        RECT 119.150 181.750 119.470 181.810 ;
        RECT 37.745 180.930 38.035 180.975 ;
        RECT 40.950 180.930 41.270 180.990 ;
        RECT 37.745 180.790 41.270 180.930 ;
        RECT 37.745 180.745 38.035 180.790 ;
        RECT 40.950 180.730 41.270 180.790 ;
        RECT 49.690 180.730 50.010 180.990 ;
        RECT 54.290 180.930 54.610 180.990 ;
        RECT 55.225 180.930 55.515 180.975 ;
        RECT 73.610 180.930 73.930 180.990 ;
        RECT 54.290 180.790 55.515 180.930 ;
        RECT 54.290 180.730 54.610 180.790 ;
        RECT 55.225 180.745 55.515 180.790 ;
        RECT 70.940 180.790 73.930 180.930 ;
        RECT 25.735 180.590 26.025 180.635 ;
        RECT 27.625 180.590 27.915 180.635 ;
        RECT 30.745 180.590 31.035 180.635 ;
        RECT 25.735 180.450 31.035 180.590 ;
        RECT 25.735 180.405 26.025 180.450 ;
        RECT 27.625 180.405 27.915 180.450 ;
        RECT 30.745 180.405 31.035 180.450 ;
        RECT 49.230 180.590 49.550 180.650 ;
        RECT 58.085 180.590 58.375 180.635 ;
        RECT 61.205 180.590 61.495 180.635 ;
        RECT 63.095 180.590 63.385 180.635 ;
        RECT 49.230 180.450 55.900 180.590 ;
        RECT 49.230 180.390 49.550 180.450 ;
        RECT 33.605 180.250 33.895 180.295 ;
        RECT 34.510 180.250 34.830 180.310 ;
        RECT 33.605 180.110 34.830 180.250 ;
        RECT 33.605 180.065 33.895 180.110 ;
        RECT 34.510 180.050 34.830 180.110 ;
        RECT 52.005 180.250 52.295 180.295 ;
        RECT 52.910 180.250 53.230 180.310 ;
        RECT 52.005 180.110 53.230 180.250 ;
        RECT 55.760 180.250 55.900 180.450 ;
        RECT 58.085 180.450 63.385 180.590 ;
        RECT 58.085 180.405 58.375 180.450 ;
        RECT 61.205 180.405 61.495 180.450 ;
        RECT 63.095 180.405 63.385 180.450 ;
        RECT 66.725 180.590 67.015 180.635 ;
        RECT 68.550 180.590 68.870 180.650 ;
        RECT 70.940 180.590 71.080 180.790 ;
        RECT 73.610 180.730 73.930 180.790 ;
        RECT 83.270 180.730 83.590 180.990 ;
        RECT 87.410 180.930 87.730 180.990 ;
        RECT 90.185 180.930 90.475 180.975 ;
        RECT 87.410 180.790 90.475 180.930 ;
        RECT 87.410 180.730 87.730 180.790 ;
        RECT 90.185 180.745 90.475 180.790 ;
        RECT 97.545 180.930 97.835 180.975 ;
        RECT 99.370 180.930 99.690 180.990 ;
        RECT 97.545 180.790 99.690 180.930 ;
        RECT 97.545 180.745 97.835 180.790 ;
        RECT 99.370 180.730 99.690 180.790 ;
        RECT 99.830 180.930 100.150 180.990 ;
        RECT 102.145 180.930 102.435 180.975 ;
        RECT 99.830 180.790 102.435 180.930 ;
        RECT 99.830 180.730 100.150 180.790 ;
        RECT 102.145 180.745 102.435 180.790 ;
        RECT 123.305 180.930 123.595 180.975 ;
        RECT 124.210 180.930 124.530 180.990 ;
        RECT 123.305 180.790 124.530 180.930 ;
        RECT 123.305 180.745 123.595 180.790 ;
        RECT 124.210 180.730 124.530 180.790 ;
        RECT 74.990 180.590 75.310 180.650 ;
        RECT 75.910 180.590 76.230 180.650 ;
        RECT 85.570 180.590 85.890 180.650 ;
        RECT 66.725 180.450 68.870 180.590 ;
        RECT 66.725 180.405 67.015 180.450 ;
        RECT 66.800 180.250 66.940 180.405 ;
        RECT 68.550 180.390 68.870 180.450 ;
        RECT 69.100 180.450 71.080 180.590 ;
        RECT 72.320 180.450 73.840 180.590 ;
        RECT 69.100 180.295 69.240 180.450 ;
        RECT 72.320 180.310 72.460 180.450 ;
        RECT 55.760 180.110 66.940 180.250 ;
        RECT 52.005 180.065 52.295 180.110 ;
        RECT 52.910 180.050 53.230 180.110 ;
        RECT 69.025 180.065 69.315 180.295 ;
        RECT 69.470 180.050 69.790 180.310 ;
        RECT 70.405 180.250 70.695 180.295 ;
        RECT 72.230 180.250 72.550 180.310 ;
        RECT 70.405 180.110 72.550 180.250 ;
        RECT 70.405 180.065 70.695 180.110 ;
        RECT 72.230 180.050 72.550 180.110 ;
        RECT 72.705 180.250 72.995 180.295 ;
        RECT 73.150 180.250 73.470 180.310 ;
        RECT 72.705 180.110 73.470 180.250 ;
        RECT 73.700 180.250 73.840 180.450 ;
        RECT 74.990 180.450 78.900 180.590 ;
        RECT 74.990 180.390 75.310 180.450 ;
        RECT 75.910 180.390 76.230 180.450 ;
        RECT 76.830 180.250 77.150 180.310 ;
        RECT 78.760 180.295 78.900 180.450 ;
        RECT 80.600 180.450 85.890 180.590 ;
        RECT 80.600 180.295 80.740 180.450 ;
        RECT 85.570 180.390 85.890 180.450 ;
        RECT 105.810 180.590 106.130 180.650 ;
        RECT 105.810 180.450 108.340 180.590 ;
        RECT 105.810 180.390 106.130 180.450 ;
        RECT 73.700 180.110 77.150 180.250 ;
        RECT 72.705 180.065 72.995 180.110 ;
        RECT 73.150 180.050 73.470 180.110 ;
        RECT 76.830 180.050 77.150 180.110 ;
        RECT 77.305 180.065 77.595 180.295 ;
        RECT 78.685 180.065 78.975 180.295 ;
        RECT 80.525 180.065 80.815 180.295 ;
        RECT 24.865 179.725 25.155 179.955 ;
        RECT 25.330 179.910 25.620 179.955 ;
        RECT 27.165 179.910 27.455 179.955 ;
        RECT 30.745 179.910 31.035 179.955 ;
        RECT 25.330 179.770 31.035 179.910 ;
        RECT 25.330 179.725 25.620 179.770 ;
        RECT 27.165 179.725 27.455 179.770 ;
        RECT 30.745 179.725 31.035 179.770 ;
        RECT 24.940 179.230 25.080 179.725 ;
        RECT 26.230 179.370 26.550 179.630 ;
        RECT 27.610 179.570 27.930 179.630 ;
        RECT 31.825 179.615 32.115 179.930 ;
        RECT 34.985 179.910 35.275 179.955 ;
        RECT 36.350 179.910 36.670 179.970 ;
        RECT 34.985 179.770 36.670 179.910 ;
        RECT 34.985 179.725 35.275 179.770 ;
        RECT 36.350 179.710 36.670 179.770 ;
        RECT 39.110 179.910 39.430 179.970 ;
        RECT 39.585 179.910 39.875 179.955 ;
        RECT 39.110 179.770 39.875 179.910 ;
        RECT 39.110 179.710 39.430 179.770 ;
        RECT 39.585 179.725 39.875 179.770 ;
        RECT 43.710 179.910 44.030 179.970 ;
        RECT 46.485 179.910 46.775 179.955 ;
        RECT 54.290 179.910 54.610 179.970 ;
        RECT 43.710 179.770 54.610 179.910 ;
        RECT 43.710 179.710 44.030 179.770 ;
        RECT 46.485 179.725 46.775 179.770 ;
        RECT 54.290 179.710 54.610 179.770 ;
        RECT 28.525 179.570 29.175 179.615 ;
        RECT 31.825 179.570 32.415 179.615 ;
        RECT 27.610 179.430 32.415 179.570 ;
        RECT 27.610 179.370 27.930 179.430 ;
        RECT 28.525 179.385 29.175 179.430 ;
        RECT 32.125 179.385 32.415 179.430 ;
        RECT 37.270 179.570 37.590 179.630 ;
        RECT 45.550 179.570 45.870 179.630 ;
        RECT 55.670 179.570 55.990 179.630 ;
        RECT 57.005 179.615 57.295 179.930 ;
        RECT 58.085 179.910 58.375 179.955 ;
        RECT 61.665 179.910 61.955 179.955 ;
        RECT 63.500 179.910 63.790 179.955 ;
        RECT 58.085 179.770 63.790 179.910 ;
        RECT 58.085 179.725 58.375 179.770 ;
        RECT 61.665 179.725 61.955 179.770 ;
        RECT 63.500 179.725 63.790 179.770 ;
        RECT 63.950 179.710 64.270 179.970 ;
        RECT 65.790 179.710 66.110 179.970 ;
        RECT 67.645 179.910 67.935 179.955 ;
        RECT 66.800 179.770 67.935 179.910 ;
        RECT 56.705 179.570 57.295 179.615 ;
        RECT 59.945 179.570 60.595 179.615 ;
        RECT 37.270 179.430 55.440 179.570 ;
        RECT 37.270 179.370 37.590 179.430 ;
        RECT 45.550 179.370 45.870 179.430 ;
        RECT 25.770 179.230 26.090 179.290 ;
        RECT 37.730 179.230 38.050 179.290 ;
        RECT 24.940 179.090 38.050 179.230 ;
        RECT 25.770 179.030 26.090 179.090 ;
        RECT 37.730 179.030 38.050 179.090 ;
        RECT 38.650 179.030 38.970 179.290 ;
        RECT 54.750 179.030 55.070 179.290 ;
        RECT 55.300 179.230 55.440 179.430 ;
        RECT 55.670 179.430 60.595 179.570 ;
        RECT 55.670 179.370 55.990 179.430 ;
        RECT 56.705 179.385 56.995 179.430 ;
        RECT 59.945 179.385 60.595 179.430 ;
        RECT 61.190 179.570 61.510 179.630 ;
        RECT 62.585 179.570 62.875 179.615 ;
        RECT 66.250 179.570 66.570 179.630 ;
        RECT 61.190 179.430 62.875 179.570 ;
        RECT 61.190 179.370 61.510 179.430 ;
        RECT 62.585 179.385 62.875 179.430 ;
        RECT 63.120 179.430 66.570 179.570 ;
        RECT 63.120 179.230 63.260 179.430 ;
        RECT 66.250 179.370 66.570 179.430 ;
        RECT 55.300 179.090 63.260 179.230 ;
        RECT 65.330 179.030 65.650 179.290 ;
        RECT 66.800 179.230 66.940 179.770 ;
        RECT 67.645 179.725 67.935 179.770 ;
        RECT 68.105 179.910 68.395 179.955 ;
        RECT 68.550 179.910 68.870 179.970 ;
        RECT 68.105 179.770 68.870 179.910 ;
        RECT 68.105 179.725 68.395 179.770 ;
        RECT 68.550 179.710 68.870 179.770 ;
        RECT 69.930 179.710 70.250 179.970 ;
        RECT 74.530 179.910 74.850 179.970 ;
        RECT 77.380 179.910 77.520 180.065 ;
        RECT 80.970 180.050 81.290 180.310 ;
        RECT 94.770 180.050 95.090 180.310 ;
        RECT 98.450 180.050 98.770 180.310 ;
        RECT 108.200 180.295 108.340 180.450 ;
        RECT 111.345 180.405 111.635 180.635 ;
        RECT 114.665 180.590 114.955 180.635 ;
        RECT 117.785 180.590 118.075 180.635 ;
        RECT 119.675 180.590 119.965 180.635 ;
        RECT 114.665 180.450 119.965 180.590 ;
        RECT 114.665 180.405 114.955 180.450 ;
        RECT 117.785 180.405 118.075 180.450 ;
        RECT 119.675 180.405 119.965 180.450 ;
        RECT 120.160 180.450 122.140 180.590 ;
        RECT 100.840 180.110 106.040 180.250 ;
        RECT 100.840 179.970 100.980 180.110 ;
        RECT 105.900 179.970 106.040 180.110 ;
        RECT 108.125 180.065 108.415 180.295 ;
        RECT 109.030 180.050 109.350 180.310 ;
        RECT 111.420 180.250 111.560 180.405 ;
        RECT 120.160 180.250 120.300 180.450 ;
        RECT 111.420 180.110 120.300 180.250 ;
        RECT 120.545 180.250 120.835 180.295 ;
        RECT 120.990 180.250 121.310 180.310 ;
        RECT 120.545 180.110 121.310 180.250 ;
        RECT 120.545 180.065 120.835 180.110 ;
        RECT 120.990 180.050 121.310 180.110 ;
        RECT 70.940 179.770 74.850 179.910 ;
        RECT 70.940 179.630 71.080 179.770 ;
        RECT 74.530 179.710 74.850 179.770 ;
        RECT 75.080 179.770 77.520 179.910 ;
        RECT 70.850 179.370 71.170 179.630 ;
        RECT 71.325 179.570 71.615 179.615 ;
        RECT 71.770 179.570 72.090 179.630 ;
        RECT 71.325 179.430 72.090 179.570 ;
        RECT 71.325 179.385 71.615 179.430 ;
        RECT 71.770 179.370 72.090 179.430 ;
        RECT 73.610 179.570 73.930 179.630 ;
        RECT 75.080 179.615 75.220 179.770 ;
        RECT 77.765 179.725 78.055 179.955 ;
        RECT 78.225 179.725 78.515 179.955 ;
        RECT 95.690 179.910 96.010 179.970 ;
        RECT 100.750 179.910 101.070 179.970 ;
        RECT 95.690 179.770 101.070 179.910 ;
        RECT 75.005 179.570 75.295 179.615 ;
        RECT 73.610 179.430 75.295 179.570 ;
        RECT 73.610 179.370 73.930 179.430 ;
        RECT 75.005 179.385 75.295 179.430 ;
        RECT 76.385 179.385 76.675 179.615 ;
        RECT 77.290 179.570 77.610 179.630 ;
        RECT 77.840 179.570 77.980 179.725 ;
        RECT 77.290 179.430 77.980 179.570 ;
        RECT 68.090 179.230 68.410 179.290 ;
        RECT 76.460 179.230 76.600 179.385 ;
        RECT 77.290 179.370 77.610 179.430 ;
        RECT 66.800 179.090 76.600 179.230 ;
        RECT 76.830 179.230 77.150 179.290 ;
        RECT 78.300 179.230 78.440 179.725 ;
        RECT 95.690 179.710 96.010 179.770 ;
        RECT 100.750 179.710 101.070 179.770 ;
        RECT 101.225 179.910 101.515 179.955 ;
        RECT 103.065 179.910 103.355 179.955 ;
        RECT 101.225 179.770 103.355 179.910 ;
        RECT 101.225 179.725 101.515 179.770 ;
        RECT 103.065 179.725 103.355 179.770 ;
        RECT 105.365 179.725 105.655 179.955 ;
        RECT 83.730 179.370 84.050 179.630 ;
        RECT 76.830 179.090 78.440 179.230 ;
        RECT 68.090 179.030 68.410 179.090 ;
        RECT 76.830 179.030 77.150 179.090 ;
        RECT 81.430 179.030 81.750 179.290 ;
        RECT 103.050 179.230 103.370 179.290 ;
        RECT 103.985 179.230 104.275 179.275 ;
        RECT 103.050 179.090 104.275 179.230 ;
        RECT 105.440 179.230 105.580 179.725 ;
        RECT 105.810 179.710 106.130 179.970 ;
        RECT 106.285 179.725 106.575 179.955 ;
        RECT 106.360 179.570 106.500 179.725 ;
        RECT 107.190 179.710 107.510 179.970 ;
        RECT 113.630 179.930 113.950 179.970 ;
        RECT 122.000 179.955 122.140 180.450 ;
        RECT 113.585 179.710 113.950 179.930 ;
        RECT 114.665 179.910 114.955 179.955 ;
        RECT 118.245 179.910 118.535 179.955 ;
        RECT 120.080 179.910 120.370 179.955 ;
        RECT 114.665 179.770 120.370 179.910 ;
        RECT 114.665 179.725 114.955 179.770 ;
        RECT 118.245 179.725 118.535 179.770 ;
        RECT 120.080 179.725 120.370 179.770 ;
        RECT 121.925 179.725 122.215 179.955 ;
        RECT 122.385 179.725 122.675 179.955 ;
        RECT 109.950 179.570 110.270 179.630 ;
        RECT 113.585 179.615 113.875 179.710 ;
        RECT 113.285 179.570 113.875 179.615 ;
        RECT 116.525 179.570 117.175 179.615 ;
        RECT 106.360 179.430 112.020 179.570 ;
        RECT 109.950 179.370 110.270 179.430 ;
        RECT 106.730 179.230 107.050 179.290 ;
        RECT 105.440 179.090 107.050 179.230 ;
        RECT 103.050 179.030 103.370 179.090 ;
        RECT 103.985 179.045 104.275 179.090 ;
        RECT 106.730 179.030 107.050 179.090 ;
        RECT 109.030 179.230 109.350 179.290 ;
        RECT 111.880 179.275 112.020 179.430 ;
        RECT 113.285 179.430 117.175 179.570 ;
        RECT 113.285 179.385 113.575 179.430 ;
        RECT 116.525 179.385 117.175 179.430 ;
        RECT 119.165 179.385 119.455 179.615 ;
        RECT 119.610 179.570 119.930 179.630 ;
        RECT 122.460 179.570 122.600 179.725 ;
        RECT 119.610 179.430 122.600 179.570 ;
        RECT 109.505 179.230 109.795 179.275 ;
        RECT 109.030 179.090 109.795 179.230 ;
        RECT 109.030 179.030 109.350 179.090 ;
        RECT 109.505 179.045 109.795 179.090 ;
        RECT 111.805 179.045 112.095 179.275 ;
        RECT 119.240 179.230 119.380 179.385 ;
        RECT 119.610 179.370 119.930 179.430 ;
        RECT 121.005 179.230 121.295 179.275 ;
        RECT 119.240 179.090 121.295 179.230 ;
        RECT 121.005 179.045 121.295 179.090 ;
        RECT 26.230 178.210 26.550 178.270 ;
        RECT 26.705 178.210 26.995 178.255 ;
        RECT 26.230 178.070 26.995 178.210 ;
        RECT 26.230 178.010 26.550 178.070 ;
        RECT 26.705 178.025 26.995 178.070 ;
        RECT 27.610 178.010 27.930 178.270 ;
        RECT 37.745 178.210 38.035 178.255 ;
        RECT 39.110 178.210 39.430 178.270 ;
        RECT 37.745 178.070 39.430 178.210 ;
        RECT 37.745 178.025 38.035 178.070 ;
        RECT 39.110 178.010 39.430 178.070 ;
        RECT 39.570 178.010 39.890 178.270 ;
        RECT 49.230 178.210 49.550 178.270 ;
        RECT 52.910 178.210 53.230 178.270 ;
        RECT 49.230 178.070 53.230 178.210 ;
        RECT 49.230 178.010 49.550 178.070 ;
        RECT 52.910 178.010 53.230 178.070 ;
        RECT 54.290 178.210 54.610 178.270 ;
        RECT 57.065 178.210 57.355 178.255 ;
        RECT 54.290 178.070 57.355 178.210 ;
        RECT 54.290 178.010 54.610 178.070 ;
        RECT 57.065 178.025 57.355 178.070 ;
        RECT 62.200 178.070 70.620 178.210 ;
        RECT 25.785 177.870 26.075 177.915 ;
        RECT 27.700 177.870 27.840 178.010 ;
        RECT 25.785 177.730 27.840 177.870 ;
        RECT 29.565 177.870 29.855 177.915 ;
        RECT 32.805 177.870 33.455 177.915 ;
        RECT 29.565 177.730 33.455 177.870 ;
        RECT 25.785 177.685 26.075 177.730 ;
        RECT 29.565 177.685 30.155 177.730 ;
        RECT 32.805 177.685 33.455 177.730 ;
        RECT 35.445 177.870 35.735 177.915 ;
        RECT 38.650 177.870 38.970 177.930 ;
        RECT 35.445 177.730 38.970 177.870 ;
        RECT 35.445 177.685 35.735 177.730 ;
        RECT 29.865 177.590 30.155 177.685 ;
        RECT 38.650 177.670 38.970 177.730 ;
        RECT 40.030 177.870 40.350 177.930 ;
        RECT 48.310 177.870 48.630 177.930 ;
        RECT 62.200 177.915 62.340 178.070 ;
        RECT 70.480 177.915 70.620 178.070 ;
        RECT 71.310 178.010 71.630 178.270 ;
        RECT 72.230 178.210 72.550 178.270 ;
        RECT 74.070 178.210 74.390 178.270 ;
        RECT 95.690 178.210 96.010 178.270 ;
        RECT 72.230 178.070 72.920 178.210 ;
        RECT 72.230 178.010 72.550 178.070 ;
        RECT 40.030 177.730 44.860 177.870 ;
        RECT 40.030 177.670 40.350 177.730 ;
        RECT 26.230 177.330 26.550 177.590 ;
        RECT 27.625 177.530 27.915 177.575 ;
        RECT 28.070 177.530 28.390 177.590 ;
        RECT 27.625 177.390 28.390 177.530 ;
        RECT 27.625 177.345 27.915 177.390 ;
        RECT 28.070 177.330 28.390 177.390 ;
        RECT 29.865 177.370 30.230 177.590 ;
        RECT 29.910 177.330 30.230 177.370 ;
        RECT 30.945 177.530 31.235 177.575 ;
        RECT 34.525 177.530 34.815 177.575 ;
        RECT 36.360 177.530 36.650 177.575 ;
        RECT 30.945 177.390 36.650 177.530 ;
        RECT 30.945 177.345 31.235 177.390 ;
        RECT 34.525 177.345 34.815 177.390 ;
        RECT 36.360 177.345 36.650 177.390 ;
        RECT 36.825 177.530 37.115 177.575 ;
        RECT 37.730 177.530 38.050 177.590 ;
        RECT 36.825 177.390 38.050 177.530 ;
        RECT 36.825 177.345 37.115 177.390 ;
        RECT 37.730 177.330 38.050 177.390 ;
        RECT 43.250 177.530 43.570 177.590 ;
        RECT 44.720 177.575 44.860 177.730 ;
        RECT 48.310 177.730 56.820 177.870 ;
        RECT 48.310 177.670 48.630 177.730 ;
        RECT 43.725 177.530 44.015 177.575 ;
        RECT 43.250 177.390 44.015 177.530 ;
        RECT 43.250 177.330 43.570 177.390 ;
        RECT 43.725 177.345 44.015 177.390 ;
        RECT 44.645 177.345 44.935 177.575 ;
        RECT 45.105 177.345 45.395 177.575 ;
        RECT 34.970 177.190 35.290 177.250 ;
        RECT 40.045 177.190 40.335 177.235 ;
        RECT 34.970 177.050 40.335 177.190 ;
        RECT 34.970 176.990 35.290 177.050 ;
        RECT 40.045 177.005 40.335 177.050 ;
        RECT 40.505 177.005 40.795 177.235 ;
        RECT 30.945 176.850 31.235 176.895 ;
        RECT 34.065 176.850 34.355 176.895 ;
        RECT 35.955 176.850 36.245 176.895 ;
        RECT 40.580 176.850 40.720 177.005 ;
        RECT 30.945 176.710 36.245 176.850 ;
        RECT 30.945 176.665 31.235 176.710 ;
        RECT 34.065 176.665 34.355 176.710 ;
        RECT 35.955 176.665 36.245 176.710 ;
        RECT 39.660 176.710 40.720 176.850 ;
        RECT 45.180 176.850 45.320 177.345 ;
        RECT 45.550 177.330 45.870 177.590 ;
        RECT 49.230 177.330 49.550 177.590 ;
        RECT 49.780 177.575 49.920 177.730 ;
        RECT 49.705 177.345 49.995 177.575 ;
        RECT 50.165 177.530 50.455 177.575 ;
        RECT 50.610 177.530 50.930 177.590 ;
        RECT 50.165 177.390 50.930 177.530 ;
        RECT 50.165 177.345 50.455 177.390 ;
        RECT 50.610 177.330 50.930 177.390 ;
        RECT 51.085 177.345 51.375 177.575 ;
        RECT 51.160 177.190 51.300 177.345 ;
        RECT 52.910 177.330 53.230 177.590 ;
        RECT 53.460 177.575 53.600 177.730 ;
        RECT 53.385 177.345 53.675 177.575 ;
        RECT 53.830 177.330 54.150 177.590 ;
        RECT 54.765 177.530 55.055 177.575 ;
        RECT 55.210 177.530 55.530 177.590 ;
        RECT 54.765 177.390 55.530 177.530 ;
        RECT 54.765 177.345 55.055 177.390 ;
        RECT 54.840 177.190 54.980 177.345 ;
        RECT 55.210 177.330 55.530 177.390 ;
        RECT 51.160 177.050 54.980 177.190 ;
        RECT 56.130 176.990 56.450 177.250 ;
        RECT 56.680 177.190 56.820 177.730 ;
        RECT 62.125 177.685 62.415 177.915 ;
        RECT 70.405 177.870 70.695 177.915 ;
        RECT 70.850 177.870 71.170 177.930 ;
        RECT 70.405 177.730 71.170 177.870 ;
        RECT 71.400 177.870 71.540 178.010 ;
        RECT 71.400 177.730 72.000 177.870 ;
        RECT 70.405 177.685 70.695 177.730 ;
        RECT 70.850 177.670 71.170 177.730 ;
        RECT 57.525 177.530 57.815 177.575 ;
        RECT 57.970 177.530 58.290 177.590 ;
        RECT 57.525 177.390 58.290 177.530 ;
        RECT 57.525 177.345 57.815 177.390 ;
        RECT 57.970 177.330 58.290 177.390 ;
        RECT 65.345 177.345 65.635 177.575 ;
        RECT 67.185 177.530 67.475 177.575 ;
        RECT 68.090 177.530 68.410 177.590 ;
        RECT 67.185 177.390 68.410 177.530 ;
        RECT 67.185 177.345 67.475 177.390 ;
        RECT 65.420 177.190 65.560 177.345 ;
        RECT 68.090 177.330 68.410 177.390 ;
        RECT 69.010 177.545 69.330 177.590 ;
        RECT 69.945 177.545 70.235 177.575 ;
        RECT 69.010 177.530 70.235 177.545 ;
        RECT 71.310 177.530 71.630 177.590 ;
        RECT 71.860 177.575 72.000 177.730 ;
        RECT 69.010 177.405 71.630 177.530 ;
        RECT 69.010 177.330 69.330 177.405 ;
        RECT 69.945 177.390 71.630 177.405 ;
        RECT 69.945 177.345 70.235 177.390 ;
        RECT 71.310 177.330 71.630 177.390 ;
        RECT 71.785 177.345 72.075 177.575 ;
        RECT 72.230 177.330 72.550 177.590 ;
        RECT 72.780 177.575 72.920 178.070 ;
        RECT 74.070 178.070 96.010 178.210 ;
        RECT 74.070 178.010 74.390 178.070 ;
        RECT 95.690 178.010 96.010 178.070 ;
        RECT 96.150 178.010 96.470 178.270 ;
        RECT 101.670 178.210 101.990 178.270 ;
        RECT 107.190 178.210 107.510 178.270 ;
        RECT 101.670 178.070 108.800 178.210 ;
        RECT 101.670 178.010 101.990 178.070 ;
        RECT 107.190 178.010 107.510 178.070 ;
        RECT 73.610 177.870 73.930 177.930 ;
        RECT 86.490 177.870 86.810 177.930 ;
        RECT 73.240 177.730 73.930 177.870 ;
        RECT 73.240 177.575 73.380 177.730 ;
        RECT 73.610 177.670 73.930 177.730 ;
        RECT 75.080 177.730 86.810 177.870 ;
        RECT 75.080 177.575 75.220 177.730 ;
        RECT 86.490 177.670 86.810 177.730 ;
        RECT 72.705 177.345 72.995 177.575 ;
        RECT 73.165 177.345 73.455 177.575 ;
        RECT 74.085 177.345 74.375 177.575 ;
        RECT 75.005 177.345 75.295 177.575 ;
        RECT 56.680 177.050 64.640 177.190 ;
        RECT 65.420 177.050 68.780 177.190 ;
        RECT 57.050 176.850 57.370 176.910 ;
        RECT 59.365 176.850 59.655 176.895 ;
        RECT 45.180 176.710 52.220 176.850 ;
        RECT 27.610 176.510 27.930 176.570 ;
        RECT 28.085 176.510 28.375 176.555 ;
        RECT 27.610 176.370 28.375 176.510 ;
        RECT 27.610 176.310 27.930 176.370 ;
        RECT 28.085 176.325 28.375 176.370 ;
        RECT 35.430 176.510 35.750 176.570 ;
        RECT 39.660 176.510 39.800 176.710 ;
        RECT 35.430 176.370 39.800 176.510 ;
        RECT 40.030 176.510 40.350 176.570 ;
        RECT 45.180 176.510 45.320 176.710 ;
        RECT 40.030 176.370 45.320 176.510 ;
        RECT 46.945 176.510 47.235 176.555 ;
        RECT 47.390 176.510 47.710 176.570 ;
        RECT 46.945 176.370 47.710 176.510 ;
        RECT 35.430 176.310 35.750 176.370 ;
        RECT 40.030 176.310 40.350 176.370 ;
        RECT 46.945 176.325 47.235 176.370 ;
        RECT 47.390 176.310 47.710 176.370 ;
        RECT 47.850 176.310 48.170 176.570 ;
        RECT 49.690 176.510 50.010 176.570 ;
        RECT 51.545 176.510 51.835 176.555 ;
        RECT 49.690 176.370 51.835 176.510 ;
        RECT 52.080 176.510 52.220 176.710 ;
        RECT 57.050 176.710 59.655 176.850 ;
        RECT 57.050 176.650 57.370 176.710 ;
        RECT 59.365 176.665 59.655 176.710 ;
        RECT 64.500 176.570 64.640 177.050 ;
        RECT 66.250 176.650 66.570 176.910 ;
        RECT 57.510 176.510 57.830 176.570 ;
        RECT 52.080 176.370 57.830 176.510 ;
        RECT 49.690 176.310 50.010 176.370 ;
        RECT 51.545 176.325 51.835 176.370 ;
        RECT 57.510 176.310 57.830 176.370 ;
        RECT 59.810 176.510 60.130 176.570 ;
        RECT 60.745 176.510 61.035 176.555 ;
        RECT 59.810 176.370 61.035 176.510 ;
        RECT 59.810 176.310 60.130 176.370 ;
        RECT 60.745 176.325 61.035 176.370 ;
        RECT 64.410 176.310 64.730 176.570 ;
        RECT 68.640 176.555 68.780 177.050 ;
        RECT 69.485 177.005 69.775 177.235 ;
        RECT 70.865 177.190 71.155 177.235 ;
        RECT 73.610 177.190 73.930 177.250 ;
        RECT 74.160 177.190 74.300 177.345 ;
        RECT 75.450 177.330 75.770 177.590 ;
        RECT 75.910 177.530 76.230 177.590 ;
        RECT 77.750 177.530 78.070 177.590 ;
        RECT 75.910 177.390 78.070 177.530 ;
        RECT 75.910 177.330 76.230 177.390 ;
        RECT 77.750 177.330 78.070 177.390 ;
        RECT 87.410 177.330 87.730 177.590 ;
        RECT 96.625 177.530 96.915 177.575 ;
        RECT 97.070 177.530 97.390 177.590 ;
        RECT 100.075 177.530 100.365 177.575 ;
        RECT 100.750 177.545 101.070 177.590 ;
        RECT 96.625 177.390 97.390 177.530 ;
        RECT 96.625 177.345 96.915 177.390 ;
        RECT 97.070 177.330 97.390 177.390 ;
        RECT 99.460 177.390 100.365 177.530 ;
        RECT 100.570 177.405 101.070 177.545 ;
        RECT 76.370 177.190 76.690 177.250 ;
        RECT 77.290 177.190 77.610 177.250 ;
        RECT 70.865 177.050 73.380 177.190 ;
        RECT 70.865 177.005 71.155 177.050 ;
        RECT 69.010 176.850 69.330 176.910 ;
        RECT 69.560 176.850 69.700 177.005 ;
        RECT 69.010 176.710 69.700 176.850 ;
        RECT 69.010 176.650 69.330 176.710 ;
        RECT 68.565 176.510 68.855 176.555 ;
        RECT 70.940 176.510 71.080 177.005 ;
        RECT 73.240 176.910 73.380 177.050 ;
        RECT 73.610 177.050 77.610 177.190 ;
        RECT 73.610 176.990 73.930 177.050 ;
        RECT 76.370 176.990 76.690 177.050 ;
        RECT 77.290 176.990 77.610 177.050 ;
        RECT 73.150 176.650 73.470 176.910 ;
        RECT 74.530 176.850 74.850 176.910 ;
        RECT 99.460 176.850 99.600 177.390 ;
        RECT 100.075 177.345 100.365 177.390 ;
        RECT 100.750 177.330 101.070 177.405 ;
        RECT 101.210 177.345 101.530 177.605 ;
        RECT 108.660 177.590 108.800 178.070 ;
        RECT 109.030 178.010 109.350 178.270 ;
        RECT 113.630 178.010 113.950 178.270 ;
        RECT 117.310 178.010 117.630 178.270 ;
        RECT 101.670 177.530 101.990 177.590 ;
        RECT 102.145 177.530 102.435 177.575 ;
        RECT 101.670 177.390 102.435 177.530 ;
        RECT 101.670 177.330 101.990 177.390 ;
        RECT 102.145 177.345 102.435 177.390 ;
        RECT 106.730 177.330 107.050 177.590 ;
        RECT 107.205 177.345 107.495 177.575 ;
        RECT 105.810 177.190 106.130 177.250 ;
        RECT 107.280 177.190 107.420 177.345 ;
        RECT 107.650 177.330 107.970 177.590 ;
        RECT 108.570 177.330 108.890 177.590 ;
        RECT 112.265 177.530 112.555 177.575 ;
        RECT 112.710 177.530 113.030 177.590 ;
        RECT 112.265 177.390 113.030 177.530 ;
        RECT 112.265 177.345 112.555 177.390 ;
        RECT 112.710 177.330 113.030 177.390 ;
        RECT 113.185 177.530 113.475 177.575 ;
        RECT 115.930 177.530 116.250 177.590 ;
        RECT 116.865 177.530 117.155 177.575 ;
        RECT 113.185 177.390 117.155 177.530 ;
        RECT 113.185 177.345 113.475 177.390 ;
        RECT 115.930 177.330 116.250 177.390 ;
        RECT 116.865 177.345 117.155 177.390 ;
        RECT 109.950 177.190 110.270 177.250 ;
        RECT 105.810 177.050 110.270 177.190 ;
        RECT 112.800 177.190 112.940 177.330 ;
        RECT 115.470 177.190 115.790 177.250 ;
        RECT 112.800 177.050 115.790 177.190 ;
        RECT 105.810 176.990 106.130 177.050 ;
        RECT 109.950 176.990 110.270 177.050 ;
        RECT 115.470 176.990 115.790 177.050 ;
        RECT 106.730 176.850 107.050 176.910 ;
        RECT 109.490 176.850 109.810 176.910 ;
        RECT 74.530 176.710 109.810 176.850 ;
        RECT 74.530 176.650 74.850 176.710 ;
        RECT 106.730 176.650 107.050 176.710 ;
        RECT 109.490 176.650 109.810 176.710 ;
        RECT 68.565 176.370 71.080 176.510 ;
        RECT 68.565 176.325 68.855 176.370 ;
        RECT 77.290 176.310 77.610 176.570 ;
        RECT 77.750 176.510 78.070 176.570 ;
        RECT 84.190 176.510 84.510 176.570 ;
        RECT 77.750 176.370 84.510 176.510 ;
        RECT 77.750 176.310 78.070 176.370 ;
        RECT 84.190 176.310 84.510 176.370 ;
        RECT 98.925 176.510 99.215 176.555 ;
        RECT 99.830 176.510 100.150 176.570 ;
        RECT 98.925 176.370 100.150 176.510 ;
        RECT 98.925 176.325 99.215 176.370 ;
        RECT 99.830 176.310 100.150 176.370 ;
        RECT 104.890 176.510 105.210 176.570 ;
        RECT 105.365 176.510 105.655 176.555 ;
        RECT 104.890 176.370 105.655 176.510 ;
        RECT 104.890 176.310 105.210 176.370 ;
        RECT 105.365 176.325 105.655 176.370 ;
        RECT 110.870 176.510 111.190 176.570 ;
        RECT 113.630 176.510 113.950 176.570 ;
        RECT 110.870 176.370 113.950 176.510 ;
        RECT 110.870 176.310 111.190 176.370 ;
        RECT 113.630 176.310 113.950 176.370 ;
        RECT 26.245 175.490 26.535 175.535 ;
        RECT 29.910 175.490 30.230 175.550 ;
        RECT 26.245 175.350 30.230 175.490 ;
        RECT 26.245 175.305 26.535 175.350 ;
        RECT 29.910 175.290 30.230 175.350 ;
        RECT 55.210 175.490 55.530 175.550 ;
        RECT 71.785 175.490 72.075 175.535 ;
        RECT 73.610 175.490 73.930 175.550 ;
        RECT 55.210 175.350 73.930 175.490 ;
        RECT 55.210 175.290 55.530 175.350 ;
        RECT 71.785 175.305 72.075 175.350 ;
        RECT 73.610 175.290 73.930 175.350 ;
        RECT 74.070 175.290 74.390 175.550 ;
        RECT 75.450 175.490 75.770 175.550 ;
        RECT 78.670 175.490 78.990 175.550 ;
        RECT 75.450 175.350 78.990 175.490 ;
        RECT 75.450 175.290 75.770 175.350 ;
        RECT 78.670 175.290 78.990 175.350 ;
        RECT 81.430 175.490 81.750 175.550 ;
        RECT 84.665 175.490 84.955 175.535 ;
        RECT 81.430 175.350 84.955 175.490 ;
        RECT 81.430 175.290 81.750 175.350 ;
        RECT 84.665 175.305 84.955 175.350 ;
        RECT 85.570 175.490 85.890 175.550 ;
        RECT 89.265 175.490 89.555 175.535 ;
        RECT 85.570 175.350 89.555 175.490 ;
        RECT 85.570 175.290 85.890 175.350 ;
        RECT 89.265 175.305 89.555 175.350 ;
        RECT 112.250 175.490 112.570 175.550 ;
        RECT 118.245 175.490 118.535 175.535 ;
        RECT 112.250 175.350 118.535 175.490 ;
        RECT 112.250 175.290 112.570 175.350 ;
        RECT 118.245 175.305 118.535 175.350 ;
        RECT 28.070 175.150 28.390 175.210 ;
        RECT 31.305 175.150 31.595 175.195 ;
        RECT 35.430 175.150 35.750 175.210 ;
        RECT 28.070 175.010 31.595 175.150 ;
        RECT 28.070 174.950 28.390 175.010 ;
        RECT 31.305 174.965 31.595 175.010 ;
        RECT 34.600 175.010 35.750 175.150 ;
        RECT 33.605 174.810 33.895 174.855 ;
        RECT 34.050 174.810 34.370 174.870 ;
        RECT 34.600 174.855 34.740 175.010 ;
        RECT 35.430 174.950 35.750 175.010 ;
        RECT 38.665 175.150 38.955 175.195 ;
        RECT 40.490 175.150 40.810 175.210 ;
        RECT 44.630 175.150 44.950 175.210 ;
        RECT 49.230 175.150 49.550 175.210 ;
        RECT 38.665 175.010 40.810 175.150 ;
        RECT 38.665 174.965 38.955 175.010 ;
        RECT 40.490 174.950 40.810 175.010 ;
        RECT 41.040 175.010 49.550 175.150 ;
        RECT 33.605 174.670 34.370 174.810 ;
        RECT 33.605 174.625 33.895 174.670 ;
        RECT 34.050 174.610 34.370 174.670 ;
        RECT 34.525 174.625 34.815 174.855 ;
        RECT 40.030 174.810 40.350 174.870 ;
        RECT 41.040 174.810 41.180 175.010 ;
        RECT 44.630 174.950 44.950 175.010 ;
        RECT 43.250 174.810 43.570 174.870 ;
        RECT 36.900 174.670 40.350 174.810 ;
        RECT 26.230 174.470 26.550 174.530 ;
        RECT 26.705 174.470 26.995 174.515 ;
        RECT 26.230 174.330 26.995 174.470 ;
        RECT 26.230 174.270 26.550 174.330 ;
        RECT 26.705 174.285 26.995 174.330 ;
        RECT 26.780 173.790 26.920 174.285 ;
        RECT 27.610 174.270 27.930 174.530 ;
        RECT 30.385 174.470 30.675 174.515 ;
        RECT 33.145 174.470 33.435 174.515 ;
        RECT 34.970 174.470 35.290 174.530 ;
        RECT 30.385 174.330 35.290 174.470 ;
        RECT 30.385 174.285 30.675 174.330 ;
        RECT 33.145 174.285 33.435 174.330 ;
        RECT 34.970 174.270 35.290 174.330 ;
        RECT 35.445 174.470 35.735 174.515 ;
        RECT 35.890 174.470 36.210 174.530 ;
        RECT 36.900 174.515 37.040 174.670 ;
        RECT 40.030 174.610 40.350 174.670 ;
        RECT 40.580 174.670 41.180 174.810 ;
        RECT 42.880 174.670 47.160 174.810 ;
        RECT 35.445 174.330 36.210 174.470 ;
        RECT 35.445 174.285 35.735 174.330 ;
        RECT 35.890 174.270 36.210 174.330 ;
        RECT 36.365 174.285 36.655 174.515 ;
        RECT 36.825 174.285 37.115 174.515 ;
        RECT 27.700 174.130 27.840 174.270 ;
        RECT 36.440 174.130 36.580 174.285 ;
        RECT 37.270 174.270 37.590 174.530 ;
        RECT 40.580 174.515 40.720 174.670 ;
        RECT 40.505 174.285 40.795 174.515 ;
        RECT 40.965 174.285 41.255 174.515 ;
        RECT 41.425 174.470 41.715 174.515 ;
        RECT 41.870 174.470 42.190 174.530 ;
        RECT 42.880 174.515 43.020 174.670 ;
        RECT 43.250 174.610 43.570 174.670 ;
        RECT 41.425 174.330 42.190 174.470 ;
        RECT 41.425 174.285 41.715 174.330 ;
        RECT 27.700 173.990 36.580 174.130 ;
        RECT 38.190 174.130 38.510 174.190 ;
        RECT 39.125 174.130 39.415 174.175 ;
        RECT 38.190 173.990 39.415 174.130 ;
        RECT 41.040 174.130 41.180 174.285 ;
        RECT 41.870 174.270 42.190 174.330 ;
        RECT 42.345 174.470 42.635 174.515 ;
        RECT 42.805 174.470 43.095 174.515 ;
        RECT 42.345 174.330 43.095 174.470 ;
        RECT 42.345 174.285 42.635 174.330 ;
        RECT 42.805 174.285 43.095 174.330 ;
        RECT 43.710 174.270 44.030 174.530 ;
        RECT 44.185 174.285 44.475 174.515 ;
        RECT 44.260 174.130 44.400 174.285 ;
        RECT 44.630 174.270 44.950 174.530 ;
        RECT 41.040 173.990 44.400 174.130 ;
        RECT 38.190 173.930 38.510 173.990 ;
        RECT 39.125 173.945 39.415 173.990 ;
        RECT 31.290 173.790 31.610 173.850 ;
        RECT 26.780 173.650 31.610 173.790 ;
        RECT 44.260 173.790 44.400 173.990 ;
        RECT 46.010 173.930 46.330 174.190 ;
        RECT 46.470 173.930 46.790 174.190 ;
        RECT 47.020 174.130 47.160 174.670 ;
        RECT 47.940 174.515 48.080 175.010 ;
        RECT 49.230 174.950 49.550 175.010 ;
        RECT 55.300 174.810 55.440 175.290 ;
        RECT 60.285 174.965 60.575 175.195 ;
        RECT 64.410 175.150 64.730 175.210 ;
        RECT 69.930 175.150 70.250 175.210 ;
        RECT 75.910 175.150 76.230 175.210 ;
        RECT 64.410 175.010 69.700 175.150 ;
        RECT 48.860 174.670 52.680 174.810 ;
        RECT 47.865 174.285 48.155 174.515 ;
        RECT 48.310 174.270 48.630 174.530 ;
        RECT 48.860 174.515 49.000 174.670 ;
        RECT 52.540 174.530 52.680 174.670 ;
        RECT 53.000 174.670 55.440 174.810 ;
        RECT 56.130 174.810 56.450 174.870 ;
        RECT 57.525 174.810 57.815 174.855 ;
        RECT 59.810 174.810 60.130 174.870 ;
        RECT 56.130 174.670 60.130 174.810 ;
        RECT 48.785 174.285 49.075 174.515 ;
        RECT 49.705 174.285 49.995 174.515 ;
        RECT 49.780 174.130 49.920 174.285 ;
        RECT 52.450 174.270 52.770 174.530 ;
        RECT 53.000 174.130 53.140 174.670 ;
        RECT 56.130 174.610 56.450 174.670 ;
        RECT 57.525 174.625 57.815 174.670 ;
        RECT 59.810 174.610 60.130 174.670 ;
        RECT 55.225 174.470 55.515 174.515 ;
        RECT 57.970 174.470 58.290 174.530 ;
        RECT 55.225 174.330 58.290 174.470 ;
        RECT 60.360 174.470 60.500 174.965 ;
        RECT 64.410 174.950 64.730 175.010 ;
        RECT 66.710 174.810 67.030 174.870 ;
        RECT 69.025 174.810 69.315 174.855 ;
        RECT 66.710 174.670 69.315 174.810 ;
        RECT 69.560 174.810 69.700 175.010 ;
        RECT 69.930 175.010 76.230 175.150 ;
        RECT 78.760 175.150 78.900 175.290 ;
        RECT 82.810 175.150 83.130 175.210 ;
        RECT 78.760 175.010 83.130 175.150 ;
        RECT 69.930 174.950 70.250 175.010 ;
        RECT 75.910 174.950 76.230 175.010 ;
        RECT 82.810 174.950 83.130 175.010 ;
        RECT 109.950 175.150 110.270 175.210 ;
        RECT 109.950 175.010 113.400 175.150 ;
        RECT 109.950 174.950 110.270 175.010 ;
        RECT 70.850 174.810 71.170 174.870 ;
        RECT 87.885 174.810 88.175 174.855 ;
        RECT 90.630 174.810 90.950 174.870 ;
        RECT 69.560 174.670 70.620 174.810 ;
        RECT 66.710 174.610 67.030 174.670 ;
        RECT 69.025 174.625 69.315 174.670 ;
        RECT 63.505 174.470 63.795 174.515 ;
        RECT 60.360 174.330 63.795 174.470 ;
        RECT 55.225 174.285 55.515 174.330 ;
        RECT 57.970 174.270 58.290 174.330 ;
        RECT 63.505 174.285 63.795 174.330 ;
        RECT 68.105 174.480 68.395 174.515 ;
        RECT 68.105 174.470 68.780 174.480 ;
        RECT 68.105 174.340 69.240 174.470 ;
        RECT 68.105 174.285 68.395 174.340 ;
        RECT 68.640 174.330 69.240 174.340 ;
        RECT 69.100 174.190 69.240 174.330 ;
        RECT 47.020 173.990 53.140 174.130 ;
        RECT 54.750 174.130 55.070 174.190 ;
        RECT 58.445 174.130 58.735 174.175 ;
        RECT 54.750 173.990 58.735 174.130 ;
        RECT 54.750 173.930 55.070 173.990 ;
        RECT 58.445 173.945 58.735 173.990 ;
        RECT 69.010 173.930 69.330 174.190 ;
        RECT 70.480 174.130 70.620 174.670 ;
        RECT 70.850 174.670 85.110 174.810 ;
        RECT 70.850 174.610 71.170 174.670 ;
        RECT 71.310 174.470 71.630 174.530 ;
        RECT 72.705 174.470 72.995 174.515 ;
        RECT 71.310 174.330 72.995 174.470 ;
        RECT 71.310 174.270 71.630 174.330 ;
        RECT 72.705 174.285 72.995 174.330 ;
        RECT 73.150 174.270 73.470 174.530 ;
        RECT 77.305 174.470 77.595 174.515 ;
        RECT 77.750 174.470 78.070 174.530 ;
        RECT 77.305 174.330 78.070 174.470 ;
        RECT 77.305 174.285 77.595 174.330 ;
        RECT 77.750 174.270 78.070 174.330 ;
        RECT 78.210 174.270 78.530 174.530 ;
        RECT 78.670 174.270 78.990 174.530 ;
        RECT 79.145 174.470 79.435 174.515 ;
        RECT 82.365 174.470 82.655 174.515 ;
        RECT 79.145 174.330 82.655 174.470 ;
        RECT 79.145 174.285 79.435 174.330 ;
        RECT 82.365 174.285 82.655 174.330 ;
        RECT 75.450 174.130 75.770 174.190 ;
        RECT 70.480 173.990 75.770 174.130 ;
        RECT 75.450 173.930 75.770 173.990 ;
        RECT 75.910 174.130 76.230 174.190 ;
        RECT 79.220 174.130 79.360 174.285 ;
        RECT 82.810 174.270 83.130 174.530 ;
        RECT 83.285 174.285 83.575 174.515 ;
        RECT 75.910 173.990 79.360 174.130 ;
        RECT 80.050 174.130 80.370 174.190 ;
        RECT 80.525 174.130 80.815 174.175 ;
        RECT 80.050 173.990 80.815 174.130 ;
        RECT 75.910 173.930 76.230 173.990 ;
        RECT 80.050 173.930 80.370 173.990 ;
        RECT 80.525 173.945 80.815 173.990 ;
        RECT 80.985 174.130 81.275 174.175 ;
        RECT 81.890 174.130 82.210 174.190 ;
        RECT 80.985 173.990 82.210 174.130 ;
        RECT 83.360 174.130 83.500 174.285 ;
        RECT 84.190 174.270 84.510 174.530 ;
        RECT 84.970 174.470 85.110 174.670 ;
        RECT 87.885 174.670 90.950 174.810 ;
        RECT 87.885 174.625 88.175 174.670 ;
        RECT 88.805 174.470 89.095 174.515 ;
        RECT 84.970 174.330 89.095 174.470 ;
        RECT 88.805 174.285 89.095 174.330 ;
        RECT 89.340 174.130 89.480 174.670 ;
        RECT 90.630 174.610 90.950 174.670 ;
        RECT 106.730 174.810 107.050 174.870 ;
        RECT 111.345 174.810 111.635 174.855 ;
        RECT 113.260 174.810 113.400 175.010 ;
        RECT 106.730 174.670 111.635 174.810 ;
        RECT 106.730 174.610 107.050 174.670 ;
        RECT 111.345 174.625 111.635 174.670 ;
        RECT 111.880 174.670 112.840 174.810 ;
        RECT 102.130 174.270 102.450 174.530 ;
        RECT 83.360 173.990 89.480 174.130 ;
        RECT 110.885 174.130 111.175 174.175 ;
        RECT 111.330 174.130 111.650 174.190 ;
        RECT 110.885 173.990 111.650 174.130 ;
        RECT 111.880 174.130 112.020 174.670 ;
        RECT 112.700 174.515 112.840 174.670 ;
        RECT 113.260 174.670 116.620 174.810 ;
        RECT 113.260 174.515 113.400 174.670 ;
        RECT 112.495 174.330 112.840 174.515 ;
        RECT 112.495 174.285 112.785 174.330 ;
        RECT 113.185 174.285 113.475 174.515 ;
        RECT 113.630 174.270 113.950 174.530 ;
        RECT 114.550 174.470 114.870 174.530 ;
        RECT 115.025 174.470 115.315 174.515 ;
        RECT 114.550 174.330 115.315 174.470 ;
        RECT 114.550 174.270 114.870 174.330 ;
        RECT 115.025 174.285 115.315 174.330 ;
        RECT 115.470 174.470 115.790 174.530 ;
        RECT 116.480 174.515 116.620 174.670 ;
        RECT 115.945 174.470 116.235 174.515 ;
        RECT 115.470 174.330 116.235 174.470 ;
        RECT 115.470 174.270 115.790 174.330 ;
        RECT 115.945 174.285 116.235 174.330 ;
        RECT 116.405 174.285 116.695 174.515 ;
        RECT 116.865 174.285 117.155 174.515 ;
        RECT 119.625 174.285 119.915 174.515 ;
        RECT 116.940 174.130 117.080 174.285 ;
        RECT 111.880 173.990 112.480 174.130 ;
        RECT 80.985 173.945 81.275 173.990 ;
        RECT 81.890 173.930 82.210 173.990 ;
        RECT 110.885 173.945 111.175 173.990 ;
        RECT 111.330 173.930 111.650 173.990 ;
        RECT 48.310 173.790 48.630 173.850 ;
        RECT 44.260 173.650 48.630 173.790 ;
        RECT 31.290 173.590 31.610 173.650 ;
        RECT 48.310 173.590 48.630 173.650 ;
        RECT 61.190 173.790 61.510 173.850 ;
        RECT 62.585 173.790 62.875 173.835 ;
        RECT 61.190 173.650 62.875 173.790 ;
        RECT 61.190 173.590 61.510 173.650 ;
        RECT 62.585 173.605 62.875 173.650 ;
        RECT 78.210 173.790 78.530 173.850 ;
        RECT 101.670 173.790 101.990 173.850 ;
        RECT 78.210 173.650 101.990 173.790 ;
        RECT 78.210 173.590 78.530 173.650 ;
        RECT 101.670 173.590 101.990 173.650 ;
        RECT 109.490 173.790 109.810 173.850 ;
        RECT 112.340 173.790 112.480 173.990 ;
        RECT 113.260 173.990 117.080 174.130 ;
        RECT 117.770 174.130 118.090 174.190 ;
        RECT 119.165 174.130 119.455 174.175 ;
        RECT 117.770 173.990 119.455 174.130 ;
        RECT 113.260 173.790 113.400 173.990 ;
        RECT 117.770 173.930 118.090 173.990 ;
        RECT 119.165 173.945 119.455 173.990 ;
        RECT 109.490 173.650 113.400 173.790 ;
        RECT 117.310 173.790 117.630 173.850 ;
        RECT 119.700 173.790 119.840 174.285 ;
        RECT 117.310 173.650 119.840 173.790 ;
        RECT 109.490 173.590 109.810 173.650 ;
        RECT 117.310 173.590 117.630 173.650 ;
        RECT 52.450 172.770 52.770 172.830 ;
        RECT 53.845 172.770 54.135 172.815 ;
        RECT 63.965 172.770 64.255 172.815 ;
        RECT 97.070 172.770 97.390 172.830 ;
        RECT 108.110 172.770 108.430 172.830 ;
        RECT 112.250 172.770 112.570 172.830 ;
        RECT 52.450 172.630 54.135 172.770 ;
        RECT 52.450 172.570 52.770 172.630 ;
        RECT 53.845 172.585 54.135 172.630 ;
        RECT 60.820 172.630 64.255 172.770 ;
        RECT 35.890 172.430 36.210 172.490 ;
        RECT 55.325 172.430 55.615 172.475 ;
        RECT 58.565 172.430 59.215 172.475 ;
        RECT 60.820 172.430 60.960 172.630 ;
        RECT 63.965 172.585 64.255 172.630 ;
        RECT 89.800 172.630 112.570 172.770 ;
        RECT 33.680 172.290 41.640 172.430 ;
        RECT 33.680 172.135 33.820 172.290 ;
        RECT 35.890 172.230 36.210 172.290 ;
        RECT 41.500 172.150 41.640 172.290 ;
        RECT 55.325 172.290 60.960 172.430 ;
        RECT 55.325 172.245 55.915 172.290 ;
        RECT 58.565 172.245 59.215 172.290 ;
        RECT 33.605 171.905 33.895 172.135 ;
        RECT 34.510 171.890 34.830 172.150 ;
        RECT 34.985 171.905 35.275 172.135 ;
        RECT 35.445 172.090 35.735 172.135 ;
        RECT 37.270 172.090 37.590 172.150 ;
        RECT 39.585 172.090 39.875 172.135 ;
        RECT 35.445 171.950 39.875 172.090 ;
        RECT 35.445 171.905 35.735 171.950 ;
        RECT 35.060 171.750 35.200 171.905 ;
        RECT 37.270 171.890 37.590 171.950 ;
        RECT 39.585 171.905 39.875 171.950 ;
        RECT 40.030 171.890 40.350 172.150 ;
        RECT 40.505 172.090 40.795 172.135 ;
        RECT 40.950 172.090 41.270 172.150 ;
        RECT 40.505 171.950 41.270 172.090 ;
        RECT 40.505 171.905 40.795 171.950 ;
        RECT 40.950 171.890 41.270 171.950 ;
        RECT 41.410 171.890 41.730 172.150 ;
        RECT 53.370 171.890 53.690 172.150 ;
        RECT 55.625 171.930 55.915 172.245 ;
        RECT 61.190 172.230 61.510 172.490 ;
        RECT 83.745 172.430 84.035 172.475 ;
        RECT 89.800 172.430 89.940 172.630 ;
        RECT 97.070 172.570 97.390 172.630 ;
        RECT 108.110 172.570 108.430 172.630 ;
        RECT 112.250 172.570 112.570 172.630 ;
        RECT 83.745 172.290 89.940 172.430 ;
        RECT 83.745 172.245 84.035 172.290 ;
        RECT 56.705 172.090 56.995 172.135 ;
        RECT 60.285 172.090 60.575 172.135 ;
        RECT 62.120 172.090 62.410 172.135 ;
        RECT 56.705 171.950 62.410 172.090 ;
        RECT 56.705 171.905 56.995 171.950 ;
        RECT 60.285 171.905 60.575 171.950 ;
        RECT 62.120 171.905 62.410 171.950 ;
        RECT 64.410 171.890 64.730 172.150 ;
        RECT 69.010 172.090 69.330 172.150 ;
        RECT 89.800 172.135 89.940 172.290 ;
        RECT 90.185 172.430 90.475 172.475 ;
        RECT 92.585 172.430 92.875 172.475 ;
        RECT 95.825 172.430 96.475 172.475 ;
        RECT 90.185 172.290 96.475 172.430 ;
        RECT 90.185 172.245 90.475 172.290 ;
        RECT 92.585 172.245 93.175 172.290 ;
        RECT 95.825 172.245 96.475 172.290 ;
        RECT 82.365 172.090 82.655 172.135 ;
        RECT 69.010 171.950 82.655 172.090 ;
        RECT 69.010 171.890 69.330 171.950 ;
        RECT 82.365 171.905 82.655 171.950 ;
        RECT 89.725 171.905 90.015 172.135 ;
        RECT 92.885 171.930 93.175 172.245 ;
        RECT 98.450 172.230 98.770 172.490 ;
        RECT 108.570 172.430 108.890 172.490 ;
        RECT 114.550 172.430 114.870 172.490 ;
        RECT 108.570 172.290 114.870 172.430 ;
        RECT 108.570 172.230 108.890 172.290 ;
        RECT 93.965 172.090 94.255 172.135 ;
        RECT 97.545 172.090 97.835 172.135 ;
        RECT 99.380 172.090 99.670 172.135 ;
        RECT 93.965 171.950 99.670 172.090 ;
        RECT 93.965 171.905 94.255 171.950 ;
        RECT 97.545 171.905 97.835 171.950 ;
        RECT 99.380 171.905 99.670 171.950 ;
        RECT 107.205 171.905 107.495 172.135 ;
        RECT 40.120 171.750 40.260 171.890 ;
        RECT 35.060 171.610 40.260 171.750 ;
        RECT 62.585 171.750 62.875 171.795 ;
        RECT 63.950 171.750 64.270 171.810 ;
        RECT 62.585 171.610 64.270 171.750 ;
        RECT 62.585 171.565 62.875 171.610 ;
        RECT 63.950 171.550 64.270 171.610 ;
        RECT 85.585 171.565 85.875 171.795 ;
        RECT 87.410 171.750 87.730 171.810 ;
        RECT 90.170 171.750 90.490 171.810 ;
        RECT 99.845 171.750 100.135 171.795 ;
        RECT 87.410 171.610 100.135 171.750 ;
        RECT 35.430 171.410 35.750 171.470 ;
        RECT 38.205 171.410 38.495 171.455 ;
        RECT 35.430 171.270 38.495 171.410 ;
        RECT 35.430 171.210 35.750 171.270 ;
        RECT 38.205 171.225 38.495 171.270 ;
        RECT 56.705 171.410 56.995 171.455 ;
        RECT 59.825 171.410 60.115 171.455 ;
        RECT 61.715 171.410 62.005 171.455 ;
        RECT 56.705 171.270 62.005 171.410 ;
        RECT 85.660 171.410 85.800 171.565 ;
        RECT 87.410 171.550 87.730 171.610 ;
        RECT 90.170 171.550 90.490 171.610 ;
        RECT 99.845 171.565 100.135 171.610 ;
        RECT 106.270 171.750 106.590 171.810 ;
        RECT 107.280 171.750 107.420 171.905 ;
        RECT 109.490 171.890 109.810 172.150 ;
        RECT 109.950 171.890 110.270 172.150 ;
        RECT 110.410 171.890 110.730 172.150 ;
        RECT 111.420 172.135 111.560 172.290 ;
        RECT 114.550 172.230 114.870 172.290 ;
        RECT 117.425 172.430 117.715 172.475 ;
        RECT 120.665 172.430 121.315 172.475 ;
        RECT 117.425 172.290 121.315 172.430 ;
        RECT 117.425 172.245 118.015 172.290 ;
        RECT 120.665 172.245 121.315 172.290 ;
        RECT 117.725 172.150 118.015 172.245 ;
        RECT 111.345 171.905 111.635 172.135 ;
        RECT 112.250 172.090 112.570 172.150 ;
        RECT 113.185 172.090 113.475 172.135 ;
        RECT 112.250 171.950 113.475 172.090 ;
        RECT 112.250 171.890 112.570 171.950 ;
        RECT 113.185 171.905 113.475 171.950 ;
        RECT 117.725 171.930 118.090 172.150 ;
        RECT 110.870 171.750 111.190 171.810 ;
        RECT 106.270 171.610 111.190 171.750 ;
        RECT 113.260 171.750 113.400 171.905 ;
        RECT 117.770 171.890 118.090 171.930 ;
        RECT 118.805 172.090 119.095 172.135 ;
        RECT 122.385 172.090 122.675 172.135 ;
        RECT 124.220 172.090 124.510 172.135 ;
        RECT 118.805 171.950 124.510 172.090 ;
        RECT 118.805 171.905 119.095 171.950 ;
        RECT 122.385 171.905 122.675 171.950 ;
        RECT 124.220 171.905 124.510 171.950 ;
        RECT 124.670 171.890 124.990 172.150 ;
        RECT 117.310 171.750 117.630 171.810 ;
        RECT 120.530 171.750 120.850 171.810 ;
        RECT 113.260 171.610 120.850 171.750 ;
        RECT 106.270 171.550 106.590 171.610 ;
        RECT 110.870 171.550 111.190 171.610 ;
        RECT 117.310 171.550 117.630 171.610 ;
        RECT 120.530 171.550 120.850 171.610 ;
        RECT 123.305 171.750 123.595 171.795 ;
        RECT 123.305 171.610 124.440 171.750 ;
        RECT 123.305 171.565 123.595 171.610 ;
        RECT 91.105 171.410 91.395 171.455 ;
        RECT 85.660 171.270 91.395 171.410 ;
        RECT 56.705 171.225 56.995 171.270 ;
        RECT 59.825 171.225 60.115 171.270 ;
        RECT 61.715 171.225 62.005 171.270 ;
        RECT 91.105 171.225 91.395 171.270 ;
        RECT 93.965 171.410 94.255 171.455 ;
        RECT 97.085 171.410 97.375 171.455 ;
        RECT 98.975 171.410 99.265 171.455 ;
        RECT 112.250 171.410 112.570 171.470 ;
        RECT 93.965 171.270 99.265 171.410 ;
        RECT 93.965 171.225 94.255 171.270 ;
        RECT 97.085 171.225 97.375 171.270 ;
        RECT 98.975 171.225 99.265 171.270 ;
        RECT 107.740 171.270 112.570 171.410 ;
        RECT 35.890 171.070 36.210 171.130 ;
        RECT 36.825 171.070 37.115 171.115 ;
        RECT 35.890 170.930 37.115 171.070 ;
        RECT 35.890 170.870 36.210 170.930 ;
        RECT 36.825 170.885 37.115 170.930 ;
        RECT 46.945 171.070 47.235 171.115 ;
        RECT 57.510 171.070 57.830 171.130 ;
        RECT 46.945 170.930 57.830 171.070 ;
        RECT 46.945 170.885 47.235 170.930 ;
        RECT 57.510 170.870 57.830 170.930 ;
        RECT 88.345 171.070 88.635 171.115 ;
        RECT 90.630 171.070 90.950 171.130 ;
        RECT 88.345 170.930 90.950 171.070 ;
        RECT 91.180 171.070 91.320 171.225 ;
        RECT 107.740 171.130 107.880 171.270 ;
        RECT 112.250 171.210 112.570 171.270 ;
        RECT 118.805 171.410 119.095 171.455 ;
        RECT 121.925 171.410 122.215 171.455 ;
        RECT 123.815 171.410 124.105 171.455 ;
        RECT 118.805 171.270 124.105 171.410 ;
        RECT 118.805 171.225 119.095 171.270 ;
        RECT 121.925 171.225 122.215 171.270 ;
        RECT 123.815 171.225 124.105 171.270 ;
        RECT 124.300 171.130 124.440 171.610 ;
        RECT 107.650 171.070 107.970 171.130 ;
        RECT 91.180 170.930 107.970 171.070 ;
        RECT 88.345 170.885 88.635 170.930 ;
        RECT 90.630 170.870 90.950 170.930 ;
        RECT 107.650 170.870 107.970 170.930 ;
        RECT 108.125 171.070 108.415 171.115 ;
        RECT 109.030 171.070 109.350 171.130 ;
        RECT 108.125 170.930 109.350 171.070 ;
        RECT 108.125 170.885 108.415 170.930 ;
        RECT 109.030 170.870 109.350 170.930 ;
        RECT 113.630 170.870 113.950 171.130 ;
        RECT 115.470 171.070 115.790 171.130 ;
        RECT 115.945 171.070 116.235 171.115 ;
        RECT 115.470 170.930 116.235 171.070 ;
        RECT 115.470 170.870 115.790 170.930 ;
        RECT 115.945 170.885 116.235 170.930 ;
        RECT 124.210 170.870 124.530 171.130 ;
        RECT 56.590 170.050 56.910 170.110 ;
        RECT 64.410 170.050 64.730 170.110 ;
        RECT 56.590 169.910 64.730 170.050 ;
        RECT 56.590 169.850 56.910 169.910 ;
        RECT 64.410 169.850 64.730 169.910 ;
        RECT 70.865 170.050 71.155 170.095 ;
        RECT 78.210 170.050 78.530 170.110 ;
        RECT 92.010 170.050 92.330 170.110 ;
        RECT 93.850 170.050 94.170 170.110 ;
        RECT 70.865 169.910 78.530 170.050 ;
        RECT 70.865 169.865 71.155 169.910 ;
        RECT 41.410 169.710 41.730 169.770 ;
        RECT 43.250 169.710 43.570 169.770 ;
        RECT 70.940 169.710 71.080 169.865 ;
        RECT 78.210 169.850 78.530 169.910 ;
        RECT 78.760 169.910 94.170 170.050 ;
        RECT 41.410 169.570 71.080 169.710 ;
        RECT 41.410 169.510 41.730 169.570 ;
        RECT 43.250 169.510 43.570 169.570 ;
        RECT 78.760 169.430 78.900 169.910 ;
        RECT 92.010 169.850 92.330 169.910 ;
        RECT 93.850 169.850 94.170 169.910 ;
        RECT 97.085 170.050 97.375 170.095 ;
        RECT 98.450 170.050 98.770 170.110 ;
        RECT 97.085 169.910 98.770 170.050 ;
        RECT 97.085 169.865 97.375 169.910 ;
        RECT 98.450 169.850 98.770 169.910 ;
        RECT 123.765 170.050 124.055 170.095 ;
        RECT 124.210 170.050 124.530 170.110 ;
        RECT 123.765 169.910 124.530 170.050 ;
        RECT 123.765 169.865 124.055 169.910 ;
        RECT 124.210 169.850 124.530 169.910 ;
        RECT 84.620 169.710 84.910 169.755 ;
        RECT 87.400 169.710 87.690 169.755 ;
        RECT 89.260 169.710 89.550 169.755 ;
        RECT 84.620 169.570 89.550 169.710 ;
        RECT 84.620 169.525 84.910 169.570 ;
        RECT 87.400 169.525 87.690 169.570 ;
        RECT 89.260 169.525 89.550 169.570 ;
        RECT 90.630 169.710 90.950 169.770 ;
        RECT 105.465 169.710 105.755 169.755 ;
        RECT 108.585 169.710 108.875 169.755 ;
        RECT 110.475 169.710 110.765 169.755 ;
        RECT 124.670 169.710 124.990 169.770 ;
        RECT 90.630 169.570 92.700 169.710 ;
        RECT 90.630 169.510 90.950 169.570 ;
        RECT 36.350 169.370 36.670 169.430 ;
        RECT 73.150 169.370 73.470 169.430 ;
        RECT 36.350 169.230 48.080 169.370 ;
        RECT 36.350 169.170 36.670 169.230 ;
        RECT 22.550 169.030 22.870 169.090 ;
        RECT 27.625 169.030 27.915 169.075 ;
        RECT 22.550 168.890 27.915 169.030 ;
        RECT 22.550 168.830 22.870 168.890 ;
        RECT 27.625 168.845 27.915 168.890 ;
        RECT 28.085 169.030 28.375 169.075 ;
        RECT 31.290 169.030 31.610 169.090 ;
        RECT 28.085 168.890 31.610 169.030 ;
        RECT 28.085 168.845 28.375 168.890 ;
        RECT 31.290 168.830 31.610 168.890 ;
        RECT 32.225 169.030 32.515 169.075 ;
        RECT 34.050 169.030 34.370 169.090 ;
        RECT 32.225 168.890 34.370 169.030 ;
        RECT 32.225 168.845 32.515 168.890 ;
        RECT 34.050 168.830 34.370 168.890 ;
        RECT 37.730 168.830 38.050 169.090 ;
        RECT 44.630 169.030 44.950 169.090 ;
        RECT 47.940 169.075 48.080 169.230 ;
        RECT 71.860 169.230 73.470 169.370 ;
        RECT 46.945 169.030 47.235 169.075 ;
        RECT 44.630 168.890 47.235 169.030 ;
        RECT 44.630 168.830 44.950 168.890 ;
        RECT 46.945 168.845 47.235 168.890 ;
        RECT 47.405 168.845 47.695 169.075 ;
        RECT 47.865 168.845 48.155 169.075 ;
        RECT 48.785 168.845 49.075 169.075 ;
        RECT 54.765 169.030 55.055 169.075 ;
        RECT 57.510 169.030 57.830 169.090 ;
        RECT 54.765 168.890 57.830 169.030 ;
        RECT 54.765 168.845 55.055 168.890 ;
        RECT 47.480 168.690 47.620 168.845 ;
        RECT 48.310 168.690 48.630 168.750 ;
        RECT 47.480 168.550 48.630 168.690 ;
        RECT 48.310 168.490 48.630 168.550 ;
        RECT 27.610 168.350 27.930 168.410 ;
        RECT 30.845 168.350 31.135 168.395 ;
        RECT 27.610 168.210 31.135 168.350 ;
        RECT 27.610 168.150 27.930 168.210 ;
        RECT 30.845 168.165 31.135 168.210 ;
        RECT 34.970 168.150 35.290 168.410 ;
        RECT 41.410 168.350 41.730 168.410 ;
        RECT 45.565 168.350 45.855 168.395 ;
        RECT 41.410 168.210 45.855 168.350 ;
        RECT 48.860 168.350 49.000 168.845 ;
        RECT 57.510 168.830 57.830 168.890 ;
        RECT 68.565 169.030 68.855 169.075 ;
        RECT 71.310 169.030 71.630 169.090 ;
        RECT 71.860 169.075 72.000 169.230 ;
        RECT 73.150 169.170 73.470 169.230 ;
        RECT 74.545 169.370 74.835 169.415 ;
        RECT 76.845 169.370 77.135 169.415 ;
        RECT 78.670 169.370 78.990 169.430 ;
        RECT 89.725 169.370 90.015 169.415 ;
        RECT 90.170 169.370 90.490 169.430 ;
        RECT 74.545 169.230 78.990 169.370 ;
        RECT 74.545 169.185 74.835 169.230 ;
        RECT 76.845 169.185 77.135 169.230 ;
        RECT 78.670 169.170 78.990 169.230 ;
        RECT 80.830 169.230 88.560 169.370 ;
        RECT 71.785 169.030 72.075 169.075 ;
        RECT 68.565 168.890 72.075 169.030 ;
        RECT 68.565 168.845 68.855 168.890 ;
        RECT 71.310 168.830 71.630 168.890 ;
        RECT 71.785 168.845 72.075 168.890 ;
        RECT 72.230 168.690 72.550 168.750 ;
        RECT 80.830 168.735 80.970 169.230 ;
        RECT 84.620 169.030 84.910 169.075 ;
        RECT 87.410 169.030 87.730 169.090 ;
        RECT 87.885 169.030 88.175 169.075 ;
        RECT 84.620 168.890 87.155 169.030 ;
        RECT 84.620 168.845 84.910 168.890 ;
        RECT 73.165 168.690 73.455 168.735 ;
        RECT 80.755 168.690 81.045 168.735 ;
        RECT 72.230 168.550 73.455 168.690 ;
        RECT 72.230 168.490 72.550 168.550 ;
        RECT 73.165 168.505 73.455 168.550 ;
        RECT 77.840 168.550 81.045 168.690 ;
        RECT 64.870 168.350 65.190 168.410 ;
        RECT 69.485 168.350 69.775 168.395 ;
        RECT 48.860 168.210 69.775 168.350 ;
        RECT 41.410 168.150 41.730 168.210 ;
        RECT 45.565 168.165 45.855 168.210 ;
        RECT 64.870 168.150 65.190 168.210 ;
        RECT 69.485 168.165 69.775 168.210 ;
        RECT 76.370 168.350 76.690 168.410 ;
        RECT 77.840 168.395 77.980 168.550 ;
        RECT 80.755 168.505 81.045 168.550 ;
        RECT 82.760 168.690 83.050 168.735 ;
        RECT 84.190 168.690 84.510 168.750 ;
        RECT 86.940 168.735 87.155 168.890 ;
        RECT 87.410 168.890 88.175 169.030 ;
        RECT 88.420 169.030 88.560 169.230 ;
        RECT 89.725 169.230 90.490 169.370 ;
        RECT 89.725 169.185 90.015 169.230 ;
        RECT 90.170 169.170 90.490 169.230 ;
        RECT 92.010 169.170 92.330 169.430 ;
        RECT 92.560 169.415 92.700 169.570 ;
        RECT 105.465 169.570 110.765 169.710 ;
        RECT 105.465 169.525 105.755 169.570 ;
        RECT 108.585 169.525 108.875 169.570 ;
        RECT 110.475 169.525 110.765 169.570 ;
        RECT 111.880 169.570 124.990 169.710 ;
        RECT 92.485 169.185 92.775 169.415 ;
        RECT 111.330 169.370 111.650 169.430 ;
        RECT 111.880 169.370 112.020 169.570 ;
        RECT 124.670 169.510 124.990 169.570 ;
        RECT 111.330 169.230 112.020 169.370 ;
        RECT 112.710 169.370 113.030 169.430 ;
        RECT 115.485 169.370 115.775 169.415 ;
        RECT 112.710 169.230 115.775 169.370 ;
        RECT 111.330 169.170 111.650 169.230 ;
        RECT 112.710 169.170 113.030 169.230 ;
        RECT 115.485 169.185 115.775 169.230 ;
        RECT 116.390 169.370 116.710 169.430 ;
        RECT 119.625 169.370 119.915 169.415 ;
        RECT 116.390 169.230 119.915 169.370 ;
        RECT 116.390 169.170 116.710 169.230 ;
        RECT 119.625 169.185 119.915 169.230 ;
        RECT 92.945 169.030 93.235 169.075 ;
        RECT 96.165 169.030 96.455 169.075 ;
        RECT 104.430 169.050 104.750 169.090 ;
        RECT 88.420 168.890 93.235 169.030 ;
        RECT 87.410 168.830 87.730 168.890 ;
        RECT 87.885 168.845 88.175 168.890 ;
        RECT 92.945 168.845 93.235 168.890 ;
        RECT 94.860 168.890 96.455 169.030 ;
        RECT 86.020 168.690 86.310 168.735 ;
        RECT 82.760 168.550 86.310 168.690 ;
        RECT 82.760 168.505 83.050 168.550 ;
        RECT 84.190 168.490 84.510 168.550 ;
        RECT 86.020 168.505 86.310 168.550 ;
        RECT 86.940 168.690 87.230 168.735 ;
        RECT 88.800 168.690 89.090 168.735 ;
        RECT 86.940 168.550 89.090 168.690 ;
        RECT 86.940 168.505 87.230 168.550 ;
        RECT 88.800 168.505 89.090 168.550 ;
        RECT 77.765 168.350 78.055 168.395 ;
        RECT 76.370 168.210 78.055 168.350 ;
        RECT 76.370 168.150 76.690 168.210 ;
        RECT 77.765 168.165 78.055 168.210 ;
        RECT 78.210 168.150 78.530 168.410 ;
        RECT 80.065 168.350 80.355 168.395 ;
        RECT 83.270 168.350 83.590 168.410 ;
        RECT 94.860 168.395 95.000 168.890 ;
        RECT 96.165 168.845 96.455 168.890 ;
        RECT 104.385 168.830 104.750 169.050 ;
        RECT 105.465 169.030 105.755 169.075 ;
        RECT 109.045 169.030 109.335 169.075 ;
        RECT 110.880 169.030 111.170 169.075 ;
        RECT 105.465 168.890 111.170 169.030 ;
        RECT 105.465 168.845 105.755 168.890 ;
        RECT 109.045 168.845 109.335 168.890 ;
        RECT 110.880 168.845 111.170 168.890 ;
        RECT 112.250 169.030 112.570 169.090 ;
        RECT 114.565 169.030 114.855 169.075 ;
        RECT 112.250 168.890 114.855 169.030 ;
        RECT 112.250 168.830 112.570 168.890 ;
        RECT 114.565 168.845 114.855 168.890 ;
        RECT 115.025 169.030 115.315 169.075 ;
        RECT 116.865 169.030 117.155 169.075 ;
        RECT 115.025 168.890 117.155 169.030 ;
        RECT 115.025 168.845 115.315 168.890 ;
        RECT 116.865 168.845 117.155 168.890 ;
        RECT 120.530 168.830 120.850 169.090 ;
        RECT 124.685 169.030 124.975 169.075 ;
        RECT 121.080 168.890 124.975 169.030 ;
        RECT 104.385 168.735 104.675 168.830 ;
        RECT 104.085 168.690 104.675 168.735 ;
        RECT 107.325 168.690 107.975 168.735 ;
        RECT 104.085 168.550 107.975 168.690 ;
        RECT 104.085 168.505 104.375 168.550 ;
        RECT 107.325 168.505 107.975 168.550 ;
        RECT 109.950 168.490 110.270 168.750 ;
        RECT 110.410 168.690 110.730 168.750 ;
        RECT 121.080 168.690 121.220 168.890 ;
        RECT 124.685 168.845 124.975 168.890 ;
        RECT 110.410 168.550 121.220 168.690 ;
        RECT 121.450 168.690 121.770 168.750 ;
        RECT 121.925 168.690 122.215 168.735 ;
        RECT 121.450 168.550 122.215 168.690 ;
        RECT 110.410 168.490 110.730 168.550 ;
        RECT 121.450 168.490 121.770 168.550 ;
        RECT 121.925 168.505 122.215 168.550 ;
        RECT 80.065 168.210 83.590 168.350 ;
        RECT 80.065 168.165 80.355 168.210 ;
        RECT 83.270 168.150 83.590 168.210 ;
        RECT 94.785 168.165 95.075 168.395 ;
        RECT 102.590 168.150 102.910 168.410 ;
        RECT 112.250 168.350 112.570 168.410 ;
        RECT 112.725 168.350 113.015 168.395 ;
        RECT 112.250 168.210 113.015 168.350 ;
        RECT 112.250 168.150 112.570 168.210 ;
        RECT 112.725 168.165 113.015 168.210 ;
        RECT 120.990 168.150 121.310 168.410 ;
        RECT 31.290 167.330 31.610 167.390 ;
        RECT 31.290 167.190 37.040 167.330 ;
        RECT 31.290 167.130 31.610 167.190 ;
        RECT 19.905 166.990 20.195 167.035 ;
        RECT 22.550 166.990 22.870 167.050 ;
        RECT 23.145 166.990 23.795 167.035 ;
        RECT 19.905 166.850 23.795 166.990 ;
        RECT 19.905 166.805 20.495 166.850 ;
        RECT 20.205 166.490 20.495 166.805 ;
        RECT 22.550 166.790 22.870 166.850 ;
        RECT 23.145 166.805 23.795 166.850 ;
        RECT 21.285 166.650 21.575 166.695 ;
        RECT 24.865 166.650 25.155 166.695 ;
        RECT 26.700 166.650 26.990 166.695 ;
        RECT 21.285 166.510 26.990 166.650 ;
        RECT 21.285 166.465 21.575 166.510 ;
        RECT 24.865 166.465 25.155 166.510 ;
        RECT 26.700 166.465 26.990 166.510 ;
        RECT 36.350 166.450 36.670 166.710 ;
        RECT 36.900 166.650 37.040 167.190 ;
        RECT 37.745 167.145 38.035 167.375 ;
        RECT 64.410 167.330 64.730 167.390 ;
        RECT 64.410 167.190 71.310 167.330 ;
        RECT 37.270 166.990 37.590 167.050 ;
        RECT 37.820 166.990 37.960 167.145 ;
        RECT 64.410 167.130 64.730 167.190 ;
        RECT 42.805 166.990 43.095 167.035 ;
        RECT 48.885 166.990 49.175 167.035 ;
        RECT 52.125 166.990 52.775 167.035 ;
        RECT 37.270 166.850 37.960 166.990 ;
        RECT 38.280 166.850 40.260 166.990 ;
        RECT 37.270 166.790 37.590 166.850 ;
        RECT 38.280 166.650 38.420 166.850 ;
        RECT 36.900 166.510 38.420 166.650 ;
        RECT 38.650 166.450 38.970 166.710 ;
        RECT 40.120 166.695 40.260 166.850 ;
        RECT 42.805 166.850 52.775 166.990 ;
        RECT 42.805 166.805 43.095 166.850 ;
        RECT 48.885 166.805 49.475 166.850 ;
        RECT 52.125 166.805 52.775 166.850 ;
        RECT 54.290 166.990 54.610 167.050 ;
        RECT 65.420 167.035 65.560 167.190 ;
        RECT 54.290 166.850 58.660 166.990 ;
        RECT 40.045 166.465 40.335 166.695 ;
        RECT 25.770 166.110 26.090 166.370 ;
        RECT 27.150 166.310 27.470 166.370 ;
        RECT 34.970 166.310 35.290 166.370 ;
        RECT 40.120 166.310 40.260 166.465 ;
        RECT 40.950 166.450 41.270 166.710 ;
        RECT 42.345 166.650 42.635 166.695 ;
        RECT 42.345 166.510 48.080 166.650 ;
        RECT 42.345 166.465 42.635 166.510 ;
        RECT 42.420 166.310 42.560 166.465 ;
        RECT 27.150 166.170 30.140 166.310 ;
        RECT 27.150 166.110 27.470 166.170 ;
        RECT 30.000 166.015 30.140 166.170 ;
        RECT 34.970 166.170 38.420 166.310 ;
        RECT 40.120 166.170 42.560 166.310 ;
        RECT 44.185 166.310 44.475 166.355 ;
        RECT 47.940 166.310 48.080 166.510 ;
        RECT 49.185 166.490 49.475 166.805 ;
        RECT 54.290 166.790 54.610 166.850 ;
        RECT 58.520 166.695 58.660 166.850 ;
        RECT 65.345 166.805 65.635 167.035 ;
        RECT 68.550 166.990 68.870 167.050 ;
        RECT 71.170 166.990 71.310 167.190 ;
        RECT 110.410 167.130 110.730 167.390 ;
        RECT 73.610 166.990 73.930 167.050 ;
        RECT 68.550 166.850 69.700 166.990 ;
        RECT 71.170 166.850 73.930 166.990 ;
        RECT 68.550 166.790 68.870 166.850 ;
        RECT 50.265 166.650 50.555 166.695 ;
        RECT 53.845 166.650 54.135 166.695 ;
        RECT 55.680 166.650 55.970 166.695 ;
        RECT 50.265 166.510 55.970 166.650 ;
        RECT 50.265 166.465 50.555 166.510 ;
        RECT 53.845 166.465 54.135 166.510 ;
        RECT 55.680 166.465 55.970 166.510 ;
        RECT 58.445 166.650 58.735 166.695 ;
        RECT 60.745 166.650 61.035 166.695 ;
        RECT 58.445 166.510 61.035 166.650 ;
        RECT 58.445 166.465 58.735 166.510 ;
        RECT 60.745 166.465 61.035 166.510 ;
        RECT 62.125 166.650 62.415 166.695 ;
        RECT 64.410 166.650 64.730 166.710 ;
        RECT 66.725 166.650 67.015 166.695 ;
        RECT 69.025 166.650 69.315 166.695 ;
        RECT 62.125 166.510 69.315 166.650 ;
        RECT 69.560 166.650 69.700 166.850 ;
        RECT 73.610 166.790 73.930 166.850 ;
        RECT 77.700 166.990 77.990 167.035 ;
        RECT 80.960 166.990 81.250 167.035 ;
        RECT 77.700 166.850 81.250 166.990 ;
        RECT 77.700 166.805 77.990 166.850 ;
        RECT 69.930 166.650 70.250 166.710 ;
        RECT 71.325 166.650 71.615 166.695 ;
        RECT 69.560 166.510 71.615 166.650 ;
        RECT 62.125 166.465 62.415 166.510 ;
        RECT 64.410 166.450 64.730 166.510 ;
        RECT 66.725 166.465 67.015 166.510 ;
        RECT 69.025 166.465 69.315 166.510 ;
        RECT 69.930 166.450 70.250 166.510 ;
        RECT 71.325 166.465 71.615 166.510 ;
        RECT 73.150 166.450 73.470 166.710 ;
        RECT 54.290 166.310 54.610 166.370 ;
        RECT 44.185 166.170 47.620 166.310 ;
        RECT 47.940 166.170 54.610 166.310 ;
        RECT 34.970 166.110 35.290 166.170 ;
        RECT 21.285 165.970 21.575 166.015 ;
        RECT 24.405 165.970 24.695 166.015 ;
        RECT 26.295 165.970 26.585 166.015 ;
        RECT 21.285 165.830 26.585 165.970 ;
        RECT 21.285 165.785 21.575 165.830 ;
        RECT 24.405 165.785 24.695 165.830 ;
        RECT 26.295 165.785 26.585 165.830 ;
        RECT 29.925 165.970 30.215 166.015 ;
        RECT 37.730 165.970 38.050 166.030 ;
        RECT 29.925 165.830 38.050 165.970 ;
        RECT 38.280 165.970 38.420 166.170 ;
        RECT 44.185 166.125 44.475 166.170 ;
        RECT 45.550 165.970 45.870 166.030 ;
        RECT 38.280 165.830 45.870 165.970 ;
        RECT 29.925 165.785 30.215 165.830 ;
        RECT 37.730 165.770 38.050 165.830 ;
        RECT 45.550 165.770 45.870 165.830 ;
        RECT 18.425 165.630 18.715 165.675 ;
        RECT 34.050 165.630 34.370 165.690 ;
        RECT 18.425 165.490 34.370 165.630 ;
        RECT 18.425 165.445 18.715 165.490 ;
        RECT 34.050 165.430 34.370 165.490 ;
        RECT 39.585 165.630 39.875 165.675 ;
        RECT 40.030 165.630 40.350 165.690 ;
        RECT 39.585 165.490 40.350 165.630 ;
        RECT 39.585 165.445 39.875 165.490 ;
        RECT 40.030 165.430 40.350 165.490 ;
        RECT 41.870 165.430 42.190 165.690 ;
        RECT 46.930 165.430 47.250 165.690 ;
        RECT 47.480 165.675 47.620 166.170 ;
        RECT 54.290 166.110 54.610 166.170 ;
        RECT 54.750 166.110 55.070 166.370 ;
        RECT 56.145 166.310 56.435 166.355 ;
        RECT 57.510 166.310 57.830 166.370 ;
        RECT 63.950 166.310 64.270 166.370 ;
        RECT 56.145 166.170 64.270 166.310 ;
        RECT 56.145 166.125 56.435 166.170 ;
        RECT 57.510 166.110 57.830 166.170 ;
        RECT 63.950 166.110 64.270 166.170 ;
        RECT 67.630 166.310 67.950 166.370 ;
        RECT 71.785 166.310 72.075 166.355 ;
        RECT 72.705 166.310 72.995 166.355 ;
        RECT 67.630 166.170 72.075 166.310 ;
        RECT 72.595 166.170 72.995 166.310 ;
        RECT 79.220 166.310 79.360 166.850 ;
        RECT 80.960 166.805 81.250 166.850 ;
        RECT 81.880 166.990 82.170 167.035 ;
        RECT 83.740 166.990 84.030 167.035 ;
        RECT 81.880 166.850 84.030 166.990 ;
        RECT 81.880 166.805 82.170 166.850 ;
        RECT 83.740 166.805 84.030 166.850 ;
        RECT 84.190 166.990 84.510 167.050 ;
        RECT 86.965 166.990 87.255 167.035 ;
        RECT 84.190 166.850 87.255 166.990 ;
        RECT 79.560 166.650 79.850 166.695 ;
        RECT 81.880 166.650 82.095 166.805 ;
        RECT 84.190 166.790 84.510 166.850 ;
        RECT 86.965 166.805 87.255 166.850 ;
        RECT 99.320 166.990 99.610 167.035 ;
        RECT 101.670 166.990 101.990 167.050 ;
        RECT 120.990 167.035 121.310 167.050 ;
        RECT 102.580 166.990 102.870 167.035 ;
        RECT 99.320 166.850 102.870 166.990 ;
        RECT 99.320 166.805 99.610 166.850 ;
        RECT 101.670 166.790 101.990 166.850 ;
        RECT 102.580 166.805 102.870 166.850 ;
        RECT 103.500 166.990 103.790 167.035 ;
        RECT 105.360 166.990 105.650 167.035 ;
        RECT 103.500 166.850 105.650 166.990 ;
        RECT 103.500 166.805 103.790 166.850 ;
        RECT 105.360 166.805 105.650 166.850 ;
        RECT 117.425 166.990 117.715 167.035 ;
        RECT 120.665 166.990 121.315 167.035 ;
        RECT 117.425 166.850 121.315 166.990 ;
        RECT 117.425 166.805 118.015 166.850 ;
        RECT 120.665 166.805 121.315 166.850 ;
        RECT 85.585 166.650 85.875 166.695 ;
        RECT 79.560 166.510 82.095 166.650 ;
        RECT 82.440 166.510 85.875 166.650 ;
        RECT 79.560 166.465 79.850 166.510 ;
        RECT 82.440 166.310 82.580 166.510 ;
        RECT 85.585 166.465 85.875 166.510 ;
        RECT 86.045 166.650 86.335 166.695 ;
        RECT 87.425 166.650 87.715 166.695 ;
        RECT 95.690 166.650 96.010 166.710 ;
        RECT 86.045 166.510 96.010 166.650 ;
        RECT 86.045 166.465 86.335 166.510 ;
        RECT 87.425 166.465 87.715 166.510 ;
        RECT 95.690 166.450 96.010 166.510 ;
        RECT 101.180 166.650 101.470 166.695 ;
        RECT 103.500 166.650 103.715 166.805 ;
        RECT 101.180 166.510 103.715 166.650 ;
        RECT 101.180 166.465 101.470 166.510 ;
        RECT 106.270 166.450 106.590 166.710 ;
        RECT 107.665 166.650 107.955 166.695 ;
        RECT 112.250 166.650 112.570 166.710 ;
        RECT 107.665 166.510 112.570 166.650 ;
        RECT 107.665 166.465 107.955 166.510 ;
        RECT 112.250 166.450 112.570 166.510 ;
        RECT 117.725 166.490 118.015 166.805 ;
        RECT 120.990 166.790 121.310 166.805 ;
        RECT 118.805 166.650 119.095 166.695 ;
        RECT 122.385 166.650 122.675 166.695 ;
        RECT 124.220 166.650 124.510 166.695 ;
        RECT 118.805 166.510 124.510 166.650 ;
        RECT 118.805 166.465 119.095 166.510 ;
        RECT 122.385 166.465 122.675 166.510 ;
        RECT 124.220 166.465 124.510 166.510 ;
        RECT 124.670 166.450 124.990 166.710 ;
        RECT 79.220 166.170 82.580 166.310 ;
        RECT 67.630 166.110 67.950 166.170 ;
        RECT 71.785 166.125 72.075 166.170 ;
        RECT 72.705 166.125 72.995 166.170 ;
        RECT 50.265 165.970 50.555 166.015 ;
        RECT 53.385 165.970 53.675 166.015 ;
        RECT 55.275 165.970 55.565 166.015 ;
        RECT 50.265 165.830 55.565 165.970 ;
        RECT 50.265 165.785 50.555 165.830 ;
        RECT 53.385 165.785 53.675 165.830 ;
        RECT 55.275 165.785 55.565 165.830 ;
        RECT 69.470 165.970 69.790 166.030 ;
        RECT 72.780 165.970 72.920 166.125 ;
        RECT 82.810 166.110 83.130 166.370 ;
        RECT 84.665 166.310 84.955 166.355 ;
        RECT 90.170 166.310 90.490 166.370 ;
        RECT 84.665 166.170 90.490 166.310 ;
        RECT 84.665 166.125 84.955 166.170 ;
        RECT 90.170 166.110 90.490 166.170 ;
        RECT 100.750 166.310 101.070 166.370 ;
        RECT 104.445 166.310 104.735 166.355 ;
        RECT 100.750 166.170 104.735 166.310 ;
        RECT 100.750 166.110 101.070 166.170 ;
        RECT 104.445 166.125 104.735 166.170 ;
        RECT 113.170 166.310 113.490 166.370 ;
        RECT 113.645 166.310 113.935 166.355 ;
        RECT 115.945 166.310 116.235 166.355 ;
        RECT 113.170 166.170 116.235 166.310 ;
        RECT 113.170 166.110 113.490 166.170 ;
        RECT 113.645 166.125 113.935 166.170 ;
        RECT 115.945 166.125 116.235 166.170 ;
        RECT 123.305 166.310 123.595 166.355 ;
        RECT 123.305 166.170 124.440 166.310 ;
        RECT 123.305 166.125 123.595 166.170 ;
        RECT 74.530 165.970 74.850 166.030 ;
        RECT 69.470 165.830 74.850 165.970 ;
        RECT 69.470 165.770 69.790 165.830 ;
        RECT 74.530 165.770 74.850 165.830 ;
        RECT 79.560 165.970 79.850 166.015 ;
        RECT 82.340 165.970 82.630 166.015 ;
        RECT 84.200 165.970 84.490 166.015 ;
        RECT 79.560 165.830 84.490 165.970 ;
        RECT 79.560 165.785 79.850 165.830 ;
        RECT 82.340 165.785 82.630 165.830 ;
        RECT 84.200 165.785 84.490 165.830 ;
        RECT 101.180 165.970 101.470 166.015 ;
        RECT 103.960 165.970 104.250 166.015 ;
        RECT 105.820 165.970 106.110 166.015 ;
        RECT 101.180 165.830 106.110 165.970 ;
        RECT 101.180 165.785 101.470 165.830 ;
        RECT 103.960 165.785 104.250 165.830 ;
        RECT 105.820 165.785 106.110 165.830 ;
        RECT 118.805 165.970 119.095 166.015 ;
        RECT 121.925 165.970 122.215 166.015 ;
        RECT 123.815 165.970 124.105 166.015 ;
        RECT 118.805 165.830 124.105 165.970 ;
        RECT 118.805 165.785 119.095 165.830 ;
        RECT 121.925 165.785 122.215 165.830 ;
        RECT 123.815 165.785 124.105 165.830 ;
        RECT 124.300 165.690 124.440 166.170 ;
        RECT 47.405 165.630 47.695 165.675 ;
        RECT 48.770 165.630 49.090 165.690 ;
        RECT 47.405 165.490 49.090 165.630 ;
        RECT 47.405 165.445 47.695 165.490 ;
        RECT 48.770 165.430 49.090 165.490 ;
        RECT 57.985 165.630 58.275 165.675 ;
        RECT 58.430 165.630 58.750 165.690 ;
        RECT 57.985 165.490 58.750 165.630 ;
        RECT 57.985 165.445 58.275 165.490 ;
        RECT 58.430 165.430 58.750 165.490 ;
        RECT 68.565 165.630 68.855 165.675 ;
        RECT 69.010 165.630 69.330 165.690 ;
        RECT 68.565 165.490 69.330 165.630 ;
        RECT 68.565 165.445 68.855 165.490 ;
        RECT 69.010 165.430 69.330 165.490 ;
        RECT 72.230 165.430 72.550 165.690 ;
        RECT 73.150 165.630 73.470 165.690 ;
        RECT 75.695 165.630 75.985 165.675 ;
        RECT 73.150 165.490 75.985 165.630 ;
        RECT 73.150 165.430 73.470 165.490 ;
        RECT 75.695 165.445 75.985 165.490 ;
        RECT 97.315 165.630 97.605 165.675 ;
        RECT 100.290 165.630 100.610 165.690 ;
        RECT 97.315 165.490 100.610 165.630 ;
        RECT 97.315 165.445 97.605 165.490 ;
        RECT 100.290 165.430 100.610 165.490 ;
        RECT 110.870 165.430 111.190 165.690 ;
        RECT 124.210 165.430 124.530 165.690 ;
        RECT 25.770 164.410 26.090 164.670 ;
        RECT 37.730 164.610 38.050 164.670 ;
        RECT 67.645 164.610 67.935 164.655 ;
        RECT 37.730 164.470 45.320 164.610 ;
        RECT 37.730 164.410 38.050 164.470 ;
        RECT 30.025 164.270 30.315 164.315 ;
        RECT 33.145 164.270 33.435 164.315 ;
        RECT 35.035 164.270 35.325 164.315 ;
        RECT 37.270 164.270 37.590 164.330 ;
        RECT 30.025 164.130 35.325 164.270 ;
        RECT 30.025 164.085 30.315 164.130 ;
        RECT 33.145 164.085 33.435 164.130 ;
        RECT 35.035 164.085 35.325 164.130 ;
        RECT 35.520 164.130 37.590 164.270 ;
        RECT 34.525 163.930 34.815 163.975 ;
        RECT 35.520 163.930 35.660 164.130 ;
        RECT 37.270 164.070 37.590 164.130 ;
        RECT 39.225 164.270 39.515 164.315 ;
        RECT 42.345 164.270 42.635 164.315 ;
        RECT 44.235 164.270 44.525 164.315 ;
        RECT 39.225 164.130 44.525 164.270 ;
        RECT 39.225 164.085 39.515 164.130 ;
        RECT 42.345 164.085 42.635 164.130 ;
        RECT 44.235 164.085 44.525 164.130 ;
        RECT 34.525 163.790 35.660 163.930 ;
        RECT 35.905 163.930 36.195 163.975 ;
        RECT 37.730 163.930 38.050 163.990 ;
        RECT 35.905 163.790 38.050 163.930 ;
        RECT 34.525 163.745 34.815 163.790 ;
        RECT 35.905 163.745 36.195 163.790 ;
        RECT 37.730 163.730 38.050 163.790 ;
        RECT 41.870 163.930 42.190 163.990 ;
        RECT 45.180 163.975 45.320 164.470 ;
        RECT 52.080 164.470 67.935 164.610 ;
        RECT 43.725 163.930 44.015 163.975 ;
        RECT 41.870 163.790 44.015 163.930 ;
        RECT 41.870 163.730 42.190 163.790 ;
        RECT 43.725 163.745 44.015 163.790 ;
        RECT 45.105 163.745 45.395 163.975 ;
        RECT 45.550 163.930 45.870 163.990 ;
        RECT 48.785 163.930 49.075 163.975 ;
        RECT 51.070 163.930 51.390 163.990 ;
        RECT 51.545 163.930 51.835 163.975 ;
        RECT 52.080 163.930 52.220 164.470 ;
        RECT 67.645 164.425 67.935 164.470 ;
        RECT 82.810 164.610 83.130 164.670 ;
        RECT 83.285 164.610 83.575 164.655 ;
        RECT 82.810 164.470 83.575 164.610 ;
        RECT 82.810 164.410 83.130 164.470 ;
        RECT 83.285 164.425 83.575 164.470 ;
        RECT 86.505 164.610 86.795 164.655 ;
        RECT 87.410 164.610 87.730 164.670 ;
        RECT 86.505 164.470 87.730 164.610 ;
        RECT 86.505 164.425 86.795 164.470 ;
        RECT 87.410 164.410 87.730 164.470 ;
        RECT 104.430 164.610 104.750 164.670 ;
        RECT 111.345 164.610 111.635 164.655 ;
        RECT 104.430 164.470 111.635 164.610 ;
        RECT 104.430 164.410 104.750 164.470 ;
        RECT 111.345 164.425 111.635 164.470 ;
        RECT 57.625 164.270 57.915 164.315 ;
        RECT 60.745 164.270 61.035 164.315 ;
        RECT 62.635 164.270 62.925 164.315 ;
        RECT 57.625 164.130 62.925 164.270 ;
        RECT 57.625 164.085 57.915 164.130 ;
        RECT 60.745 164.085 61.035 164.130 ;
        RECT 62.635 164.085 62.925 164.130 ;
        RECT 81.905 164.085 82.195 164.315 ;
        RECT 116.045 164.270 116.335 164.315 ;
        RECT 119.165 164.270 119.455 164.315 ;
        RECT 121.055 164.270 121.345 164.315 ;
        RECT 98.080 164.130 109.720 164.270 ;
        RECT 45.550 163.790 48.080 163.930 ;
        RECT 45.550 163.730 45.870 163.790 ;
        RECT 26.690 163.390 27.010 163.650 ;
        RECT 27.610 163.250 27.930 163.310 ;
        RECT 28.945 163.295 29.235 163.610 ;
        RECT 30.025 163.590 30.315 163.635 ;
        RECT 33.605 163.590 33.895 163.635 ;
        RECT 35.440 163.590 35.730 163.635 ;
        RECT 30.025 163.450 35.730 163.590 ;
        RECT 30.025 163.405 30.315 163.450 ;
        RECT 33.605 163.405 33.895 163.450 ;
        RECT 35.440 163.405 35.730 163.450 ;
        RECT 38.145 163.295 38.435 163.610 ;
        RECT 39.225 163.590 39.515 163.635 ;
        RECT 42.805 163.590 43.095 163.635 ;
        RECT 44.640 163.590 44.930 163.635 ;
        RECT 39.225 163.450 44.930 163.590 ;
        RECT 39.225 163.405 39.515 163.450 ;
        RECT 42.805 163.405 43.095 163.450 ;
        RECT 44.640 163.405 44.930 163.450 ;
        RECT 46.930 163.590 47.250 163.650 ;
        RECT 47.405 163.590 47.695 163.635 ;
        RECT 46.930 163.450 47.695 163.590 ;
        RECT 47.940 163.590 48.080 163.790 ;
        RECT 48.785 163.790 52.220 163.930 ;
        RECT 53.830 163.930 54.150 163.990 ;
        RECT 54.765 163.930 55.055 163.975 ;
        RECT 53.830 163.790 55.055 163.930 ;
        RECT 48.785 163.745 49.075 163.790 ;
        RECT 51.070 163.730 51.390 163.790 ;
        RECT 51.545 163.745 51.835 163.790 ;
        RECT 53.830 163.730 54.150 163.790 ;
        RECT 54.765 163.745 55.055 163.790 ;
        RECT 78.670 163.730 78.990 163.990 ;
        RECT 52.465 163.590 52.755 163.635 ;
        RECT 47.940 163.450 52.755 163.590 ;
        RECT 46.930 163.390 47.250 163.450 ;
        RECT 47.405 163.405 47.695 163.450 ;
        RECT 52.465 163.405 52.755 163.450 ;
        RECT 28.645 163.250 29.235 163.295 ;
        RECT 31.885 163.250 32.535 163.295 ;
        RECT 27.610 163.110 32.535 163.250 ;
        RECT 27.610 163.050 27.930 163.110 ;
        RECT 28.645 163.065 28.935 163.110 ;
        RECT 31.885 163.065 32.535 163.110 ;
        RECT 37.845 163.250 38.435 163.295 ;
        RECT 40.030 163.250 40.350 163.310 ;
        RECT 41.085 163.250 41.735 163.295 ;
        RECT 37.845 163.110 41.735 163.250 ;
        RECT 37.845 163.065 38.135 163.110 ;
        RECT 40.030 163.050 40.350 163.110 ;
        RECT 41.085 163.065 41.735 163.110 ;
        RECT 43.710 163.250 44.030 163.310 ;
        RECT 56.545 163.295 56.835 163.610 ;
        RECT 57.625 163.590 57.915 163.635 ;
        RECT 61.205 163.590 61.495 163.635 ;
        RECT 63.040 163.590 63.330 163.635 ;
        RECT 57.625 163.450 63.330 163.590 ;
        RECT 57.625 163.405 57.915 163.450 ;
        RECT 61.205 163.405 61.495 163.450 ;
        RECT 63.040 163.405 63.330 163.450 ;
        RECT 63.505 163.590 63.795 163.635 ;
        RECT 63.950 163.590 64.270 163.650 ;
        RECT 63.505 163.450 64.270 163.590 ;
        RECT 63.505 163.405 63.795 163.450 ;
        RECT 63.950 163.390 64.270 163.450 ;
        RECT 69.025 163.590 69.315 163.635 ;
        RECT 72.230 163.590 72.550 163.650 ;
        RECT 69.025 163.450 72.550 163.590 ;
        RECT 69.025 163.405 69.315 163.450 ;
        RECT 72.230 163.390 72.550 163.450 ;
        RECT 73.150 163.590 73.470 163.650 ;
        RECT 78.210 163.590 78.530 163.650 ;
        RECT 79.605 163.590 79.895 163.635 ;
        RECT 73.150 163.450 79.895 163.590 ;
        RECT 81.980 163.590 82.120 164.085 ;
        RECT 93.850 163.930 94.170 163.990 ;
        RECT 98.080 163.975 98.220 164.130 ;
        RECT 98.005 163.930 98.295 163.975 ;
        RECT 93.850 163.790 98.295 163.930 ;
        RECT 93.850 163.730 94.170 163.790 ;
        RECT 98.005 163.745 98.295 163.790 ;
        RECT 102.590 163.930 102.910 163.990 ;
        RECT 104.430 163.930 104.750 163.990 ;
        RECT 109.580 163.975 109.720 164.130 ;
        RECT 116.045 164.130 121.345 164.270 ;
        RECT 116.045 164.085 116.335 164.130 ;
        RECT 119.165 164.085 119.455 164.130 ;
        RECT 121.055 164.085 121.345 164.130 ;
        RECT 104.905 163.930 105.195 163.975 ;
        RECT 109.045 163.930 109.335 163.975 ;
        RECT 102.590 163.790 109.335 163.930 ;
        RECT 102.590 163.730 102.910 163.790 ;
        RECT 104.430 163.730 104.750 163.790 ;
        RECT 104.905 163.745 105.195 163.790 ;
        RECT 109.045 163.745 109.335 163.790 ;
        RECT 109.505 163.930 109.795 163.975 ;
        RECT 112.710 163.930 113.030 163.990 ;
        RECT 109.505 163.790 113.030 163.930 ;
        RECT 109.505 163.745 109.795 163.790 ;
        RECT 112.710 163.730 113.030 163.790 ;
        RECT 121.925 163.930 122.215 163.975 ;
        RECT 124.670 163.930 124.990 163.990 ;
        RECT 121.925 163.790 124.990 163.930 ;
        RECT 121.925 163.745 122.215 163.790 ;
        RECT 124.670 163.730 124.990 163.790 ;
        RECT 82.365 163.590 82.655 163.635 ;
        RECT 81.980 163.450 82.655 163.590 ;
        RECT 73.150 163.390 73.470 163.450 ;
        RECT 78.210 163.390 78.530 163.450 ;
        RECT 79.605 163.405 79.895 163.450 ;
        RECT 82.365 163.405 82.655 163.450 ;
        RECT 83.270 163.590 83.590 163.650 ;
        RECT 85.585 163.590 85.875 163.635 ;
        RECT 83.270 163.450 85.875 163.590 ;
        RECT 83.270 163.390 83.590 163.450 ;
        RECT 85.585 163.405 85.875 163.450 ;
        RECT 99.385 163.590 99.675 163.635 ;
        RECT 102.145 163.590 102.435 163.635 ;
        RECT 99.385 163.450 102.435 163.590 ;
        RECT 99.385 163.405 99.675 163.450 ;
        RECT 102.145 163.405 102.435 163.450 ;
        RECT 108.110 163.590 108.430 163.650 ;
        RECT 111.805 163.590 112.095 163.635 ;
        RECT 108.110 163.450 112.095 163.590 ;
        RECT 108.110 163.390 108.430 163.450 ;
        RECT 111.805 163.405 112.095 163.450 ;
        RECT 47.865 163.250 48.155 163.295 ;
        RECT 43.710 163.110 48.155 163.250 ;
        RECT 43.710 163.050 44.030 163.110 ;
        RECT 47.865 163.065 48.155 163.110 ;
        RECT 56.245 163.250 56.835 163.295 ;
        RECT 58.430 163.250 58.750 163.310 ;
        RECT 59.485 163.250 60.135 163.295 ;
        RECT 56.245 163.110 60.135 163.250 ;
        RECT 56.245 163.065 56.535 163.110 ;
        RECT 58.430 163.050 58.750 163.110 ;
        RECT 59.485 163.065 60.135 163.110 ;
        RECT 62.110 163.050 62.430 163.310 ;
        RECT 95.245 163.250 95.535 163.295 ;
        RECT 113.630 163.250 113.950 163.310 ;
        RECT 114.965 163.295 115.255 163.610 ;
        RECT 116.045 163.590 116.335 163.635 ;
        RECT 119.625 163.590 119.915 163.635 ;
        RECT 121.460 163.590 121.750 163.635 ;
        RECT 116.045 163.450 121.750 163.590 ;
        RECT 116.045 163.405 116.335 163.450 ;
        RECT 119.625 163.405 119.915 163.450 ;
        RECT 121.460 163.405 121.750 163.450 ;
        RECT 123.290 163.390 123.610 163.650 ;
        RECT 114.665 163.250 115.255 163.295 ;
        RECT 117.905 163.250 118.555 163.295 ;
        RECT 95.245 163.110 99.140 163.250 ;
        RECT 95.245 163.065 95.535 163.110 ;
        RECT 26.230 162.910 26.550 162.970 ;
        RECT 27.165 162.910 27.455 162.955 ;
        RECT 26.230 162.770 27.455 162.910 ;
        RECT 26.230 162.710 26.550 162.770 ;
        RECT 27.165 162.725 27.455 162.770 ;
        RECT 35.890 162.910 36.210 162.970 ;
        RECT 36.365 162.910 36.655 162.955 ;
        RECT 43.800 162.910 43.940 163.050 ;
        RECT 35.890 162.770 43.940 162.910 ;
        RECT 35.890 162.710 36.210 162.770 ;
        RECT 36.365 162.725 36.655 162.770 ;
        RECT 45.550 162.710 45.870 162.970 ;
        RECT 51.530 162.910 51.850 162.970 ;
        RECT 52.005 162.910 52.295 162.955 ;
        RECT 51.530 162.770 52.295 162.910 ;
        RECT 51.530 162.710 51.850 162.770 ;
        RECT 52.005 162.725 52.295 162.770 ;
        RECT 54.290 162.710 54.610 162.970 ;
        RECT 80.065 162.910 80.355 162.955 ;
        RECT 80.510 162.910 80.830 162.970 ;
        RECT 80.065 162.770 80.830 162.910 ;
        RECT 80.065 162.725 80.355 162.770 ;
        RECT 80.510 162.710 80.830 162.770 ;
        RECT 90.630 162.910 90.950 162.970 ;
        RECT 94.785 162.910 95.075 162.955 ;
        RECT 90.630 162.770 95.075 162.910 ;
        RECT 90.630 162.710 90.950 162.770 ;
        RECT 94.785 162.725 95.075 162.770 ;
        RECT 97.070 162.710 97.390 162.970 ;
        RECT 99.000 162.955 99.140 163.110 ;
        RECT 113.630 163.110 118.555 163.250 ;
        RECT 113.630 163.050 113.950 163.110 ;
        RECT 114.665 163.065 114.955 163.110 ;
        RECT 117.905 163.065 118.555 163.110 ;
        RECT 120.545 163.065 120.835 163.295 ;
        RECT 98.925 162.910 99.215 162.955 ;
        RECT 100.290 162.910 100.610 162.970 ;
        RECT 98.925 162.770 100.610 162.910 ;
        RECT 98.925 162.725 99.215 162.770 ;
        RECT 100.290 162.710 100.610 162.770 ;
        RECT 101.210 162.710 101.530 162.970 ;
        RECT 106.730 162.710 107.050 162.970 ;
        RECT 108.570 162.710 108.890 162.970 ;
        RECT 109.490 162.910 109.810 162.970 ;
        RECT 113.185 162.910 113.475 162.955 ;
        RECT 109.490 162.770 113.475 162.910 ;
        RECT 120.620 162.910 120.760 163.065 ;
        RECT 122.385 162.910 122.675 162.955 ;
        RECT 120.620 162.770 122.675 162.910 ;
        RECT 109.490 162.710 109.810 162.770 ;
        RECT 113.185 162.725 113.475 162.770 ;
        RECT 122.385 162.725 122.675 162.770 ;
        RECT 26.690 161.890 27.010 161.950 ;
        RECT 27.625 161.890 27.915 161.935 ;
        RECT 26.690 161.750 27.915 161.890 ;
        RECT 26.690 161.690 27.010 161.750 ;
        RECT 27.625 161.705 27.915 161.750 ;
        RECT 29.925 161.890 30.215 161.935 ;
        RECT 34.970 161.890 35.290 161.950 ;
        RECT 29.925 161.750 35.290 161.890 ;
        RECT 29.925 161.705 30.215 161.750 ;
        RECT 34.970 161.690 35.290 161.750 ;
        RECT 36.825 161.890 37.115 161.935 ;
        RECT 38.650 161.890 38.970 161.950 ;
        RECT 36.825 161.750 38.970 161.890 ;
        RECT 36.825 161.705 37.115 161.750 ;
        RECT 38.650 161.690 38.970 161.750 ;
        RECT 40.950 161.890 41.270 161.950 ;
        RECT 41.885 161.890 42.175 161.935 ;
        RECT 40.950 161.750 42.175 161.890 ;
        RECT 40.950 161.690 41.270 161.750 ;
        RECT 41.885 161.705 42.175 161.750 ;
        RECT 59.825 161.890 60.115 161.935 ;
        RECT 62.110 161.890 62.430 161.950 ;
        RECT 59.825 161.750 62.430 161.890 ;
        RECT 59.825 161.705 60.115 161.750 ;
        RECT 62.110 161.690 62.430 161.750 ;
        RECT 80.510 161.890 80.830 161.950 ;
        RECT 83.285 161.890 83.575 161.935 ;
        RECT 80.510 161.750 83.575 161.890 ;
        RECT 80.510 161.690 80.830 161.750 ;
        RECT 83.285 161.705 83.575 161.750 ;
        RECT 85.585 161.705 85.875 161.935 ;
        RECT 89.495 161.890 89.785 161.935 ;
        RECT 90.630 161.890 90.950 161.950 ;
        RECT 87.960 161.750 90.950 161.890 ;
        RECT 18.870 161.550 19.190 161.610 ;
        RECT 20.200 161.550 20.490 161.595 ;
        RECT 23.460 161.550 23.750 161.595 ;
        RECT 18.870 161.410 23.750 161.550 ;
        RECT 18.870 161.350 19.190 161.410 ;
        RECT 20.200 161.365 20.490 161.410 ;
        RECT 23.460 161.365 23.750 161.410 ;
        RECT 24.380 161.550 24.670 161.595 ;
        RECT 26.240 161.550 26.530 161.595 ;
        RECT 24.380 161.410 26.530 161.550 ;
        RECT 24.380 161.365 24.670 161.410 ;
        RECT 26.240 161.365 26.530 161.410 ;
        RECT 50.165 161.550 50.455 161.595 ;
        RECT 51.530 161.550 51.850 161.610 ;
        RECT 52.465 161.550 52.755 161.595 ;
        RECT 50.165 161.410 52.755 161.550 ;
        RECT 50.165 161.365 50.455 161.410 ;
        RECT 22.060 161.210 22.350 161.255 ;
        RECT 24.380 161.210 24.595 161.365 ;
        RECT 51.530 161.350 51.850 161.410 ;
        RECT 52.465 161.365 52.755 161.410 ;
        RECT 67.630 161.550 67.950 161.610 ;
        RECT 78.670 161.550 78.990 161.610 ;
        RECT 67.630 161.410 68.780 161.550 ;
        RECT 67.630 161.350 67.950 161.410 ;
        RECT 22.060 161.070 24.595 161.210 ;
        RECT 22.060 161.025 22.350 161.070 ;
        RECT 27.150 161.010 27.470 161.270 ;
        RECT 29.465 161.025 29.755 161.255 ;
        RECT 25.325 160.870 25.615 160.915 ;
        RECT 25.770 160.870 26.090 160.930 ;
        RECT 25.325 160.730 26.090 160.870 ;
        RECT 25.325 160.685 25.615 160.730 ;
        RECT 25.770 160.670 26.090 160.730 ;
        RECT 22.060 160.530 22.350 160.575 ;
        RECT 24.840 160.530 25.130 160.575 ;
        RECT 26.700 160.530 26.990 160.575 ;
        RECT 22.060 160.390 26.990 160.530 ;
        RECT 22.060 160.345 22.350 160.390 ;
        RECT 24.840 160.345 25.130 160.390 ;
        RECT 26.700 160.345 26.990 160.390 ;
        RECT 18.195 160.190 18.485 160.235 ;
        RECT 21.630 160.190 21.950 160.250 ;
        RECT 29.540 160.190 29.680 161.025 ;
        RECT 34.970 161.010 35.290 161.270 ;
        RECT 45.105 161.210 45.395 161.255 ;
        RECT 45.550 161.210 45.870 161.270 ;
        RECT 45.105 161.070 45.870 161.210 ;
        RECT 45.105 161.025 45.395 161.070 ;
        RECT 45.550 161.010 45.870 161.070 ;
        RECT 47.405 161.210 47.695 161.255 ;
        RECT 52.910 161.210 53.230 161.270 ;
        RECT 53.830 161.210 54.150 161.270 ;
        RECT 47.405 161.070 54.150 161.210 ;
        RECT 47.405 161.025 47.695 161.070 ;
        RECT 52.910 161.010 53.230 161.070 ;
        RECT 53.830 161.010 54.150 161.070 ;
        RECT 54.290 161.210 54.610 161.270 ;
        RECT 58.905 161.210 59.195 161.255 ;
        RECT 54.290 161.070 59.195 161.210 ;
        RECT 54.290 161.010 54.610 161.070 ;
        RECT 58.905 161.025 59.195 161.070 ;
        RECT 66.265 161.210 66.555 161.255 ;
        RECT 67.720 161.210 67.860 161.350 ;
        RECT 68.640 161.255 68.780 161.410 ;
        RECT 78.670 161.410 82.580 161.550 ;
        RECT 78.670 161.350 78.990 161.410 ;
        RECT 66.265 161.070 67.860 161.210 ;
        RECT 66.265 161.025 66.555 161.070 ;
        RECT 68.105 161.025 68.395 161.255 ;
        RECT 68.565 161.025 68.855 161.255 ;
        RECT 69.930 161.210 70.250 161.270 ;
        RECT 70.405 161.210 70.695 161.255 ;
        RECT 69.930 161.070 70.695 161.210 ;
        RECT 30.845 160.870 31.135 160.915 ;
        RECT 30.845 160.730 31.520 160.870 ;
        RECT 30.845 160.685 31.135 160.730 ;
        RECT 31.380 160.590 31.520 160.730 ;
        RECT 34.065 160.685 34.355 160.915 ;
        RECT 31.290 160.530 31.610 160.590 ;
        RECT 34.140 160.530 34.280 160.685 ;
        RECT 34.510 160.670 34.830 160.930 ;
        RECT 51.070 160.870 51.390 160.930 ;
        RECT 35.060 160.730 51.390 160.870 ;
        RECT 35.060 160.530 35.200 160.730 ;
        RECT 51.070 160.670 51.390 160.730 ;
        RECT 52.005 160.685 52.295 160.915 ;
        RECT 54.765 160.685 55.055 160.915 ;
        RECT 68.180 160.870 68.320 161.025 ;
        RECT 69.930 161.010 70.250 161.070 ;
        RECT 70.405 161.025 70.695 161.070 ;
        RECT 81.445 161.025 81.735 161.255 ;
        RECT 70.020 160.870 70.160 161.010 ;
        RECT 68.180 160.730 70.160 160.870 ;
        RECT 31.290 160.390 35.200 160.530 ;
        RECT 48.770 160.530 49.090 160.590 ;
        RECT 52.080 160.530 52.220 160.685 ;
        RECT 48.770 160.390 52.220 160.530 ;
        RECT 54.305 160.530 54.595 160.575 ;
        RECT 54.840 160.530 54.980 160.685 ;
        RECT 72.230 160.530 72.550 160.590 ;
        RECT 54.305 160.390 54.980 160.530 ;
        RECT 67.260 160.390 72.550 160.530 ;
        RECT 81.520 160.530 81.660 161.025 ;
        RECT 82.440 160.915 82.580 161.410 ;
        RECT 83.745 161.025 84.035 161.255 ;
        RECT 85.660 161.210 85.800 161.705 ;
        RECT 86.505 161.210 86.795 161.255 ;
        RECT 85.660 161.070 86.795 161.210 ;
        RECT 86.505 161.025 86.795 161.070 ;
        RECT 82.365 160.685 82.655 160.915 ;
        RECT 83.270 160.870 83.590 160.930 ;
        RECT 83.820 160.870 83.960 161.025 ;
        RECT 87.960 160.870 88.100 161.750 ;
        RECT 89.495 161.705 89.785 161.750 ;
        RECT 90.630 161.690 90.950 161.750 ;
        RECT 100.750 161.690 101.070 161.950 ;
        RECT 101.670 161.690 101.990 161.950 ;
        RECT 108.570 161.890 108.890 161.950 ;
        RECT 109.965 161.890 110.255 161.935 ;
        RECT 111.805 161.890 112.095 161.935 ;
        RECT 108.570 161.750 112.095 161.890 ;
        RECT 108.570 161.690 108.890 161.750 ;
        RECT 109.965 161.705 110.255 161.750 ;
        RECT 111.805 161.705 112.095 161.750 ;
        RECT 114.105 161.705 114.395 161.935 ;
        RECT 115.470 161.890 115.790 161.950 ;
        RECT 116.865 161.890 117.155 161.935 ;
        RECT 115.470 161.750 117.155 161.890 ;
        RECT 91.500 161.550 91.790 161.595 ;
        RECT 93.850 161.550 94.170 161.610 ;
        RECT 94.760 161.550 95.050 161.595 ;
        RECT 91.500 161.410 95.050 161.550 ;
        RECT 91.500 161.365 91.790 161.410 ;
        RECT 93.850 161.350 94.170 161.410 ;
        RECT 94.760 161.365 95.050 161.410 ;
        RECT 95.680 161.550 95.970 161.595 ;
        RECT 97.540 161.550 97.830 161.595 ;
        RECT 95.680 161.410 97.830 161.550 ;
        RECT 114.180 161.550 114.320 161.705 ;
        RECT 115.470 161.690 115.790 161.750 ;
        RECT 116.865 161.705 117.155 161.750 ;
        RECT 123.765 161.890 124.055 161.935 ;
        RECT 124.210 161.890 124.530 161.950 ;
        RECT 123.765 161.750 124.530 161.890 ;
        RECT 123.765 161.705 124.055 161.750 ;
        RECT 124.210 161.690 124.530 161.750 ;
        RECT 123.290 161.550 123.610 161.610 ;
        RECT 114.180 161.410 123.610 161.550 ;
        RECT 95.680 161.365 95.970 161.410 ;
        RECT 97.540 161.365 97.830 161.410 ;
        RECT 93.360 161.210 93.650 161.255 ;
        RECT 95.680 161.210 95.895 161.365 ;
        RECT 123.290 161.350 123.610 161.410 ;
        RECT 93.360 161.070 95.895 161.210 ;
        RECT 93.360 161.025 93.650 161.070 ;
        RECT 96.610 161.010 96.930 161.270 ;
        RECT 99.845 161.210 100.135 161.255 ;
        RECT 101.210 161.210 101.530 161.270 ;
        RECT 99.845 161.070 101.530 161.210 ;
        RECT 99.845 161.025 100.135 161.070 ;
        RECT 101.210 161.010 101.530 161.070 ;
        RECT 102.145 161.025 102.435 161.255 ;
        RECT 105.825 161.210 106.115 161.255 ;
        RECT 106.730 161.210 107.050 161.270 ;
        RECT 105.825 161.070 107.050 161.210 ;
        RECT 105.825 161.025 106.115 161.070 ;
        RECT 83.270 160.730 88.100 160.870 ;
        RECT 90.170 160.870 90.490 160.930 ;
        RECT 98.465 160.870 98.755 160.915 ;
        RECT 90.170 160.730 98.755 160.870 ;
        RECT 83.270 160.670 83.590 160.730 ;
        RECT 90.170 160.670 90.490 160.730 ;
        RECT 98.465 160.685 98.755 160.730 ;
        RECT 93.360 160.530 93.650 160.575 ;
        RECT 96.140 160.530 96.430 160.575 ;
        RECT 98.000 160.530 98.290 160.575 ;
        RECT 81.520 160.390 88.560 160.530 ;
        RECT 31.290 160.330 31.610 160.390 ;
        RECT 48.770 160.330 49.090 160.390 ;
        RECT 54.305 160.345 54.595 160.390 ;
        RECT 30.370 160.190 30.690 160.250 ;
        RECT 18.195 160.050 30.690 160.190 ;
        RECT 18.195 160.005 18.485 160.050 ;
        RECT 21.630 159.990 21.950 160.050 ;
        RECT 30.370 159.990 30.690 160.050 ;
        RECT 55.670 160.190 55.990 160.250 ;
        RECT 57.985 160.190 58.275 160.235 ;
        RECT 55.670 160.050 58.275 160.190 ;
        RECT 55.670 159.990 55.990 160.050 ;
        RECT 57.985 160.005 58.275 160.050 ;
        RECT 65.330 159.990 65.650 160.250 ;
        RECT 66.250 160.190 66.570 160.250 ;
        RECT 67.260 160.235 67.400 160.390 ;
        RECT 72.230 160.330 72.550 160.390 ;
        RECT 67.185 160.190 67.475 160.235 ;
        RECT 66.250 160.050 67.475 160.190 ;
        RECT 66.250 159.990 66.570 160.050 ;
        RECT 67.185 160.005 67.475 160.050 ;
        RECT 69.470 159.990 69.790 160.250 ;
        RECT 71.325 160.190 71.615 160.235 ;
        RECT 74.070 160.190 74.390 160.250 ;
        RECT 71.325 160.050 74.390 160.190 ;
        RECT 71.325 160.005 71.615 160.050 ;
        RECT 74.070 159.990 74.390 160.050 ;
        RECT 80.970 159.990 81.290 160.250 ;
        RECT 87.425 160.190 87.715 160.235 ;
        RECT 87.870 160.190 88.190 160.250 ;
        RECT 87.425 160.050 88.190 160.190 ;
        RECT 88.420 160.190 88.560 160.390 ;
        RECT 93.360 160.390 98.290 160.530 ;
        RECT 93.360 160.345 93.650 160.390 ;
        RECT 96.140 160.345 96.430 160.390 ;
        RECT 98.000 160.345 98.290 160.390 ;
        RECT 95.690 160.190 96.010 160.250 ;
        RECT 102.220 160.190 102.360 161.025 ;
        RECT 106.730 161.010 107.050 161.070 ;
        RECT 107.205 161.210 107.495 161.255 ;
        RECT 108.110 161.210 108.430 161.270 ;
        RECT 109.490 161.210 109.810 161.270 ;
        RECT 107.205 161.070 109.810 161.210 ;
        RECT 107.205 161.025 107.495 161.070 ;
        RECT 108.110 161.010 108.430 161.070 ;
        RECT 109.490 161.010 109.810 161.070 ;
        RECT 110.870 161.210 111.190 161.270 ;
        RECT 112.265 161.210 112.555 161.255 ;
        RECT 116.405 161.210 116.695 161.255 ;
        RECT 110.870 161.070 116.695 161.210 ;
        RECT 110.870 161.010 111.190 161.070 ;
        RECT 112.265 161.025 112.555 161.070 ;
        RECT 116.405 161.025 116.695 161.070 ;
        RECT 122.385 161.210 122.675 161.255 ;
        RECT 122.845 161.210 123.135 161.255 ;
        RECT 122.385 161.070 123.135 161.210 ;
        RECT 122.385 161.025 122.675 161.070 ;
        RECT 122.845 161.025 123.135 161.070 ;
        RECT 111.345 160.870 111.635 160.915 ;
        RECT 112.710 160.870 113.030 160.930 ;
        RECT 115.485 160.870 115.775 160.915 ;
        RECT 111.345 160.730 115.775 160.870 ;
        RECT 111.345 160.685 111.635 160.730 ;
        RECT 112.710 160.670 113.030 160.730 ;
        RECT 115.485 160.685 115.775 160.730 ;
        RECT 119.165 160.685 119.455 160.915 ;
        RECT 118.705 160.530 118.995 160.575 ;
        RECT 119.240 160.530 119.380 160.685 ;
        RECT 118.705 160.390 119.380 160.530 ;
        RECT 118.705 160.345 118.995 160.390 ;
        RECT 88.420 160.050 102.360 160.190 ;
        RECT 102.605 160.190 102.895 160.235 ;
        RECT 105.350 160.190 105.670 160.250 ;
        RECT 102.605 160.050 105.670 160.190 ;
        RECT 87.425 160.005 87.715 160.050 ;
        RECT 87.870 159.990 88.190 160.050 ;
        RECT 95.690 159.990 96.010 160.050 ;
        RECT 102.605 160.005 102.895 160.050 ;
        RECT 105.350 159.990 105.670 160.050 ;
        RECT 17.965 159.170 18.255 159.215 ;
        RECT 18.870 159.170 19.190 159.230 ;
        RECT 17.965 159.030 19.190 159.170 ;
        RECT 17.965 158.985 18.255 159.030 ;
        RECT 18.870 158.970 19.190 159.030 ;
        RECT 25.770 158.970 26.090 159.230 ;
        RECT 32.225 159.170 32.515 159.215 ;
        RECT 34.970 159.170 35.290 159.230 ;
        RECT 32.225 159.030 35.290 159.170 ;
        RECT 32.225 158.985 32.515 159.030 ;
        RECT 34.970 158.970 35.290 159.030 ;
        RECT 54.750 158.970 55.070 159.230 ;
        RECT 72.230 159.170 72.550 159.230 ;
        RECT 93.405 159.170 93.695 159.215 ;
        RECT 93.850 159.170 94.170 159.230 ;
        RECT 72.230 159.030 93.160 159.170 ;
        RECT 72.230 158.970 72.550 159.030 ;
        RECT 31.290 158.830 31.610 158.890 ;
        RECT 49.230 158.830 49.550 158.890 ;
        RECT 21.260 158.690 31.610 158.830 ;
        RECT 21.260 158.550 21.400 158.690 ;
        RECT 31.290 158.630 31.610 158.690 ;
        RECT 42.880 158.690 49.550 158.830 ;
        RECT 21.170 158.290 21.490 158.550 ;
        RECT 21.630 158.290 21.950 158.550 ;
        RECT 35.445 158.490 35.735 158.535 ;
        RECT 35.890 158.490 36.210 158.550 ;
        RECT 22.870 158.350 32.900 158.490 ;
        RECT 18.425 158.150 18.715 158.195 ;
        RECT 18.870 158.150 19.190 158.210 ;
        RECT 18.425 158.010 19.190 158.150 ;
        RECT 18.425 157.965 18.715 158.010 ;
        RECT 18.870 157.950 19.190 158.010 ;
        RECT 19.330 157.270 19.650 157.530 ;
        RECT 21.630 157.470 21.950 157.530 ;
        RECT 22.105 157.470 22.395 157.515 ;
        RECT 22.870 157.470 23.010 158.350 ;
        RECT 24.865 158.150 25.155 158.195 ;
        RECT 24.020 158.010 25.155 158.150 ;
        RECT 32.760 158.150 32.900 158.350 ;
        RECT 35.445 158.350 36.210 158.490 ;
        RECT 35.445 158.305 35.735 158.350 ;
        RECT 35.890 158.290 36.210 158.350 ;
        RECT 40.950 158.490 41.270 158.550 ;
        RECT 42.880 158.490 43.020 158.690 ;
        RECT 49.230 158.630 49.550 158.690 ;
        RECT 51.990 158.830 52.310 158.890 ;
        RECT 74.070 158.830 74.390 158.890 ;
        RECT 51.990 158.690 74.390 158.830 ;
        RECT 51.990 158.630 52.310 158.690 ;
        RECT 74.070 158.630 74.390 158.690 ;
        RECT 84.620 158.830 84.910 158.875 ;
        RECT 87.400 158.830 87.690 158.875 ;
        RECT 89.260 158.830 89.550 158.875 ;
        RECT 84.620 158.690 89.550 158.830 ;
        RECT 93.020 158.830 93.160 159.030 ;
        RECT 93.405 159.030 94.170 159.170 ;
        RECT 93.405 158.985 93.695 159.030 ;
        RECT 93.850 158.970 94.170 159.030 ;
        RECT 96.165 159.170 96.455 159.215 ;
        RECT 96.610 159.170 96.930 159.230 ;
        RECT 96.165 159.030 96.930 159.170 ;
        RECT 96.165 158.985 96.455 159.030 ;
        RECT 96.610 158.970 96.930 159.030 ;
        RECT 106.285 159.170 106.575 159.215 ;
        RECT 109.950 159.170 110.270 159.230 ;
        RECT 106.285 159.030 110.270 159.170 ;
        RECT 106.285 158.985 106.575 159.030 ;
        RECT 109.950 158.970 110.270 159.030 ;
        RECT 98.910 158.830 99.230 158.890 ;
        RECT 105.810 158.830 106.130 158.890 ;
        RECT 93.020 158.690 106.130 158.830 ;
        RECT 84.620 158.645 84.910 158.690 ;
        RECT 87.400 158.645 87.690 158.690 ;
        RECT 89.260 158.645 89.550 158.690 ;
        RECT 98.910 158.630 99.230 158.690 ;
        RECT 105.810 158.630 106.130 158.690 ;
        RECT 65.330 158.490 65.650 158.550 ;
        RECT 80.510 158.535 80.830 158.550 ;
        RECT 80.510 158.490 81.045 158.535 ;
        RECT 40.950 158.350 43.020 158.490 ;
        RECT 40.950 158.290 41.270 158.350 ;
        RECT 42.330 158.150 42.650 158.210 ;
        RECT 42.880 158.195 43.020 158.350 ;
        RECT 44.260 158.350 78.900 158.490 ;
        RECT 32.760 158.010 42.650 158.150 ;
        RECT 24.020 157.515 24.160 158.010 ;
        RECT 24.865 157.965 25.155 158.010 ;
        RECT 42.330 157.950 42.650 158.010 ;
        RECT 42.805 157.965 43.095 158.195 ;
        RECT 43.710 157.950 44.030 158.210 ;
        RECT 44.260 158.195 44.400 158.350 ;
        RECT 48.400 158.210 48.540 158.350 ;
        RECT 44.185 157.965 44.475 158.195 ;
        RECT 44.645 158.150 44.935 158.195 ;
        RECT 44.645 158.010 45.320 158.150 ;
        RECT 44.645 157.965 44.935 158.010 ;
        RECT 41.870 157.810 42.190 157.870 ;
        RECT 44.260 157.810 44.400 157.965 ;
        RECT 41.870 157.670 44.400 157.810 ;
        RECT 45.180 157.810 45.320 158.010 ;
        RECT 47.865 157.965 48.155 158.195 ;
        RECT 47.940 157.810 48.080 157.965 ;
        RECT 48.310 157.950 48.630 158.210 ;
        RECT 48.770 157.950 49.090 158.210 ;
        RECT 49.230 158.150 49.550 158.210 ;
        RECT 49.705 158.150 49.995 158.195 ;
        RECT 49.230 158.010 51.760 158.150 ;
        RECT 49.230 157.950 49.550 158.010 ;
        RECT 49.705 157.965 49.995 158.010 ;
        RECT 51.620 157.810 51.760 158.010 ;
        RECT 51.990 157.950 52.310 158.210 ;
        RECT 52.540 158.195 52.680 158.350 ;
        RECT 65.330 158.290 65.650 158.350 ;
        RECT 52.465 157.965 52.755 158.195 ;
        RECT 52.910 157.950 53.230 158.210 ;
        RECT 53.845 157.965 54.135 158.195 ;
        RECT 53.920 157.810 54.060 157.965 ;
        RECT 55.670 157.950 55.990 158.210 ;
        RECT 57.050 158.150 57.370 158.210 ;
        RECT 62.585 158.150 62.875 158.195 ;
        RECT 63.490 158.150 63.810 158.210 ;
        RECT 57.050 158.010 63.810 158.150 ;
        RECT 57.050 157.950 57.370 158.010 ;
        RECT 62.585 157.965 62.875 158.010 ;
        RECT 63.490 157.950 63.810 158.010 ;
        RECT 63.965 158.150 64.255 158.195 ;
        RECT 64.410 158.150 64.730 158.210 ;
        RECT 63.965 158.010 64.730 158.150 ;
        RECT 63.965 157.965 64.255 158.010 ;
        RECT 64.410 157.950 64.730 158.010 ;
        RECT 68.565 158.150 68.855 158.195 ;
        RECT 70.405 158.150 70.695 158.195 ;
        RECT 70.850 158.150 71.170 158.210 ;
        RECT 68.565 158.010 71.170 158.150 ;
        RECT 68.565 157.965 68.855 158.010 ;
        RECT 70.405 157.965 70.695 158.010 ;
        RECT 70.850 157.950 71.170 158.010 ;
        RECT 72.245 157.965 72.535 158.195 ;
        RECT 72.320 157.810 72.460 157.965 ;
        RECT 73.150 157.950 73.470 158.210 ;
        RECT 73.700 158.195 73.840 158.350 ;
        RECT 78.760 158.210 78.900 158.350 ;
        RECT 79.220 158.350 81.265 158.490 ;
        RECT 73.625 157.965 73.915 158.195 ;
        RECT 74.070 158.150 74.390 158.210 ;
        RECT 78.210 158.150 78.530 158.210 ;
        RECT 74.070 158.010 78.530 158.150 ;
        RECT 74.070 157.950 74.390 158.010 ;
        RECT 78.210 157.950 78.530 158.010 ;
        RECT 78.670 157.950 78.990 158.210 ;
        RECT 79.220 158.195 79.360 158.350 ;
        RECT 80.510 158.305 81.045 158.350 ;
        RECT 80.510 158.290 80.830 158.305 ;
        RECT 87.870 158.290 88.190 158.550 ;
        RECT 79.145 157.965 79.435 158.195 ;
        RECT 80.065 158.150 80.355 158.195 ;
        RECT 83.730 158.150 84.050 158.210 ;
        RECT 80.065 158.010 84.050 158.150 ;
        RECT 80.065 157.965 80.355 158.010 ;
        RECT 74.990 157.810 75.310 157.870 ;
        RECT 80.140 157.810 80.280 157.965 ;
        RECT 83.730 157.950 84.050 158.010 ;
        RECT 84.620 158.150 84.910 158.195 ;
        RECT 89.725 158.150 90.015 158.195 ;
        RECT 90.170 158.150 90.490 158.210 ;
        RECT 84.620 158.010 87.155 158.150 ;
        RECT 84.620 157.965 84.910 158.010 ;
        RECT 45.180 157.670 51.300 157.810 ;
        RECT 51.620 157.670 80.280 157.810 ;
        RECT 80.970 157.810 81.290 157.870 ;
        RECT 86.940 157.855 87.155 158.010 ;
        RECT 89.725 158.010 90.490 158.150 ;
        RECT 89.725 157.965 90.015 158.010 ;
        RECT 90.170 157.950 90.490 158.010 ;
        RECT 93.850 158.150 94.170 158.210 ;
        RECT 95.690 158.150 96.010 158.210 ;
        RECT 93.850 158.010 96.010 158.150 ;
        RECT 93.850 157.950 94.170 158.010 ;
        RECT 95.690 157.950 96.010 158.010 ;
        RECT 97.070 157.950 97.390 158.210 ;
        RECT 105.350 157.950 105.670 158.210 ;
        RECT 121.450 157.950 121.770 158.210 ;
        RECT 82.760 157.810 83.050 157.855 ;
        RECT 86.020 157.810 86.310 157.855 ;
        RECT 80.970 157.670 86.310 157.810 ;
        RECT 41.870 157.610 42.190 157.670 ;
        RECT 45.180 157.530 45.320 157.670 ;
        RECT 21.630 157.330 23.010 157.470 ;
        RECT 21.630 157.270 21.950 157.330 ;
        RECT 22.105 157.285 22.395 157.330 ;
        RECT 23.945 157.285 24.235 157.515 ;
        RECT 42.790 157.470 43.110 157.530 ;
        RECT 45.090 157.470 45.410 157.530 ;
        RECT 42.790 157.330 45.410 157.470 ;
        RECT 42.790 157.270 43.110 157.330 ;
        RECT 45.090 157.270 45.410 157.330 ;
        RECT 45.550 157.470 45.870 157.530 ;
        RECT 46.025 157.470 46.315 157.515 ;
        RECT 45.550 157.330 46.315 157.470 ;
        RECT 45.550 157.270 45.870 157.330 ;
        RECT 46.025 157.285 46.315 157.330 ;
        RECT 46.485 157.470 46.775 157.515 ;
        RECT 47.390 157.470 47.710 157.530 ;
        RECT 46.485 157.330 47.710 157.470 ;
        RECT 46.485 157.285 46.775 157.330 ;
        RECT 47.390 157.270 47.710 157.330 ;
        RECT 50.150 157.470 50.470 157.530 ;
        RECT 50.625 157.470 50.915 157.515 ;
        RECT 50.150 157.330 50.915 157.470 ;
        RECT 51.160 157.470 51.300 157.670 ;
        RECT 51.990 157.470 52.310 157.530 ;
        RECT 69.560 157.515 69.700 157.670 ;
        RECT 74.990 157.610 75.310 157.670 ;
        RECT 80.970 157.610 81.290 157.670 ;
        RECT 82.760 157.625 83.050 157.670 ;
        RECT 86.020 157.625 86.310 157.670 ;
        RECT 86.940 157.810 87.230 157.855 ;
        RECT 88.800 157.810 89.090 157.855 ;
        RECT 86.940 157.670 89.090 157.810 ;
        RECT 86.940 157.625 87.230 157.670 ;
        RECT 88.800 157.625 89.090 157.670 ;
        RECT 120.085 157.810 120.375 157.855 ;
        RECT 120.530 157.810 120.850 157.870 ;
        RECT 120.085 157.670 120.850 157.810 ;
        RECT 120.085 157.625 120.375 157.670 ;
        RECT 120.530 157.610 120.850 157.670 ;
        RECT 51.160 157.330 52.310 157.470 ;
        RECT 50.150 157.270 50.470 157.330 ;
        RECT 50.625 157.285 50.915 157.330 ;
        RECT 51.990 157.270 52.310 157.330 ;
        RECT 69.485 157.285 69.775 157.515 ;
        RECT 71.325 157.470 71.615 157.515 ;
        RECT 72.230 157.470 72.550 157.530 ;
        RECT 71.325 157.330 72.550 157.470 ;
        RECT 71.325 157.285 71.615 157.330 ;
        RECT 72.230 157.270 72.550 157.330 ;
        RECT 75.465 157.470 75.755 157.515 ;
        RECT 75.910 157.470 76.230 157.530 ;
        RECT 75.465 157.330 76.230 157.470 ;
        RECT 75.465 157.285 75.755 157.330 ;
        RECT 75.910 157.270 76.230 157.330 ;
        RECT 76.830 157.270 77.150 157.530 ;
        RECT 16.815 156.450 17.105 156.495 ;
        RECT 21.630 156.450 21.950 156.510 ;
        RECT 16.815 156.310 21.950 156.450 ;
        RECT 16.815 156.265 17.105 156.310 ;
        RECT 21.630 156.250 21.950 156.310 ;
        RECT 26.245 156.265 26.535 156.495 ;
        RECT 18.820 156.110 19.110 156.155 ;
        RECT 19.330 156.110 19.650 156.170 ;
        RECT 22.080 156.110 22.370 156.155 ;
        RECT 18.820 155.970 22.370 156.110 ;
        RECT 18.820 155.925 19.110 155.970 ;
        RECT 19.330 155.910 19.650 155.970 ;
        RECT 22.080 155.925 22.370 155.970 ;
        RECT 23.000 156.110 23.290 156.155 ;
        RECT 24.860 156.110 25.150 156.155 ;
        RECT 23.000 155.970 25.150 156.110 ;
        RECT 23.000 155.925 23.290 155.970 ;
        RECT 24.860 155.925 25.150 155.970 ;
        RECT 20.680 155.770 20.970 155.815 ;
        RECT 23.000 155.770 23.215 155.925 ;
        RECT 20.680 155.630 23.215 155.770 ;
        RECT 23.945 155.770 24.235 155.815 ;
        RECT 26.320 155.770 26.460 156.265 ;
        RECT 26.690 156.250 27.010 156.510 ;
        RECT 34.510 156.450 34.830 156.510 ;
        RECT 35.445 156.450 35.735 156.495 ;
        RECT 63.965 156.450 64.255 156.495 ;
        RECT 34.510 156.310 35.735 156.450 ;
        RECT 34.510 156.250 34.830 156.310 ;
        RECT 35.445 156.265 35.735 156.310 ;
        RECT 36.670 156.310 48.540 156.450 ;
        RECT 26.780 156.110 26.920 156.250 ;
        RECT 26.780 155.970 32.440 156.110 ;
        RECT 32.300 155.815 32.440 155.970 ;
        RECT 27.165 155.770 27.455 155.815 ;
        RECT 23.945 155.630 26.460 155.770 ;
        RECT 26.780 155.630 27.455 155.770 ;
        RECT 20.680 155.585 20.970 155.630 ;
        RECT 23.945 155.585 24.235 155.630 ;
        RECT 26.780 155.490 26.920 155.630 ;
        RECT 27.165 155.585 27.455 155.630 ;
        RECT 32.225 155.585 32.515 155.815 ;
        RECT 25.770 155.230 26.090 155.490 ;
        RECT 26.690 155.230 27.010 155.490 ;
        RECT 20.680 155.090 20.970 155.135 ;
        RECT 23.460 155.090 23.750 155.135 ;
        RECT 25.320 155.090 25.610 155.135 ;
        RECT 20.680 154.950 25.610 155.090 ;
        RECT 32.300 155.090 32.440 155.585 ;
        RECT 34.050 155.430 34.370 155.490 ;
        RECT 36.670 155.430 36.810 156.310 ;
        RECT 42.790 156.110 43.110 156.170 ;
        RECT 41.500 155.970 43.110 156.110 ;
        RECT 41.500 155.815 41.640 155.970 ;
        RECT 42.790 155.910 43.110 155.970 ;
        RECT 43.800 155.970 45.780 156.110 ;
        RECT 41.425 155.585 41.715 155.815 ;
        RECT 41.870 155.570 42.190 155.830 ;
        RECT 42.330 155.570 42.650 155.830 ;
        RECT 43.250 155.570 43.570 155.830 ;
        RECT 34.050 155.290 36.810 155.430 ;
        RECT 41.960 155.430 42.100 155.570 ;
        RECT 43.800 155.430 43.940 155.970 ;
        RECT 45.090 155.815 45.410 155.830 ;
        RECT 45.640 155.815 45.780 155.970 ;
        RECT 48.400 155.815 48.540 156.310 ;
        RECT 59.440 156.310 64.255 156.450 ;
        RECT 55.620 156.110 55.910 156.155 ;
        RECT 58.880 156.110 59.170 156.155 ;
        RECT 59.440 156.110 59.580 156.310 ;
        RECT 63.965 156.265 64.255 156.310 ;
        RECT 64.410 156.450 64.730 156.510 ;
        RECT 64.410 156.310 116.620 156.450 ;
        RECT 64.410 156.250 64.730 156.310 ;
        RECT 55.620 155.970 59.580 156.110 ;
        RECT 59.800 156.110 60.090 156.155 ;
        RECT 61.660 156.110 61.950 156.155 ;
        RECT 69.470 156.110 69.790 156.170 ;
        RECT 59.800 155.970 61.950 156.110 ;
        RECT 55.620 155.925 55.910 155.970 ;
        RECT 58.880 155.925 59.170 155.970 ;
        RECT 59.800 155.925 60.090 155.970 ;
        RECT 61.660 155.925 61.950 155.970 ;
        RECT 62.200 155.970 69.790 156.110 ;
        RECT 44.875 155.585 45.410 155.815 ;
        RECT 45.565 155.585 45.855 155.815 ;
        RECT 46.130 155.770 46.420 155.815 ;
        RECT 46.945 155.800 47.235 155.815 ;
        RECT 47.435 155.800 47.725 155.815 ;
        RECT 46.945 155.770 47.725 155.800 ;
        RECT 46.130 155.630 46.700 155.770 ;
        RECT 46.130 155.585 46.420 155.630 ;
        RECT 45.090 155.570 45.410 155.585 ;
        RECT 41.960 155.290 43.940 155.430 ;
        RECT 34.050 155.230 34.370 155.290 ;
        RECT 46.560 155.090 46.700 155.630 ;
        RECT 46.945 155.660 48.080 155.770 ;
        RECT 46.945 155.585 47.235 155.660 ;
        RECT 47.435 155.630 48.080 155.660 ;
        RECT 47.435 155.585 47.725 155.630 ;
        RECT 47.940 155.430 48.080 155.630 ;
        RECT 48.325 155.585 48.615 155.815 ;
        RECT 48.770 155.570 49.090 155.830 ;
        RECT 49.245 155.770 49.535 155.815 ;
        RECT 51.990 155.770 52.310 155.830 ;
        RECT 49.245 155.630 52.310 155.770 ;
        RECT 49.245 155.585 49.535 155.630 ;
        RECT 51.990 155.570 52.310 155.630 ;
        RECT 57.480 155.770 57.770 155.815 ;
        RECT 59.800 155.770 60.015 155.925 ;
        RECT 57.480 155.630 60.015 155.770 ;
        RECT 60.270 155.770 60.590 155.830 ;
        RECT 62.200 155.770 62.340 155.970 ;
        RECT 69.470 155.910 69.790 155.970 ;
        RECT 74.990 156.110 75.310 156.170 ;
        RECT 78.670 156.110 78.990 156.170 ;
        RECT 106.730 156.110 107.050 156.170 ;
        RECT 74.990 155.970 76.140 156.110 ;
        RECT 74.990 155.910 75.310 155.970 ;
        RECT 60.270 155.630 62.340 155.770 ;
        RECT 57.480 155.585 57.770 155.630 ;
        RECT 60.270 155.570 60.590 155.630 ;
        RECT 63.490 155.570 63.810 155.830 ;
        RECT 76.000 155.815 76.140 155.970 ;
        RECT 77.380 155.970 82.580 156.110 ;
        RECT 75.925 155.585 76.215 155.815 ;
        RECT 76.370 155.770 76.690 155.830 ;
        RECT 77.380 155.815 77.520 155.970 ;
        RECT 78.670 155.910 78.990 155.970 ;
        RECT 76.845 155.770 77.135 155.815 ;
        RECT 76.370 155.630 77.135 155.770 ;
        RECT 76.370 155.570 76.690 155.630 ;
        RECT 76.845 155.585 77.135 155.630 ;
        RECT 77.305 155.585 77.595 155.815 ;
        RECT 77.765 155.770 78.055 155.815 ;
        RECT 78.210 155.770 78.530 155.830 ;
        RECT 82.440 155.815 82.580 155.970 ;
        RECT 99.460 155.970 112.940 156.110 ;
        RECT 99.460 155.830 99.600 155.970 ;
        RECT 81.905 155.770 82.195 155.815 ;
        RECT 77.765 155.630 82.195 155.770 ;
        RECT 77.765 155.585 78.055 155.630 ;
        RECT 78.210 155.570 78.530 155.630 ;
        RECT 81.905 155.585 82.195 155.630 ;
        RECT 82.365 155.585 82.655 155.815 ;
        RECT 82.825 155.770 83.115 155.815 ;
        RECT 83.270 155.770 83.590 155.830 ;
        RECT 82.825 155.630 83.590 155.770 ;
        RECT 82.825 155.585 83.115 155.630 ;
        RECT 83.270 155.570 83.590 155.630 ;
        RECT 83.730 155.570 84.050 155.830 ;
        RECT 98.910 155.570 99.230 155.830 ;
        RECT 99.370 155.570 99.690 155.830 ;
        RECT 99.845 155.770 100.135 155.815 ;
        RECT 100.290 155.770 100.610 155.830 ;
        RECT 99.845 155.630 100.610 155.770 ;
        RECT 99.845 155.585 100.135 155.630 ;
        RECT 100.290 155.570 100.610 155.630 ;
        RECT 100.765 155.770 101.055 155.815 ;
        RECT 103.525 155.770 103.815 155.815 ;
        RECT 100.765 155.630 103.815 155.770 ;
        RECT 100.765 155.585 101.055 155.630 ;
        RECT 47.940 155.290 49.460 155.430 ;
        RECT 49.320 155.150 49.460 155.290 ;
        RECT 60.730 155.230 61.050 155.490 ;
        RECT 62.585 155.430 62.875 155.475 ;
        RECT 63.950 155.430 64.270 155.490 ;
        RECT 62.585 155.290 64.270 155.430 ;
        RECT 62.585 155.245 62.875 155.290 ;
        RECT 63.950 155.230 64.270 155.290 ;
        RECT 66.710 155.230 67.030 155.490 ;
        RECT 32.300 154.950 46.700 155.090 ;
        RECT 20.680 154.905 20.970 154.950 ;
        RECT 23.460 154.905 23.750 154.950 ;
        RECT 25.320 154.905 25.610 154.950 ;
        RECT 49.230 154.890 49.550 155.150 ;
        RECT 57.480 155.090 57.770 155.135 ;
        RECT 60.260 155.090 60.550 155.135 ;
        RECT 62.120 155.090 62.410 155.135 ;
        RECT 57.480 154.950 62.410 155.090 ;
        RECT 57.480 154.905 57.770 154.950 ;
        RECT 60.260 154.905 60.550 154.950 ;
        RECT 62.120 154.905 62.410 154.950 ;
        RECT 78.670 155.090 78.990 155.150 ;
        RECT 79.145 155.090 79.435 155.135 ;
        RECT 78.670 154.950 79.435 155.090 ;
        RECT 78.670 154.890 78.990 154.950 ;
        RECT 79.145 154.905 79.435 154.950 ;
        RECT 80.525 155.090 80.815 155.135 ;
        RECT 82.810 155.090 83.130 155.150 ;
        RECT 80.525 154.950 83.130 155.090 ;
        RECT 80.525 154.905 80.815 154.950 ;
        RECT 82.810 154.890 83.130 154.950 ;
        RECT 97.160 154.950 100.520 155.090 ;
        RECT 40.030 154.550 40.350 154.810 ;
        RECT 43.710 154.550 44.030 154.810 ;
        RECT 50.610 154.550 50.930 154.810 ;
        RECT 53.830 154.795 54.150 154.810 ;
        RECT 53.615 154.565 54.150 154.795 ;
        RECT 53.830 154.550 54.150 154.565 ;
        RECT 67.170 154.750 67.490 154.810 ;
        RECT 72.230 154.750 72.550 154.810 ;
        RECT 97.160 154.750 97.300 154.950 ;
        RECT 67.170 154.610 97.300 154.750 ;
        RECT 67.170 154.550 67.490 154.610 ;
        RECT 72.230 154.550 72.550 154.610 ;
        RECT 97.530 154.550 97.850 154.810 ;
        RECT 100.380 154.750 100.520 154.950 ;
        RECT 101.300 154.750 101.440 155.630 ;
        RECT 103.525 155.585 103.815 155.630 ;
        RECT 103.600 155.430 103.740 155.585 ;
        RECT 104.430 155.570 104.750 155.830 ;
        RECT 104.980 155.815 105.120 155.970 ;
        RECT 106.730 155.910 107.050 155.970 ;
        RECT 104.905 155.585 105.195 155.815 ;
        RECT 105.365 155.770 105.655 155.815 ;
        RECT 105.810 155.770 106.130 155.830 ;
        RECT 105.365 155.630 106.130 155.770 ;
        RECT 105.365 155.585 105.655 155.630 ;
        RECT 105.810 155.570 106.130 155.630 ;
        RECT 107.205 155.585 107.495 155.815 ;
        RECT 107.280 155.430 107.420 155.585 ;
        RECT 108.110 155.570 108.430 155.830 ;
        RECT 108.660 155.815 108.800 155.970 ;
        RECT 108.585 155.585 108.875 155.815 ;
        RECT 109.045 155.770 109.335 155.815 ;
        RECT 111.330 155.770 111.650 155.830 ;
        RECT 112.800 155.815 112.940 155.970 ;
        RECT 112.265 155.770 112.555 155.815 ;
        RECT 109.045 155.630 112.555 155.770 ;
        RECT 109.045 155.585 109.335 155.630 ;
        RECT 111.330 155.570 111.650 155.630 ;
        RECT 112.265 155.585 112.555 155.630 ;
        RECT 112.725 155.585 113.015 155.815 ;
        RECT 113.170 155.570 113.490 155.830 ;
        RECT 116.480 155.815 116.620 156.310 ;
        RECT 114.105 155.585 114.395 155.815 ;
        RECT 116.405 155.770 116.695 155.815 ;
        RECT 121.450 155.770 121.770 155.830 ;
        RECT 116.405 155.630 121.770 155.770 ;
        RECT 116.405 155.585 116.695 155.630 ;
        RECT 114.180 155.430 114.320 155.585 ;
        RECT 121.450 155.570 121.770 155.630 ;
        RECT 103.600 155.290 107.420 155.430 ;
        RECT 107.280 155.090 107.420 155.290 ;
        RECT 112.340 155.290 114.320 155.430 ;
        RECT 116.850 155.430 117.170 155.490 ;
        RECT 117.325 155.430 117.615 155.475 ;
        RECT 116.850 155.290 117.615 155.430 ;
        RECT 112.340 155.150 112.480 155.290 ;
        RECT 116.850 155.230 117.170 155.290 ;
        RECT 117.325 155.245 117.615 155.290 ;
        RECT 108.570 155.090 108.890 155.150 ;
        RECT 112.250 155.090 112.570 155.150 ;
        RECT 107.280 154.950 112.570 155.090 ;
        RECT 108.570 154.890 108.890 154.950 ;
        RECT 112.250 154.890 112.570 154.950 ;
        RECT 100.380 154.610 101.440 154.750 ;
        RECT 104.430 154.750 104.750 154.810 ;
        RECT 106.745 154.750 107.035 154.795 ;
        RECT 104.430 154.610 107.035 154.750 ;
        RECT 104.430 154.550 104.750 154.610 ;
        RECT 106.745 154.565 107.035 154.610 ;
        RECT 110.410 154.550 110.730 154.810 ;
        RECT 110.870 154.550 111.190 154.810 ;
        RECT 23.945 153.730 24.235 153.775 ;
        RECT 26.690 153.730 27.010 153.790 ;
        RECT 23.945 153.590 27.010 153.730 ;
        RECT 23.945 153.545 24.235 153.590 ;
        RECT 26.690 153.530 27.010 153.590 ;
        RECT 42.790 153.730 43.110 153.790 ;
        RECT 66.250 153.730 66.570 153.790 ;
        RECT 42.790 153.590 66.570 153.730 ;
        RECT 42.790 153.530 43.110 153.590 ;
        RECT 66.250 153.530 66.570 153.590 ;
        RECT 69.470 153.730 69.790 153.790 ;
        RECT 99.370 153.730 99.690 153.790 ;
        RECT 120.530 153.730 120.850 153.790 ;
        RECT 69.470 153.590 99.690 153.730 ;
        RECT 69.470 153.530 69.790 153.590 ;
        RECT 99.370 153.530 99.690 153.590 ;
        RECT 99.920 153.590 120.850 153.730 ;
        RECT 31.290 153.390 31.610 153.450 ;
        RECT 39.570 153.390 39.890 153.450 ;
        RECT 42.330 153.390 42.650 153.450 ;
        RECT 60.270 153.390 60.590 153.450 ;
        RECT 31.290 153.250 36.580 153.390 ;
        RECT 31.290 153.190 31.610 153.250 ;
        RECT 21.170 152.850 21.490 153.110 ;
        RECT 21.630 152.850 21.950 153.110 ;
        RECT 30.370 153.050 30.690 153.110 ;
        RECT 36.440 153.095 36.580 153.250 ;
        RECT 39.570 153.250 60.590 153.390 ;
        RECT 39.570 153.190 39.890 153.250 ;
        RECT 42.330 153.190 42.650 153.250 ;
        RECT 60.270 153.190 60.590 153.250 ;
        RECT 62.540 153.390 62.830 153.435 ;
        RECT 65.320 153.390 65.610 153.435 ;
        RECT 67.180 153.390 67.470 153.435 ;
        RECT 62.540 153.250 67.470 153.390 ;
        RECT 62.540 153.205 62.830 153.250 ;
        RECT 65.320 153.205 65.610 153.250 ;
        RECT 67.180 153.205 67.470 153.250 ;
        RECT 67.630 153.390 67.950 153.450 ;
        RECT 70.850 153.390 71.170 153.450 ;
        RECT 93.850 153.390 94.170 153.450 ;
        RECT 95.690 153.390 96.010 153.450 ;
        RECT 99.920 153.390 100.060 153.590 ;
        RECT 111.330 153.390 111.650 153.450 ;
        RECT 67.630 153.250 75.220 153.390 ;
        RECT 67.630 153.190 67.950 153.250 ;
        RECT 70.850 153.190 71.170 153.250 ;
        RECT 30.370 152.910 34.280 153.050 ;
        RECT 30.370 152.850 30.690 152.910 ;
        RECT 25.310 152.710 25.630 152.770 ;
        RECT 30.845 152.710 31.135 152.755 ;
        RECT 25.310 152.570 31.135 152.710 ;
        RECT 25.310 152.510 25.630 152.570 ;
        RECT 30.845 152.525 31.135 152.570 ;
        RECT 32.225 152.710 32.515 152.755 ;
        RECT 32.225 152.570 33.820 152.710 ;
        RECT 32.225 152.525 32.515 152.570 ;
        RECT 22.105 152.030 22.395 152.075 ;
        RECT 22.550 152.030 22.870 152.090 ;
        RECT 22.105 151.890 22.870 152.030 ;
        RECT 22.105 151.845 22.395 151.890 ;
        RECT 22.550 151.830 22.870 151.890 ;
        RECT 31.290 151.830 31.610 152.090 ;
        RECT 33.130 151.830 33.450 152.090 ;
        RECT 33.680 152.075 33.820 152.570 ;
        RECT 34.140 152.370 34.280 152.910 ;
        RECT 36.365 152.865 36.655 153.095 ;
        RECT 42.790 153.050 43.110 153.110 ;
        RECT 39.200 152.910 43.110 153.050 ;
        RECT 34.510 152.710 34.830 152.770 ;
        RECT 35.445 152.710 35.735 152.755 ;
        RECT 34.510 152.570 35.735 152.710 ;
        RECT 34.510 152.510 34.830 152.570 ;
        RECT 35.445 152.525 35.735 152.570 ;
        RECT 35.905 152.710 36.195 152.755 ;
        RECT 37.270 152.710 37.590 152.770 ;
        RECT 39.200 152.755 39.340 152.910 ;
        RECT 42.790 152.850 43.110 152.910 ;
        RECT 63.950 153.050 64.270 153.110 ;
        RECT 63.950 152.910 65.560 153.050 ;
        RECT 63.950 152.850 64.270 152.910 ;
        RECT 35.905 152.570 37.590 152.710 ;
        RECT 35.905 152.525 36.195 152.570 ;
        RECT 37.270 152.510 37.590 152.570 ;
        RECT 39.125 152.525 39.415 152.755 ;
        RECT 39.570 152.510 39.890 152.770 ;
        RECT 40.045 152.525 40.335 152.755 ;
        RECT 40.965 152.710 41.255 152.755 ;
        RECT 41.870 152.710 42.190 152.770 ;
        RECT 40.965 152.570 42.190 152.710 ;
        RECT 40.965 152.525 41.255 152.570 ;
        RECT 40.120 152.370 40.260 152.525 ;
        RECT 41.870 152.510 42.190 152.570 ;
        RECT 51.530 152.710 51.850 152.770 ;
        RECT 57.050 152.710 57.370 152.770 ;
        RECT 51.530 152.570 57.370 152.710 ;
        RECT 51.530 152.510 51.850 152.570 ;
        RECT 57.050 152.510 57.370 152.570 ;
        RECT 62.540 152.710 62.830 152.755 ;
        RECT 65.420 152.710 65.560 152.910 ;
        RECT 65.790 152.850 66.110 153.110 ;
        RECT 75.080 153.095 75.220 153.250 ;
        RECT 93.850 153.250 100.060 153.390 ;
        RECT 110.500 153.250 111.650 153.390 ;
        RECT 93.850 153.190 94.170 153.250 ;
        RECT 95.690 153.190 96.010 153.250 ;
        RECT 73.625 153.050 73.915 153.095 ;
        RECT 71.860 152.910 73.915 153.050 ;
        RECT 71.860 152.770 72.000 152.910 ;
        RECT 73.625 152.865 73.915 152.910 ;
        RECT 75.005 152.865 75.295 153.095 ;
        RECT 110.500 153.050 110.640 153.250 ;
        RECT 111.330 153.190 111.650 153.250 ;
        RECT 115.470 153.050 115.790 153.110 ;
        RECT 106.820 152.910 110.640 153.050 ;
        RECT 67.645 152.710 67.935 152.755 ;
        RECT 62.540 152.570 65.075 152.710 ;
        RECT 65.420 152.570 67.935 152.710 ;
        RECT 62.540 152.525 62.830 152.570 ;
        RECT 64.860 152.415 65.075 152.570 ;
        RECT 67.645 152.525 67.935 152.570 ;
        RECT 71.325 152.710 71.615 152.755 ;
        RECT 71.770 152.710 72.090 152.770 ;
        RECT 71.325 152.570 72.090 152.710 ;
        RECT 71.325 152.525 71.615 152.570 ;
        RECT 71.770 152.510 72.090 152.570 ;
        RECT 73.165 152.525 73.455 152.755 ;
        RECT 74.070 152.710 74.390 152.770 ;
        RECT 74.545 152.710 74.835 152.755 ;
        RECT 74.070 152.570 74.835 152.710 ;
        RECT 34.140 152.230 40.260 152.370 ;
        RECT 57.525 152.370 57.815 152.415 ;
        RECT 60.680 152.370 60.970 152.415 ;
        RECT 63.940 152.370 64.230 152.415 ;
        RECT 57.525 152.230 64.230 152.370 ;
        RECT 57.525 152.185 57.815 152.230 ;
        RECT 60.680 152.185 60.970 152.230 ;
        RECT 63.940 152.185 64.230 152.230 ;
        RECT 64.860 152.370 65.150 152.415 ;
        RECT 66.720 152.370 67.010 152.415 ;
        RECT 64.860 152.230 67.010 152.370 ;
        RECT 64.860 152.185 65.150 152.230 ;
        RECT 66.720 152.185 67.010 152.230 ;
        RECT 70.390 152.370 70.710 152.430 ;
        RECT 73.240 152.370 73.380 152.525 ;
        RECT 74.070 152.510 74.390 152.570 ;
        RECT 74.545 152.525 74.835 152.570 ;
        RECT 86.490 152.710 86.810 152.770 ;
        RECT 90.645 152.710 90.935 152.755 ;
        RECT 101.210 152.710 101.530 152.770 ;
        RECT 86.490 152.570 101.530 152.710 ;
        RECT 86.490 152.510 86.810 152.570 ;
        RECT 90.645 152.525 90.935 152.570 ;
        RECT 101.210 152.510 101.530 152.570 ;
        RECT 105.810 152.710 106.130 152.770 ;
        RECT 106.820 152.755 106.960 152.910 ;
        RECT 106.745 152.710 107.035 152.755 ;
        RECT 105.810 152.570 107.035 152.710 ;
        RECT 105.810 152.510 106.130 152.570 ;
        RECT 106.745 152.525 107.035 152.570 ;
        RECT 107.190 152.510 107.510 152.770 ;
        RECT 107.650 152.510 107.970 152.770 ;
        RECT 108.570 152.510 108.890 152.770 ;
        RECT 110.500 152.755 110.640 152.910 ;
        RECT 111.420 152.910 115.790 153.050 ;
        RECT 111.420 152.755 111.560 152.910 ;
        RECT 115.470 152.850 115.790 152.910 ;
        RECT 110.425 152.525 110.715 152.755 ;
        RECT 110.885 152.525 111.175 152.755 ;
        RECT 111.345 152.525 111.635 152.755 ;
        RECT 103.970 152.370 104.290 152.430 ;
        RECT 70.390 152.230 73.380 152.370 ;
        RECT 74.620 152.230 104.290 152.370 ;
        RECT 107.280 152.370 107.420 152.510 ;
        RECT 110.960 152.370 111.100 152.525 ;
        RECT 112.250 152.510 112.570 152.770 ;
        RECT 119.700 152.755 119.840 153.590 ;
        RECT 120.530 153.530 120.850 153.590 ;
        RECT 119.625 152.525 119.915 152.755 ;
        RECT 120.545 152.525 120.835 152.755 ;
        RECT 107.280 152.230 111.100 152.370 ;
        RECT 115.930 152.370 116.250 152.430 ;
        RECT 120.620 152.370 120.760 152.525 ;
        RECT 115.930 152.230 120.760 152.370 ;
        RECT 70.390 152.170 70.710 152.230 ;
        RECT 33.605 151.845 33.895 152.075 ;
        RECT 34.970 152.030 35.290 152.090 ;
        RECT 37.745 152.030 38.035 152.075 ;
        RECT 34.970 151.890 38.035 152.030 ;
        RECT 34.970 151.830 35.290 151.890 ;
        RECT 37.745 151.845 38.035 151.890 ;
        RECT 58.675 152.030 58.965 152.075 ;
        RECT 59.810 152.030 60.130 152.090 ;
        RECT 58.675 151.890 60.130 152.030 ;
        RECT 58.675 151.845 58.965 151.890 ;
        RECT 59.810 151.830 60.130 151.890 ;
        RECT 68.090 152.030 68.410 152.090 ;
        RECT 72.245 152.030 72.535 152.075 ;
        RECT 74.620 152.030 74.760 152.230 ;
        RECT 103.970 152.170 104.290 152.230 ;
        RECT 115.930 152.170 116.250 152.230 ;
        RECT 68.090 151.890 74.760 152.030 ;
        RECT 68.090 151.830 68.410 151.890 ;
        RECT 72.245 151.845 72.535 151.890 ;
        RECT 74.990 151.830 75.310 152.090 ;
        RECT 91.105 152.030 91.395 152.075 ;
        RECT 92.930 152.030 93.250 152.090 ;
        RECT 91.105 151.890 93.250 152.030 ;
        RECT 91.105 151.845 91.395 151.890 ;
        RECT 92.930 151.830 93.250 151.890 ;
        RECT 105.350 151.830 105.670 152.090 ;
        RECT 108.110 152.030 108.430 152.090 ;
        RECT 109.045 152.030 109.335 152.075 ;
        RECT 108.110 151.890 109.335 152.030 ;
        RECT 108.110 151.830 108.430 151.890 ;
        RECT 109.045 151.845 109.335 151.890 ;
        RECT 117.770 152.030 118.090 152.090 ;
        RECT 119.165 152.030 119.455 152.075 ;
        RECT 117.770 151.890 119.455 152.030 ;
        RECT 117.770 151.830 118.090 151.890 ;
        RECT 119.165 151.845 119.455 151.890 ;
        RECT 121.465 152.030 121.755 152.075 ;
        RECT 123.290 152.030 123.610 152.090 ;
        RECT 121.465 151.890 123.610 152.030 ;
        RECT 121.465 151.845 121.755 151.890 ;
        RECT 123.290 151.830 123.610 151.890 ;
        RECT 27.855 151.010 28.145 151.055 ;
        RECT 48.325 151.010 48.615 151.055 ;
        RECT 53.370 151.010 53.690 151.070 ;
        RECT 27.855 150.870 37.500 151.010 ;
        RECT 27.855 150.825 28.145 150.870 ;
        RECT 37.360 150.730 37.500 150.870 ;
        RECT 48.325 150.870 53.690 151.010 ;
        RECT 48.325 150.825 48.615 150.870 ;
        RECT 53.370 150.810 53.690 150.870 ;
        RECT 60.730 151.010 61.050 151.070 ;
        RECT 61.665 151.010 61.955 151.055 ;
        RECT 60.730 150.870 61.955 151.010 ;
        RECT 60.730 150.810 61.050 150.870 ;
        RECT 61.665 150.825 61.955 150.870 ;
        RECT 64.885 151.010 65.175 151.055 ;
        RECT 65.790 151.010 66.110 151.070 ;
        RECT 64.885 150.870 66.110 151.010 ;
        RECT 64.885 150.825 65.175 150.870 ;
        RECT 65.790 150.810 66.110 150.870 ;
        RECT 85.570 151.010 85.890 151.070 ;
        RECT 86.045 151.010 86.335 151.055 ;
        RECT 98.235 151.010 98.525 151.055 ;
        RECT 98.910 151.010 99.230 151.070 ;
        RECT 85.570 150.870 99.230 151.010 ;
        RECT 85.570 150.810 85.890 150.870 ;
        RECT 86.045 150.825 86.335 150.870 ;
        RECT 98.235 150.825 98.525 150.870 ;
        RECT 98.910 150.810 99.230 150.870 ;
        RECT 103.970 151.010 104.290 151.070 ;
        RECT 108.570 151.010 108.890 151.070 ;
        RECT 103.970 150.870 108.890 151.010 ;
        RECT 103.970 150.810 104.290 150.870 ;
        RECT 108.570 150.810 108.890 150.870 ;
        RECT 18.360 150.670 18.650 150.715 ;
        RECT 20.710 150.670 21.030 150.730 ;
        RECT 21.620 150.670 21.910 150.715 ;
        RECT 18.360 150.530 21.910 150.670 ;
        RECT 18.360 150.485 18.650 150.530 ;
        RECT 20.710 150.470 21.030 150.530 ;
        RECT 21.620 150.485 21.910 150.530 ;
        RECT 22.540 150.670 22.830 150.715 ;
        RECT 24.400 150.670 24.690 150.715 ;
        RECT 22.540 150.530 24.690 150.670 ;
        RECT 22.540 150.485 22.830 150.530 ;
        RECT 24.400 150.485 24.690 150.530 ;
        RECT 29.860 150.670 30.150 150.715 ;
        RECT 31.290 150.670 31.610 150.730 ;
        RECT 33.120 150.670 33.410 150.715 ;
        RECT 29.860 150.530 33.410 150.670 ;
        RECT 29.860 150.485 30.150 150.530 ;
        RECT 20.220 150.330 20.510 150.375 ;
        RECT 22.540 150.330 22.755 150.485 ;
        RECT 31.290 150.470 31.610 150.530 ;
        RECT 33.120 150.485 33.410 150.530 ;
        RECT 34.040 150.670 34.330 150.715 ;
        RECT 35.900 150.670 36.190 150.715 ;
        RECT 34.040 150.530 36.190 150.670 ;
        RECT 34.040 150.485 34.330 150.530 ;
        RECT 35.900 150.485 36.190 150.530 ;
        RECT 37.270 150.670 37.590 150.730 ;
        RECT 58.905 150.670 59.195 150.715 ;
        RECT 37.270 150.530 42.100 150.670 ;
        RECT 20.220 150.190 22.755 150.330 ;
        RECT 31.720 150.330 32.010 150.375 ;
        RECT 34.040 150.330 34.255 150.485 ;
        RECT 37.270 150.470 37.590 150.530 ;
        RECT 31.720 150.190 34.255 150.330 ;
        RECT 34.510 150.330 34.830 150.390 ;
        RECT 34.985 150.330 35.275 150.375 ;
        RECT 34.510 150.190 35.275 150.330 ;
        RECT 20.220 150.145 20.510 150.190 ;
        RECT 31.720 150.145 32.010 150.190 ;
        RECT 34.510 150.130 34.830 150.190 ;
        RECT 34.985 150.145 35.275 150.190 ;
        RECT 40.950 150.130 41.270 150.390 ;
        RECT 41.960 150.375 42.100 150.530 ;
        RECT 53.920 150.530 59.195 150.670 ;
        RECT 53.920 150.390 54.060 150.530 ;
        RECT 58.905 150.485 59.195 150.530 ;
        RECT 73.165 150.670 73.455 150.715 ;
        RECT 74.990 150.670 75.310 150.730 ;
        RECT 75.465 150.670 75.755 150.715 ;
        RECT 73.165 150.530 75.755 150.670 ;
        RECT 73.165 150.485 73.455 150.530 ;
        RECT 74.990 150.470 75.310 150.530 ;
        RECT 75.465 150.485 75.755 150.530 ;
        RECT 75.910 150.670 76.230 150.730 ;
        RECT 92.930 150.715 93.250 150.730 ;
        RECT 90.190 150.670 90.480 150.715 ;
        RECT 92.050 150.670 92.340 150.715 ;
        RECT 75.910 150.530 79.360 150.670 ;
        RECT 75.910 150.470 76.230 150.530 ;
        RECT 41.885 150.145 42.175 150.375 ;
        RECT 42.330 150.130 42.650 150.390 ;
        RECT 42.790 150.130 43.110 150.390 ;
        RECT 46.025 150.145 46.315 150.375 ;
        RECT 46.470 150.330 46.790 150.390 ;
        RECT 46.945 150.330 47.235 150.375 ;
        RECT 46.470 150.190 47.235 150.330 ;
        RECT 23.470 149.790 23.790 150.050 ;
        RECT 25.325 149.990 25.615 150.035 ;
        RECT 25.770 149.990 26.090 150.050 ;
        RECT 36.825 149.990 37.115 150.035 ;
        RECT 25.325 149.850 37.115 149.990 ;
        RECT 25.325 149.805 25.615 149.850 ;
        RECT 25.770 149.790 26.090 149.850 ;
        RECT 36.825 149.805 37.115 149.850 ;
        RECT 20.220 149.650 20.510 149.695 ;
        RECT 23.000 149.650 23.290 149.695 ;
        RECT 24.860 149.650 25.150 149.695 ;
        RECT 20.220 149.510 25.150 149.650 ;
        RECT 20.220 149.465 20.510 149.510 ;
        RECT 23.000 149.465 23.290 149.510 ;
        RECT 24.860 149.465 25.150 149.510 ;
        RECT 31.720 149.650 32.010 149.695 ;
        RECT 34.500 149.650 34.790 149.695 ;
        RECT 36.360 149.650 36.650 149.695 ;
        RECT 31.720 149.510 36.650 149.650 ;
        RECT 31.720 149.465 32.010 149.510 ;
        RECT 34.500 149.465 34.790 149.510 ;
        RECT 36.360 149.465 36.650 149.510 ;
        RECT 40.950 149.650 41.270 149.710 ;
        RECT 42.880 149.650 43.020 150.130 ;
        RECT 46.100 149.990 46.240 150.145 ;
        RECT 46.470 150.130 46.790 150.190 ;
        RECT 46.945 150.145 47.235 150.190 ;
        RECT 47.390 150.130 47.710 150.390 ;
        RECT 48.770 150.130 49.090 150.390 ;
        RECT 49.690 150.130 50.010 150.390 ;
        RECT 50.150 150.130 50.470 150.390 ;
        RECT 51.070 150.330 51.390 150.390 ;
        RECT 52.925 150.330 53.215 150.375 ;
        RECT 51.070 150.190 53.215 150.330 ;
        RECT 51.070 150.130 51.390 150.190 ;
        RECT 52.925 150.145 53.215 150.190 ;
        RECT 53.385 150.145 53.675 150.375 ;
        RECT 51.545 149.990 51.835 150.035 ;
        RECT 46.100 149.850 51.835 149.990 ;
        RECT 51.545 149.805 51.835 149.850 ;
        RECT 40.950 149.510 43.020 149.650 ;
        RECT 53.000 149.650 53.140 150.145 ;
        RECT 53.460 149.990 53.600 150.145 ;
        RECT 53.830 150.130 54.150 150.390 ;
        RECT 54.750 150.130 55.070 150.390 ;
        RECT 59.350 150.130 59.670 150.390 ;
        RECT 62.585 150.330 62.875 150.375 ;
        RECT 61.280 150.190 62.875 150.330 ;
        RECT 57.050 149.990 57.370 150.050 ;
        RECT 53.460 149.850 57.370 149.990 ;
        RECT 57.050 149.790 57.370 149.850 ;
        RECT 58.445 149.990 58.735 150.035 ;
        RECT 58.445 149.850 60.960 149.990 ;
        RECT 58.445 149.805 58.735 149.850 ;
        RECT 56.590 149.650 56.910 149.710 ;
        RECT 53.000 149.510 56.910 149.650 ;
        RECT 40.950 149.450 41.270 149.510 ;
        RECT 56.590 149.450 56.910 149.510 ;
        RECT 16.355 149.310 16.645 149.355 ;
        RECT 22.550 149.310 22.870 149.370 ;
        RECT 16.355 149.170 22.870 149.310 ;
        RECT 16.355 149.125 16.645 149.170 ;
        RECT 22.550 149.110 22.870 149.170 ;
        RECT 44.185 149.310 44.475 149.355 ;
        RECT 44.630 149.310 44.950 149.370 ;
        RECT 44.185 149.170 44.950 149.310 ;
        RECT 44.185 149.125 44.475 149.170 ;
        RECT 44.630 149.110 44.950 149.170 ;
        RECT 47.390 149.110 47.710 149.370 ;
        RECT 48.310 149.310 48.630 149.370 ;
        RECT 48.785 149.310 49.075 149.355 ;
        RECT 48.310 149.170 49.075 149.310 ;
        RECT 48.310 149.110 48.630 149.170 ;
        RECT 48.785 149.125 49.075 149.170 ;
        RECT 51.085 149.310 51.375 149.355 ;
        RECT 51.990 149.310 52.310 149.370 ;
        RECT 51.085 149.170 52.310 149.310 ;
        RECT 60.820 149.310 60.960 149.850 ;
        RECT 61.280 149.695 61.420 150.190 ;
        RECT 62.585 150.145 62.875 150.190 ;
        RECT 63.950 150.130 64.270 150.390 ;
        RECT 67.630 150.130 67.950 150.390 ;
        RECT 70.390 150.330 70.710 150.390 ;
        RECT 70.865 150.330 71.155 150.375 ;
        RECT 70.390 150.190 71.155 150.330 ;
        RECT 70.390 150.130 70.710 150.190 ;
        RECT 70.865 150.145 71.155 150.190 ;
        RECT 77.750 150.130 78.070 150.390 ;
        RECT 79.220 150.375 79.360 150.530 ;
        RECT 90.190 150.530 92.340 150.670 ;
        RECT 90.190 150.485 90.480 150.530 ;
        RECT 92.050 150.485 92.340 150.530 ;
        RECT 79.145 150.145 79.435 150.375 ;
        RECT 86.030 150.330 86.350 150.390 ;
        RECT 86.505 150.330 86.795 150.375 ;
        RECT 86.030 150.190 86.795 150.330 ;
        RECT 92.125 150.330 92.340 150.485 ;
        RECT 92.930 150.670 93.260 150.715 ;
        RECT 96.230 150.670 96.520 150.715 ;
        RECT 92.930 150.530 96.520 150.670 ;
        RECT 92.930 150.485 93.260 150.530 ;
        RECT 96.230 150.485 96.520 150.530 ;
        RECT 106.745 150.670 107.035 150.715 ;
        RECT 107.205 150.670 107.495 150.715 ;
        RECT 106.745 150.530 107.495 150.670 ;
        RECT 108.660 150.670 108.800 150.810 ;
        RECT 117.425 150.670 117.715 150.715 ;
        RECT 120.665 150.670 121.315 150.715 ;
        RECT 108.660 150.530 109.260 150.670 ;
        RECT 106.745 150.485 107.035 150.530 ;
        RECT 107.205 150.485 107.495 150.530 ;
        RECT 92.930 150.470 93.250 150.485 ;
        RECT 94.370 150.330 94.660 150.375 ;
        RECT 92.125 150.190 94.660 150.330 ;
        RECT 86.030 150.130 86.350 150.190 ;
        RECT 86.505 150.145 86.795 150.190 ;
        RECT 94.370 150.145 94.660 150.190 ;
        RECT 105.365 150.330 105.655 150.375 ;
        RECT 108.110 150.330 108.430 150.390 ;
        RECT 109.120 150.375 109.260 150.530 ;
        RECT 117.425 150.530 121.315 150.670 ;
        RECT 117.425 150.485 118.015 150.530 ;
        RECT 120.665 150.485 121.315 150.530 ;
        RECT 117.725 150.390 118.015 150.485 ;
        RECT 123.290 150.470 123.610 150.730 ;
        RECT 105.365 150.190 108.430 150.330 ;
        RECT 105.365 150.145 105.655 150.190 ;
        RECT 108.110 150.130 108.430 150.190 ;
        RECT 108.585 150.145 108.875 150.375 ;
        RECT 109.045 150.145 109.335 150.375 ;
        RECT 109.505 150.145 109.795 150.375 ;
        RECT 109.950 150.330 110.270 150.390 ;
        RECT 110.425 150.330 110.715 150.375 ;
        RECT 109.950 150.190 110.715 150.330 ;
        RECT 77.290 149.990 77.610 150.050 ;
        RECT 78.225 149.990 78.515 150.035 ;
        RECT 85.110 149.990 85.430 150.050 ;
        RECT 77.290 149.850 78.515 149.990 ;
        RECT 77.290 149.790 77.610 149.850 ;
        RECT 78.225 149.805 78.515 149.850 ;
        RECT 84.740 149.850 85.430 149.990 ;
        RECT 61.205 149.465 61.495 149.695 ;
        RECT 65.330 149.650 65.650 149.710 ;
        RECT 71.785 149.650 72.075 149.695 ;
        RECT 65.330 149.510 72.075 149.650 ;
        RECT 65.330 149.450 65.650 149.510 ;
        RECT 71.785 149.465 72.075 149.510 ;
        RECT 76.845 149.650 77.135 149.695 ;
        RECT 84.740 149.650 84.880 149.850 ;
        RECT 85.110 149.790 85.430 149.850 ;
        RECT 89.265 149.990 89.555 150.035 ;
        RECT 90.170 149.990 90.490 150.050 ;
        RECT 89.265 149.850 90.490 149.990 ;
        RECT 89.265 149.805 89.555 149.850 ;
        RECT 90.170 149.790 90.490 149.850 ;
        RECT 91.090 149.790 91.410 150.050 ;
        RECT 106.270 149.790 106.590 150.050 ;
        RECT 107.650 149.990 107.970 150.050 ;
        RECT 108.660 149.990 108.800 150.145 ;
        RECT 107.650 149.850 108.800 149.990 ;
        RECT 109.580 149.990 109.720 150.145 ;
        RECT 109.950 150.130 110.270 150.190 ;
        RECT 110.425 150.145 110.715 150.190 ;
        RECT 117.725 150.170 118.090 150.390 ;
        RECT 117.770 150.130 118.090 150.170 ;
        RECT 118.805 150.330 119.095 150.375 ;
        RECT 122.385 150.330 122.675 150.375 ;
        RECT 124.220 150.330 124.510 150.375 ;
        RECT 118.805 150.190 124.510 150.330 ;
        RECT 118.805 150.145 119.095 150.190 ;
        RECT 122.385 150.145 122.675 150.190 ;
        RECT 124.220 150.145 124.510 150.190 ;
        RECT 111.345 149.990 111.635 150.035 ;
        RECT 115.945 149.990 116.235 150.035 ;
        RECT 109.580 149.850 116.235 149.990 ;
        RECT 107.650 149.790 107.970 149.850 ;
        RECT 111.345 149.805 111.635 149.850 ;
        RECT 115.945 149.805 116.235 149.850 ;
        RECT 124.685 149.990 124.975 150.035 ;
        RECT 126.050 149.990 126.370 150.050 ;
        RECT 124.685 149.850 126.370 149.990 ;
        RECT 124.685 149.805 124.975 149.850 ;
        RECT 126.050 149.790 126.370 149.850 ;
        RECT 76.845 149.510 84.880 149.650 ;
        RECT 89.730 149.650 90.020 149.695 ;
        RECT 91.590 149.650 91.880 149.695 ;
        RECT 94.370 149.650 94.660 149.695 ;
        RECT 89.730 149.510 94.660 149.650 ;
        RECT 76.845 149.465 77.135 149.510 ;
        RECT 89.730 149.465 90.020 149.510 ;
        RECT 91.590 149.465 91.880 149.510 ;
        RECT 94.370 149.465 94.660 149.510 ;
        RECT 104.445 149.650 104.735 149.695 ;
        RECT 114.550 149.650 114.870 149.710 ;
        RECT 104.445 149.510 114.870 149.650 ;
        RECT 104.445 149.465 104.735 149.510 ;
        RECT 114.550 149.450 114.870 149.510 ;
        RECT 118.805 149.650 119.095 149.695 ;
        RECT 121.925 149.650 122.215 149.695 ;
        RECT 123.815 149.650 124.105 149.695 ;
        RECT 118.805 149.510 124.105 149.650 ;
        RECT 118.805 149.465 119.095 149.510 ;
        RECT 121.925 149.465 122.215 149.510 ;
        RECT 123.815 149.465 124.105 149.510 ;
        RECT 65.420 149.310 65.560 149.450 ;
        RECT 60.820 149.170 65.560 149.310 ;
        RECT 51.085 149.125 51.375 149.170 ;
        RECT 51.990 149.110 52.310 149.170 ;
        RECT 68.550 149.110 68.870 149.370 ;
        RECT 69.945 149.310 70.235 149.355 ;
        RECT 70.850 149.310 71.170 149.370 ;
        RECT 69.945 149.170 71.170 149.310 ;
        RECT 69.945 149.125 70.235 149.170 ;
        RECT 70.850 149.110 71.170 149.170 ;
        RECT 76.370 149.310 76.690 149.370 ;
        RECT 78.225 149.310 78.515 149.355 ;
        RECT 76.370 149.170 78.515 149.310 ;
        RECT 76.370 149.110 76.690 149.170 ;
        RECT 78.225 149.125 78.515 149.170 ;
        RECT 80.065 149.310 80.355 149.355 ;
        RECT 86.950 149.310 87.270 149.370 ;
        RECT 80.065 149.170 87.270 149.310 ;
        RECT 80.065 149.125 80.355 149.170 ;
        RECT 86.950 149.110 87.270 149.170 ;
        RECT 88.345 149.310 88.635 149.355 ;
        RECT 90.630 149.310 90.950 149.370 ;
        RECT 88.345 149.170 90.950 149.310 ;
        RECT 88.345 149.125 88.635 149.170 ;
        RECT 90.630 149.110 90.950 149.170 ;
        RECT 106.745 149.310 107.035 149.355 ;
        RECT 113.630 149.310 113.950 149.370 ;
        RECT 106.745 149.170 113.950 149.310 ;
        RECT 106.745 149.125 107.035 149.170 ;
        RECT 113.630 149.110 113.950 149.170 ;
        RECT 114.090 149.110 114.410 149.370 ;
        RECT 23.470 148.290 23.790 148.350 ;
        RECT 26.705 148.290 26.995 148.335 ;
        RECT 23.470 148.150 26.995 148.290 ;
        RECT 23.470 148.090 23.790 148.150 ;
        RECT 26.705 148.105 26.995 148.150 ;
        RECT 35.890 148.290 36.210 148.350 ;
        RECT 41.870 148.290 42.190 148.350 ;
        RECT 48.770 148.290 49.090 148.350 ;
        RECT 55.685 148.290 55.975 148.335 ;
        RECT 67.170 148.290 67.490 148.350 ;
        RECT 35.890 148.150 43.020 148.290 ;
        RECT 35.890 148.090 36.210 148.150 ;
        RECT 41.870 148.090 42.190 148.150 ;
        RECT 22.090 147.950 22.410 148.010 ;
        RECT 42.330 147.950 42.650 148.010 ;
        RECT 22.090 147.810 36.120 147.950 ;
        RECT 22.090 147.750 22.410 147.810 ;
        RECT 21.170 147.410 21.490 147.670 ;
        RECT 23.930 147.610 24.250 147.670 ;
        RECT 31.840 147.655 31.980 147.810 ;
        RECT 23.930 147.470 27.840 147.610 ;
        RECT 23.930 147.410 24.250 147.470 ;
        RECT 21.645 147.270 21.935 147.315 ;
        RECT 22.550 147.270 22.870 147.330 ;
        RECT 21.645 147.130 24.160 147.270 ;
        RECT 21.645 147.085 21.935 147.130 ;
        RECT 22.550 147.070 22.870 147.130 ;
        RECT 24.020 146.930 24.160 147.130 ;
        RECT 25.310 147.070 25.630 147.330 ;
        RECT 27.700 147.315 27.840 147.470 ;
        RECT 31.765 147.425 32.055 147.655 ;
        RECT 32.225 147.425 32.515 147.655 ;
        RECT 35.980 147.610 36.120 147.810 ;
        RECT 37.360 147.810 42.650 147.950 ;
        RECT 35.980 147.470 37.040 147.610 ;
        RECT 27.625 147.085 27.915 147.315 ;
        RECT 28.085 147.270 28.375 147.315 ;
        RECT 29.450 147.270 29.770 147.330 ;
        RECT 28.085 147.130 29.770 147.270 ;
        RECT 28.085 147.085 28.375 147.130 ;
        RECT 29.450 147.070 29.770 147.130 ;
        RECT 30.830 147.270 31.150 147.330 ;
        RECT 32.300 147.270 32.440 147.425 ;
        RECT 30.830 147.130 32.440 147.270 ;
        RECT 30.830 147.070 31.150 147.130 ;
        RECT 35.890 147.070 36.210 147.330 ;
        RECT 36.900 147.315 37.040 147.470 ;
        RECT 37.360 147.315 37.500 147.810 ;
        RECT 36.825 147.085 37.115 147.315 ;
        RECT 37.285 147.085 37.575 147.315 ;
        RECT 37.745 147.270 38.035 147.315 ;
        RECT 40.950 147.270 41.270 147.330 ;
        RECT 41.500 147.315 41.640 147.810 ;
        RECT 42.330 147.750 42.650 147.810 ;
        RECT 42.880 147.950 43.020 148.150 ;
        RECT 48.770 148.150 55.975 148.290 ;
        RECT 48.770 148.090 49.090 148.150 ;
        RECT 55.685 148.105 55.975 148.150 ;
        RECT 56.220 148.150 67.490 148.290 ;
        RECT 56.220 147.950 56.360 148.150 ;
        RECT 67.170 148.090 67.490 148.150 ;
        RECT 68.550 148.290 68.870 148.350 ;
        RECT 77.750 148.290 78.070 148.350 ;
        RECT 80.065 148.290 80.355 148.335 ;
        RECT 68.550 148.150 76.600 148.290 ;
        RECT 68.550 148.090 68.870 148.150 ;
        RECT 42.880 147.810 56.360 147.950 ;
        RECT 57.050 147.950 57.370 148.010 ;
        RECT 71.325 147.950 71.615 147.995 ;
        RECT 76.460 147.950 76.600 148.150 ;
        RECT 77.750 148.150 80.355 148.290 ;
        RECT 77.750 148.090 78.070 148.150 ;
        RECT 80.065 148.105 80.355 148.150 ;
        RECT 85.110 148.290 85.430 148.350 ;
        RECT 103.985 148.290 104.275 148.335 ;
        RECT 106.285 148.290 106.575 148.335 ;
        RECT 106.730 148.290 107.050 148.350 ;
        RECT 85.110 148.150 97.760 148.290 ;
        RECT 85.110 148.090 85.430 148.150 ;
        RECT 83.270 147.950 83.590 148.010 ;
        RECT 57.050 147.810 76.140 147.950 ;
        RECT 42.880 147.315 43.020 147.810 ;
        RECT 57.050 147.750 57.370 147.810 ;
        RECT 71.325 147.765 71.615 147.810 ;
        RECT 53.830 147.610 54.150 147.670 ;
        RECT 53.460 147.470 54.150 147.610 ;
        RECT 53.460 147.315 53.600 147.470 ;
        RECT 53.830 147.410 54.150 147.470 ;
        RECT 54.290 147.610 54.610 147.670 ;
        RECT 54.765 147.610 55.055 147.655 ;
        RECT 60.745 147.610 61.035 147.655 ;
        RECT 65.330 147.610 65.650 147.670 ;
        RECT 54.290 147.470 65.650 147.610 ;
        RECT 54.290 147.410 54.610 147.470 ;
        RECT 54.765 147.425 55.055 147.470 ;
        RECT 60.745 147.425 61.035 147.470 ;
        RECT 65.330 147.410 65.650 147.470 ;
        RECT 70.390 147.610 70.710 147.670 ;
        RECT 70.390 147.470 72.920 147.610 ;
        RECT 70.390 147.410 70.710 147.470 ;
        RECT 37.745 147.130 41.270 147.270 ;
        RECT 37.745 147.085 38.035 147.130 ;
        RECT 40.950 147.070 41.270 147.130 ;
        RECT 41.425 147.085 41.715 147.315 ;
        RECT 41.885 147.250 42.175 147.315 ;
        RECT 41.885 147.110 42.560 147.250 ;
        RECT 41.885 147.085 42.175 147.110 ;
        RECT 42.420 146.930 42.560 147.110 ;
        RECT 42.805 147.085 43.095 147.315 ;
        RECT 53.385 147.085 53.675 147.315 ;
        RECT 56.590 147.270 56.910 147.330 ;
        RECT 57.065 147.270 57.355 147.315 ;
        RECT 56.590 147.130 57.355 147.270 ;
        RECT 56.590 147.070 56.910 147.130 ;
        RECT 57.065 147.085 57.355 147.130 ;
        RECT 57.510 147.070 57.830 147.330 ;
        RECT 57.985 147.085 58.275 147.315 ;
        RECT 58.890 147.270 59.210 147.330 ;
        RECT 68.550 147.270 68.870 147.330 ;
        RECT 58.890 147.130 68.870 147.270 ;
        RECT 24.020 146.790 42.560 146.930 ;
        RECT 52.450 146.930 52.770 146.990 ;
        RECT 53.845 146.930 54.135 146.975 ;
        RECT 52.450 146.790 54.135 146.930 ;
        RECT 58.060 146.930 58.200 147.085 ;
        RECT 58.890 147.070 59.210 147.130 ;
        RECT 68.550 147.070 68.870 147.130 ;
        RECT 71.770 147.270 72.090 147.330 ;
        RECT 72.780 147.315 72.920 147.470 ;
        RECT 72.245 147.270 72.535 147.315 ;
        RECT 71.770 147.130 72.535 147.270 ;
        RECT 71.770 147.070 72.090 147.130 ;
        RECT 72.245 147.085 72.535 147.130 ;
        RECT 72.705 147.085 72.995 147.315 ;
        RECT 59.350 146.930 59.670 146.990 ;
        RECT 61.205 146.930 61.495 146.975 ;
        RECT 58.060 146.790 61.495 146.930 ;
        RECT 52.450 146.730 52.770 146.790 ;
        RECT 53.845 146.745 54.135 146.790 ;
        RECT 59.350 146.730 59.670 146.790 ;
        RECT 61.205 146.745 61.495 146.790 ;
        RECT 61.650 146.730 61.970 146.990 ;
        RECT 76.000 146.930 76.140 147.810 ;
        RECT 76.460 147.810 83.590 147.950 ;
        RECT 76.460 147.315 76.600 147.810 ;
        RECT 83.270 147.750 83.590 147.810 ;
        RECT 89.220 147.950 89.510 147.995 ;
        RECT 92.000 147.950 92.290 147.995 ;
        RECT 93.860 147.950 94.150 147.995 ;
        RECT 89.220 147.810 94.150 147.950 ;
        RECT 89.220 147.765 89.510 147.810 ;
        RECT 92.000 147.765 92.290 147.810 ;
        RECT 93.860 147.765 94.150 147.810 ;
        RECT 85.570 147.610 85.890 147.670 ;
        RECT 77.380 147.470 85.890 147.610 ;
        RECT 77.380 147.315 77.520 147.470 ;
        RECT 85.570 147.410 85.890 147.470 ;
        RECT 90.170 147.610 90.490 147.670 ;
        RECT 97.620 147.655 97.760 148.150 ;
        RECT 103.985 148.150 106.040 148.290 ;
        RECT 103.985 148.105 104.275 148.150 ;
        RECT 104.890 147.750 105.210 148.010 ;
        RECT 105.900 147.950 106.040 148.150 ;
        RECT 106.285 148.150 107.050 148.290 ;
        RECT 106.285 148.105 106.575 148.150 ;
        RECT 106.730 148.090 107.050 148.150 ;
        RECT 115.930 148.090 116.250 148.350 ;
        RECT 120.500 147.950 120.790 147.995 ;
        RECT 123.280 147.950 123.570 147.995 ;
        RECT 125.140 147.950 125.430 147.995 ;
        RECT 105.900 147.810 119.610 147.950 ;
        RECT 92.485 147.610 92.775 147.655 ;
        RECT 90.170 147.470 92.775 147.610 ;
        RECT 90.170 147.410 90.490 147.470 ;
        RECT 92.485 147.425 92.775 147.470 ;
        RECT 97.545 147.425 97.835 147.655 ;
        RECT 98.465 147.610 98.755 147.655 ;
        RECT 104.980 147.610 105.120 147.750 ;
        RECT 105.825 147.610 106.115 147.655 ;
        RECT 98.465 147.470 103.280 147.610 ;
        RECT 104.980 147.470 106.115 147.610 ;
        RECT 98.465 147.425 98.755 147.470 ;
        RECT 76.385 147.085 76.675 147.315 ;
        RECT 77.305 147.085 77.595 147.315 ;
        RECT 77.765 147.085 78.055 147.315 ;
        RECT 78.210 147.270 78.530 147.330 ;
        RECT 81.430 147.270 81.750 147.330 ;
        RECT 78.210 147.130 81.750 147.270 ;
        RECT 77.840 146.930 77.980 147.085 ;
        RECT 78.210 147.070 78.530 147.130 ;
        RECT 81.430 147.070 81.750 147.130 ;
        RECT 81.890 147.070 82.210 147.330 ;
        RECT 82.365 147.085 82.655 147.315 ;
        RECT 81.980 146.930 82.120 147.070 ;
        RECT 76.000 146.790 82.120 146.930 ;
        RECT 22.090 146.390 22.410 146.650 ;
        RECT 23.930 146.390 24.250 146.650 ;
        RECT 25.770 146.390 26.090 146.650 ;
        RECT 27.150 146.590 27.470 146.650 ;
        RECT 29.005 146.590 29.295 146.635 ;
        RECT 27.150 146.450 29.295 146.590 ;
        RECT 27.150 146.390 27.470 146.450 ;
        RECT 29.005 146.405 29.295 146.450 ;
        RECT 29.450 146.390 29.770 146.650 ;
        RECT 31.305 146.590 31.595 146.635 ;
        RECT 37.270 146.590 37.590 146.650 ;
        RECT 31.305 146.450 37.590 146.590 ;
        RECT 31.305 146.405 31.595 146.450 ;
        RECT 37.270 146.390 37.590 146.450 ;
        RECT 38.650 146.590 38.970 146.650 ;
        RECT 39.125 146.590 39.415 146.635 ;
        RECT 38.650 146.450 39.415 146.590 ;
        RECT 38.650 146.390 38.970 146.450 ;
        RECT 39.125 146.405 39.415 146.450 ;
        RECT 39.570 146.390 39.890 146.650 ;
        RECT 51.545 146.590 51.835 146.635 ;
        RECT 52.910 146.590 53.230 146.650 ;
        RECT 51.545 146.450 53.230 146.590 ;
        RECT 51.545 146.405 51.835 146.450 ;
        RECT 52.910 146.390 53.230 146.450 ;
        RECT 63.505 146.590 63.795 146.635 ;
        RECT 63.950 146.590 64.270 146.650 ;
        RECT 63.505 146.450 64.270 146.590 ;
        RECT 63.505 146.405 63.795 146.450 ;
        RECT 63.950 146.390 64.270 146.450 ;
        RECT 73.150 146.590 73.470 146.650 ;
        RECT 73.625 146.590 73.915 146.635 ;
        RECT 78.210 146.590 78.530 146.650 ;
        RECT 73.150 146.450 78.530 146.590 ;
        RECT 73.150 146.390 73.470 146.450 ;
        RECT 73.625 146.405 73.915 146.450 ;
        RECT 78.210 146.390 78.530 146.450 ;
        RECT 79.590 146.390 79.910 146.650 ;
        RECT 82.440 146.590 82.580 147.085 ;
        RECT 83.270 147.070 83.590 147.330 ;
        RECT 84.665 147.270 84.955 147.315 ;
        RECT 86.490 147.270 86.810 147.330 ;
        RECT 84.665 147.130 86.810 147.270 ;
        RECT 84.665 147.085 84.955 147.130 ;
        RECT 86.490 147.070 86.810 147.130 ;
        RECT 89.220 147.270 89.510 147.315 ;
        RECT 93.850 147.270 94.170 147.330 ;
        RECT 94.325 147.270 94.615 147.315 ;
        RECT 89.220 147.130 91.755 147.270 ;
        RECT 89.220 147.085 89.510 147.130 ;
        RECT 91.540 146.975 91.755 147.130 ;
        RECT 93.850 147.130 94.615 147.270 ;
        RECT 93.850 147.070 94.170 147.130 ;
        RECT 94.325 147.085 94.615 147.130 ;
        RECT 95.690 147.070 96.010 147.330 ;
        RECT 96.150 147.270 96.470 147.330 ;
        RECT 98.540 147.270 98.680 147.425 ;
        RECT 96.150 147.130 98.680 147.270 ;
        RECT 96.150 147.070 96.470 147.130 ;
        RECT 98.910 147.070 99.230 147.330 ;
        RECT 102.145 147.270 102.435 147.315 ;
        RECT 100.840 147.130 102.435 147.270 ;
        RECT 84.205 146.930 84.495 146.975 ;
        RECT 87.360 146.930 87.650 146.975 ;
        RECT 90.620 146.930 90.910 146.975 ;
        RECT 84.205 146.790 90.910 146.930 ;
        RECT 84.205 146.745 84.495 146.790 ;
        RECT 87.360 146.745 87.650 146.790 ;
        RECT 90.620 146.745 90.910 146.790 ;
        RECT 91.540 146.930 91.830 146.975 ;
        RECT 93.400 146.930 93.690 146.975 ;
        RECT 91.540 146.790 93.690 146.930 ;
        RECT 91.540 146.745 91.830 146.790 ;
        RECT 93.400 146.745 93.690 146.790 ;
        RECT 85.355 146.590 85.645 146.635 ;
        RECT 86.030 146.590 86.350 146.650 ;
        RECT 82.440 146.450 86.350 146.590 ;
        RECT 85.355 146.405 85.645 146.450 ;
        RECT 86.030 146.390 86.350 146.450 ;
        RECT 96.165 146.590 96.455 146.635 ;
        RECT 97.070 146.590 97.390 146.650 ;
        RECT 100.840 146.635 100.980 147.130 ;
        RECT 102.145 147.085 102.435 147.130 ;
        RECT 103.140 146.930 103.280 147.470 ;
        RECT 105.825 147.425 106.115 147.470 ;
        RECT 106.360 147.470 110.640 147.610 ;
        RECT 104.905 147.270 105.195 147.315 ;
        RECT 105.350 147.270 105.670 147.330 ;
        RECT 106.360 147.270 106.500 147.470 ;
        RECT 104.905 147.130 105.670 147.270 ;
        RECT 104.905 147.085 105.195 147.130 ;
        RECT 105.350 147.070 105.670 147.130 ;
        RECT 105.900 147.130 106.500 147.270 ;
        RECT 105.900 146.930 106.040 147.130 ;
        RECT 108.110 147.070 108.430 147.330 ;
        RECT 108.570 147.070 108.890 147.330 ;
        RECT 109.045 147.085 109.335 147.315 ;
        RECT 103.140 146.790 106.040 146.930 ;
        RECT 106.285 146.930 106.575 146.975 ;
        RECT 106.745 146.930 107.035 146.975 ;
        RECT 106.285 146.790 107.035 146.930 ;
        RECT 106.285 146.745 106.575 146.790 ;
        RECT 106.745 146.745 107.035 146.790 ;
        RECT 96.165 146.450 97.390 146.590 ;
        RECT 96.165 146.405 96.455 146.450 ;
        RECT 97.070 146.390 97.390 146.450 ;
        RECT 100.765 146.405 101.055 146.635 ;
        RECT 103.065 146.590 103.355 146.635 ;
        RECT 103.970 146.590 104.290 146.650 ;
        RECT 103.065 146.450 104.290 146.590 ;
        RECT 103.065 146.405 103.355 146.450 ;
        RECT 103.970 146.390 104.290 146.450 ;
        RECT 104.430 146.590 104.750 146.650 ;
        RECT 109.120 146.590 109.260 147.085 ;
        RECT 109.950 147.070 110.270 147.330 ;
        RECT 110.500 147.270 110.640 147.470 ;
        RECT 112.710 147.410 113.030 147.670 ;
        RECT 119.470 147.610 119.610 147.810 ;
        RECT 120.500 147.810 125.430 147.950 ;
        RECT 120.500 147.765 120.790 147.810 ;
        RECT 123.280 147.765 123.570 147.810 ;
        RECT 125.140 147.765 125.430 147.810 ;
        RECT 119.470 147.470 125.360 147.610 ;
        RECT 125.220 147.330 125.360 147.470 ;
        RECT 114.105 147.270 114.395 147.315 ;
        RECT 110.500 147.130 114.395 147.270 ;
        RECT 114.105 147.085 114.395 147.130 ;
        RECT 120.500 147.270 120.790 147.315 ;
        RECT 120.500 147.130 123.035 147.270 ;
        RECT 120.500 147.085 120.790 147.130 ;
        RECT 116.635 146.930 116.925 146.975 ;
        RECT 117.770 146.930 118.090 146.990 ;
        RECT 116.635 146.790 118.090 146.930 ;
        RECT 116.635 146.745 116.925 146.790 ;
        RECT 117.770 146.730 118.090 146.790 ;
        RECT 118.640 146.930 118.930 146.975 ;
        RECT 120.990 146.930 121.310 146.990 ;
        RECT 122.820 146.975 123.035 147.130 ;
        RECT 123.750 147.070 124.070 147.330 ;
        RECT 125.130 147.070 125.450 147.330 ;
        RECT 125.605 147.270 125.895 147.315 ;
        RECT 126.050 147.270 126.370 147.330 ;
        RECT 125.605 147.130 126.370 147.270 ;
        RECT 125.605 147.085 125.895 147.130 ;
        RECT 126.050 147.070 126.370 147.130 ;
        RECT 121.900 146.930 122.190 146.975 ;
        RECT 118.640 146.790 122.190 146.930 ;
        RECT 118.640 146.745 118.930 146.790 ;
        RECT 120.990 146.730 121.310 146.790 ;
        RECT 121.900 146.745 122.190 146.790 ;
        RECT 122.820 146.930 123.110 146.975 ;
        RECT 124.680 146.930 124.970 146.975 ;
        RECT 122.820 146.790 124.970 146.930 ;
        RECT 122.820 146.745 123.110 146.790 ;
        RECT 124.680 146.745 124.970 146.790 ;
        RECT 104.430 146.450 109.260 146.590 ;
        RECT 113.645 146.590 113.935 146.635 ;
        RECT 114.090 146.590 114.410 146.650 ;
        RECT 117.310 146.590 117.630 146.650 ;
        RECT 113.645 146.450 117.630 146.590 ;
        RECT 104.430 146.390 104.750 146.450 ;
        RECT 113.645 146.405 113.935 146.450 ;
        RECT 114.090 146.390 114.410 146.450 ;
        RECT 117.310 146.390 117.630 146.450 ;
        RECT 20.710 145.370 21.030 145.630 ;
        RECT 22.090 145.615 22.410 145.630 ;
        RECT 22.090 145.385 22.625 145.615 ;
        RECT 25.310 145.570 25.630 145.630 ;
        RECT 41.425 145.570 41.715 145.615 ;
        RECT 56.590 145.570 56.910 145.630 ;
        RECT 73.150 145.570 73.470 145.630 ;
        RECT 25.310 145.430 41.180 145.570 ;
        RECT 22.090 145.370 22.410 145.385 ;
        RECT 25.310 145.370 25.630 145.430 ;
        RECT 24.340 145.230 24.630 145.275 ;
        RECT 25.770 145.230 26.090 145.290 ;
        RECT 27.600 145.230 27.890 145.275 ;
        RECT 24.340 145.090 27.890 145.230 ;
        RECT 24.340 145.045 24.630 145.090 ;
        RECT 25.770 145.030 26.090 145.090 ;
        RECT 27.600 145.045 27.890 145.090 ;
        RECT 28.520 145.230 28.810 145.275 ;
        RECT 30.380 145.230 30.670 145.275 ;
        RECT 28.520 145.090 30.670 145.230 ;
        RECT 28.520 145.045 28.810 145.090 ;
        RECT 30.380 145.045 30.670 145.090 ;
        RECT 18.870 144.890 19.190 144.950 ;
        RECT 21.185 144.890 21.475 144.935 ;
        RECT 25.310 144.890 25.630 144.950 ;
        RECT 18.870 144.750 25.630 144.890 ;
        RECT 18.870 144.690 19.190 144.750 ;
        RECT 21.185 144.705 21.475 144.750 ;
        RECT 25.310 144.690 25.630 144.750 ;
        RECT 26.200 144.890 26.490 144.935 ;
        RECT 28.520 144.890 28.735 145.045 ;
        RECT 41.040 144.950 41.180 145.430 ;
        RECT 41.425 145.430 45.780 145.570 ;
        RECT 41.425 145.385 41.715 145.430 ;
        RECT 43.270 145.230 43.560 145.275 ;
        RECT 45.130 145.230 45.420 145.275 ;
        RECT 43.270 145.090 45.420 145.230 ;
        RECT 45.640 145.230 45.780 145.430 ;
        RECT 56.590 145.430 73.470 145.570 ;
        RECT 56.590 145.370 56.910 145.430 ;
        RECT 73.150 145.370 73.470 145.430 ;
        RECT 86.030 145.370 86.350 145.630 ;
        RECT 88.345 145.385 88.635 145.615 ;
        RECT 90.170 145.570 90.490 145.630 ;
        RECT 91.105 145.570 91.395 145.615 ;
        RECT 90.170 145.430 91.395 145.570 ;
        RECT 46.050 145.230 46.340 145.275 ;
        RECT 49.310 145.230 49.600 145.275 ;
        RECT 45.640 145.090 49.600 145.230 ;
        RECT 43.270 145.045 43.560 145.090 ;
        RECT 45.130 145.045 45.420 145.090 ;
        RECT 46.050 145.045 46.340 145.090 ;
        RECT 49.310 145.045 49.600 145.090 ;
        RECT 51.530 145.230 51.850 145.290 ;
        RECT 56.130 145.230 56.450 145.290 ;
        RECT 59.350 145.230 59.670 145.290 ;
        RECT 61.650 145.230 61.970 145.290 ;
        RECT 65.345 145.230 65.635 145.275 ;
        RECT 51.530 145.090 58.660 145.230 ;
        RECT 26.200 144.750 28.735 144.890 ;
        RECT 26.200 144.705 26.490 144.750 ;
        RECT 40.950 144.690 41.270 144.950 ;
        RECT 45.205 144.890 45.420 145.045 ;
        RECT 51.530 145.030 51.850 145.090 ;
        RECT 56.130 145.030 56.450 145.090 ;
        RECT 47.450 144.890 47.740 144.935 ;
        RECT 45.205 144.750 47.740 144.890 ;
        RECT 47.450 144.705 47.740 144.750 ;
        RECT 52.910 144.690 53.230 144.950 ;
        RECT 58.520 144.935 58.660 145.090 ;
        RECT 59.350 145.090 65.635 145.230 ;
        RECT 59.350 145.030 59.670 145.090 ;
        RECT 61.650 145.030 61.970 145.090 ;
        RECT 65.345 145.045 65.635 145.090 ;
        RECT 79.590 145.030 79.910 145.290 ;
        RECT 58.445 144.705 58.735 144.935 ;
        RECT 64.410 144.890 64.730 144.950 ;
        RECT 65.805 144.890 66.095 144.935 ;
        RECT 64.410 144.750 66.095 144.890 ;
        RECT 64.410 144.690 64.730 144.750 ;
        RECT 65.805 144.705 66.095 144.750 ;
        RECT 78.670 144.890 78.990 144.950 ;
        RECT 80.985 144.890 81.275 144.935 ;
        RECT 78.670 144.750 81.275 144.890 ;
        RECT 78.670 144.690 78.990 144.750 ;
        RECT 80.985 144.705 81.275 144.750 ;
        RECT 86.030 144.890 86.350 144.950 ;
        RECT 86.505 144.890 86.795 144.935 ;
        RECT 86.030 144.750 86.795 144.890 ;
        RECT 88.420 144.890 88.560 145.385 ;
        RECT 90.170 145.370 90.490 145.430 ;
        RECT 91.105 145.385 91.395 145.430 ;
        RECT 91.550 145.370 91.870 145.630 ;
        RECT 96.150 145.370 96.470 145.630 ;
        RECT 96.625 145.570 96.915 145.615 ;
        RECT 104.430 145.570 104.750 145.630 ;
        RECT 96.625 145.430 104.750 145.570 ;
        RECT 96.625 145.385 96.915 145.430 ;
        RECT 90.185 144.890 90.475 144.935 ;
        RECT 88.420 144.750 90.475 144.890 ;
        RECT 86.030 144.690 86.350 144.750 ;
        RECT 86.505 144.705 86.795 144.750 ;
        RECT 90.185 144.705 90.475 144.750 ;
        RECT 90.630 144.890 90.950 144.950 ;
        RECT 92.485 144.890 92.775 144.935 ;
        RECT 90.630 144.750 92.775 144.890 ;
        RECT 90.630 144.690 90.950 144.750 ;
        RECT 92.485 144.705 92.775 144.750 ;
        RECT 93.405 144.890 93.695 144.935 ;
        RECT 96.700 144.890 96.840 145.385 ;
        RECT 104.430 145.370 104.750 145.430 ;
        RECT 108.110 145.570 108.430 145.630 ;
        RECT 111.330 145.570 111.650 145.630 ;
        RECT 108.110 145.430 111.650 145.570 ;
        RECT 108.110 145.370 108.430 145.430 ;
        RECT 111.330 145.370 111.650 145.430 ;
        RECT 117.310 145.370 117.630 145.630 ;
        RECT 120.085 145.570 120.375 145.615 ;
        RECT 120.990 145.570 121.310 145.630 ;
        RECT 120.085 145.430 121.310 145.570 ;
        RECT 120.085 145.385 120.375 145.430 ;
        RECT 120.990 145.370 121.310 145.430 ;
        RECT 122.385 145.570 122.675 145.615 ;
        RECT 123.750 145.570 124.070 145.630 ;
        RECT 122.385 145.430 124.070 145.570 ;
        RECT 122.385 145.385 122.675 145.430 ;
        RECT 123.750 145.370 124.070 145.430 ;
        RECT 97.070 145.230 97.390 145.290 ;
        RECT 98.105 145.230 98.395 145.275 ;
        RECT 101.345 145.230 101.995 145.275 ;
        RECT 97.070 145.090 101.995 145.230 ;
        RECT 97.070 145.030 97.390 145.090 ;
        RECT 98.105 145.045 98.695 145.090 ;
        RECT 101.345 145.045 101.995 145.090 ;
        RECT 93.405 144.750 96.840 144.890 ;
        RECT 93.405 144.705 93.695 144.750 ;
        RECT 98.405 144.730 98.695 145.045 ;
        RECT 103.970 145.030 104.290 145.290 ;
        RECT 110.960 145.090 117.080 145.230 ;
        RECT 99.485 144.890 99.775 144.935 ;
        RECT 103.065 144.890 103.355 144.935 ;
        RECT 104.900 144.890 105.190 144.935 ;
        RECT 99.485 144.750 105.190 144.890 ;
        RECT 99.485 144.705 99.775 144.750 ;
        RECT 103.065 144.705 103.355 144.750 ;
        RECT 104.900 144.705 105.190 144.750 ;
        RECT 107.650 144.890 107.970 144.950 ;
        RECT 109.950 144.890 110.270 144.950 ;
        RECT 110.960 144.935 111.100 145.090 ;
        RECT 107.650 144.750 110.270 144.890 ;
        RECT 107.650 144.690 107.970 144.750 ;
        RECT 109.950 144.690 110.270 144.750 ;
        RECT 110.885 144.705 111.175 144.935 ;
        RECT 111.345 144.705 111.635 144.935 ;
        RECT 27.150 144.550 27.470 144.610 ;
        RECT 29.465 144.550 29.755 144.595 ;
        RECT 27.150 144.410 29.755 144.550 ;
        RECT 27.150 144.350 27.470 144.410 ;
        RECT 29.465 144.365 29.755 144.410 ;
        RECT 31.305 144.550 31.595 144.595 ;
        RECT 36.810 144.550 37.130 144.610 ;
        RECT 42.345 144.550 42.635 144.595 ;
        RECT 31.305 144.410 42.635 144.550 ;
        RECT 31.305 144.365 31.595 144.410 ;
        RECT 36.810 144.350 37.130 144.410 ;
        RECT 42.345 144.365 42.635 144.410 ;
        RECT 44.185 144.550 44.475 144.595 ;
        RECT 64.885 144.550 65.175 144.595 ;
        RECT 65.330 144.550 65.650 144.610 ;
        RECT 69.010 144.550 69.330 144.610 ;
        RECT 44.185 144.410 52.220 144.550 ;
        RECT 44.185 144.365 44.475 144.410 ;
        RECT 52.080 144.255 52.220 144.410 ;
        RECT 64.885 144.410 69.330 144.550 ;
        RECT 64.885 144.365 65.175 144.410 ;
        RECT 65.330 144.350 65.650 144.410 ;
        RECT 69.010 144.350 69.330 144.410 ;
        RECT 80.050 144.350 80.370 144.610 ;
        RECT 85.110 144.350 85.430 144.610 ;
        RECT 105.350 144.350 105.670 144.610 ;
        RECT 108.570 144.550 108.890 144.610 ;
        RECT 111.420 144.550 111.560 144.705 ;
        RECT 111.790 144.690 112.110 144.950 ;
        RECT 108.570 144.410 111.560 144.550 ;
        RECT 108.570 144.350 108.890 144.410 ;
        RECT 26.200 144.210 26.490 144.255 ;
        RECT 28.980 144.210 29.270 144.255 ;
        RECT 30.840 144.210 31.130 144.255 ;
        RECT 26.200 144.070 31.130 144.210 ;
        RECT 26.200 144.025 26.490 144.070 ;
        RECT 28.980 144.025 29.270 144.070 ;
        RECT 30.840 144.025 31.130 144.070 ;
        RECT 42.810 144.210 43.100 144.255 ;
        RECT 44.670 144.210 44.960 144.255 ;
        RECT 47.450 144.210 47.740 144.255 ;
        RECT 42.810 144.070 47.740 144.210 ;
        RECT 42.810 144.025 43.100 144.070 ;
        RECT 44.670 144.025 44.960 144.070 ;
        RECT 47.450 144.025 47.740 144.070 ;
        RECT 52.005 144.025 52.295 144.255 ;
        RECT 75.910 144.210 76.230 144.270 ;
        RECT 81.905 144.210 82.195 144.255 ;
        RECT 75.910 144.070 82.195 144.210 ;
        RECT 75.910 144.010 76.230 144.070 ;
        RECT 81.905 144.025 82.195 144.070 ;
        RECT 99.485 144.210 99.775 144.255 ;
        RECT 102.605 144.210 102.895 144.255 ;
        RECT 104.495 144.210 104.785 144.255 ;
        RECT 99.485 144.070 104.785 144.210 ;
        RECT 111.420 144.210 111.560 144.410 ;
        RECT 112.710 144.550 113.030 144.610 ;
        RECT 116.940 144.595 117.080 145.090 ;
        RECT 119.625 144.890 119.915 144.935 ;
        RECT 120.530 144.890 120.850 144.950 ;
        RECT 119.625 144.750 120.850 144.890 ;
        RECT 119.625 144.705 119.915 144.750 ;
        RECT 120.530 144.690 120.850 144.750 ;
        RECT 121.465 144.705 121.755 144.935 ;
        RECT 115.945 144.550 116.235 144.595 ;
        RECT 112.710 144.410 116.235 144.550 ;
        RECT 112.710 144.350 113.030 144.410 ;
        RECT 115.945 144.365 116.235 144.410 ;
        RECT 116.865 144.550 117.155 144.595 ;
        RECT 117.770 144.550 118.090 144.610 ;
        RECT 121.540 144.550 121.680 144.705 ;
        RECT 116.865 144.410 118.090 144.550 ;
        RECT 116.865 144.365 117.155 144.410 ;
        RECT 117.770 144.350 118.090 144.410 ;
        RECT 119.240 144.410 121.680 144.550 ;
        RECT 111.790 144.210 112.110 144.270 ;
        RECT 119.240 144.255 119.380 144.410 ;
        RECT 111.420 144.070 112.110 144.210 ;
        RECT 99.485 144.025 99.775 144.070 ;
        RECT 102.605 144.025 102.895 144.070 ;
        RECT 104.495 144.025 104.785 144.070 ;
        RECT 111.790 144.010 112.110 144.070 ;
        RECT 119.165 144.025 119.455 144.255 ;
        RECT 51.315 143.870 51.605 143.915 ;
        RECT 52.450 143.870 52.770 143.930 ;
        RECT 51.315 143.730 52.770 143.870 ;
        RECT 51.315 143.685 51.605 143.730 ;
        RECT 52.450 143.670 52.770 143.730 ;
        RECT 58.890 143.670 59.210 143.930 ;
        RECT 67.645 143.870 67.935 143.915 ;
        RECT 69.930 143.870 70.250 143.930 ;
        RECT 67.645 143.730 70.250 143.870 ;
        RECT 67.645 143.685 67.935 143.730 ;
        RECT 69.930 143.670 70.250 143.730 ;
        RECT 80.050 143.670 80.370 143.930 ;
        RECT 108.570 143.870 108.890 143.930 ;
        RECT 113.185 143.870 113.475 143.915 ;
        RECT 108.570 143.730 113.475 143.870 ;
        RECT 108.570 143.670 108.890 143.730 ;
        RECT 113.185 143.685 113.475 143.730 ;
        RECT 35.890 142.650 36.210 142.910 ;
        RECT 46.930 142.850 47.250 142.910 ;
        RECT 47.405 142.850 47.695 142.895 ;
        RECT 51.530 142.850 51.850 142.910 ;
        RECT 46.930 142.710 47.695 142.850 ;
        RECT 46.930 142.650 47.250 142.710 ;
        RECT 47.405 142.665 47.695 142.710 ;
        RECT 49.320 142.710 51.850 142.850 ;
        RECT 35.430 142.510 35.750 142.570 ;
        RECT 40.950 142.510 41.270 142.570 ;
        RECT 49.320 142.510 49.460 142.710 ;
        RECT 51.530 142.650 51.850 142.710 ;
        RECT 59.350 142.650 59.670 142.910 ;
        RECT 109.950 142.650 110.270 142.910 ;
        RECT 35.430 142.370 36.120 142.510 ;
        RECT 35.430 142.310 35.750 142.370 ;
        RECT 35.980 142.215 36.120 142.370 ;
        RECT 40.950 142.370 49.460 142.510 ;
        RECT 49.705 142.510 49.995 142.555 ;
        RECT 62.685 142.510 62.975 142.555 ;
        RECT 65.805 142.510 66.095 142.555 ;
        RECT 67.695 142.510 67.985 142.555 ;
        RECT 49.705 142.370 61.420 142.510 ;
        RECT 40.950 142.310 41.270 142.370 ;
        RECT 49.705 142.325 49.995 142.370 ;
        RECT 61.280 142.230 61.420 142.370 ;
        RECT 62.685 142.370 67.985 142.510 ;
        RECT 62.685 142.325 62.975 142.370 ;
        RECT 65.805 142.325 66.095 142.370 ;
        RECT 67.695 142.325 67.985 142.370 ;
        RECT 69.025 142.325 69.315 142.555 ;
        RECT 119.625 142.510 119.915 142.555 ;
        RECT 124.670 142.510 124.990 142.570 ;
        RECT 119.625 142.370 124.990 142.510 ;
        RECT 119.625 142.325 119.915 142.370 ;
        RECT 35.905 141.985 36.195 142.215 ;
        RECT 47.850 141.970 48.170 142.230 ;
        RECT 50.150 142.170 50.470 142.230 ;
        RECT 51.070 142.170 51.390 142.230 ;
        RECT 56.605 142.170 56.895 142.215 ;
        RECT 59.825 142.170 60.115 142.215 ;
        RECT 50.150 142.030 53.830 142.170 ;
        RECT 50.150 141.970 50.470 142.030 ;
        RECT 51.070 141.970 51.390 142.030 ;
        RECT 34.970 141.830 35.290 141.890 ;
        RECT 35.445 141.830 35.735 141.875 ;
        RECT 34.970 141.690 35.735 141.830 ;
        RECT 34.970 141.630 35.290 141.690 ;
        RECT 35.445 141.645 35.735 141.690 ;
        RECT 48.785 141.830 49.075 141.875 ;
        RECT 50.610 141.830 50.930 141.890 ;
        RECT 53.690 141.875 53.830 142.030 ;
        RECT 54.840 142.030 60.115 142.170 ;
        RECT 54.840 141.875 54.980 142.030 ;
        RECT 56.605 141.985 56.895 142.030 ;
        RECT 59.825 141.985 60.115 142.030 ;
        RECT 61.190 141.970 61.510 142.230 ;
        RECT 67.185 142.170 67.475 142.215 ;
        RECT 69.100 142.170 69.240 142.325 ;
        RECT 124.670 142.310 124.990 142.370 ;
        RECT 67.185 142.030 69.240 142.170 ;
        RECT 67.185 141.985 67.475 142.030 ;
        RECT 109.030 141.970 109.350 142.230 ;
        RECT 112.710 142.170 113.030 142.230 ;
        RECT 116.405 142.170 116.695 142.215 ;
        RECT 112.710 142.030 116.695 142.170 ;
        RECT 112.710 141.970 113.030 142.030 ;
        RECT 116.405 141.985 116.695 142.030 ;
        RECT 48.785 141.690 50.930 141.830 ;
        RECT 48.785 141.645 49.075 141.690 ;
        RECT 50.610 141.630 50.930 141.690 ;
        RECT 53.615 141.645 53.905 141.875 ;
        RECT 54.305 141.645 54.595 141.875 ;
        RECT 54.765 141.645 55.055 141.875 ;
        RECT 55.210 141.830 55.530 141.890 ;
        RECT 55.685 141.830 55.975 141.875 ;
        RECT 55.210 141.690 55.975 141.830 ;
        RECT 36.825 141.305 37.115 141.535 ;
        RECT 47.405 141.490 47.695 141.535 ;
        RECT 52.465 141.490 52.755 141.535 ;
        RECT 47.405 141.350 52.755 141.490 ;
        RECT 47.405 141.305 47.695 141.350 ;
        RECT 52.465 141.305 52.755 141.350 ;
        RECT 54.380 141.490 54.520 141.645 ;
        RECT 55.210 141.630 55.530 141.690 ;
        RECT 55.685 141.645 55.975 141.690 ;
        RECT 57.050 141.490 57.370 141.550 ;
        RECT 54.380 141.350 57.370 141.490 ;
        RECT 24.850 141.150 25.170 141.210 ;
        RECT 34.525 141.150 34.815 141.195 ;
        RECT 24.850 141.010 34.815 141.150 ;
        RECT 36.900 141.150 37.040 141.305 ;
        RECT 51.070 141.150 51.390 141.210 ;
        RECT 36.900 141.010 51.390 141.150 ;
        RECT 24.850 140.950 25.170 141.010 ;
        RECT 34.525 140.965 34.815 141.010 ;
        RECT 51.070 140.950 51.390 141.010 ;
        RECT 51.530 141.150 51.850 141.210 ;
        RECT 54.380 141.150 54.520 141.350 ;
        RECT 57.050 141.290 57.370 141.350 ;
        RECT 58.890 141.490 59.210 141.550 ;
        RECT 61.605 141.535 61.895 141.850 ;
        RECT 62.685 141.830 62.975 141.875 ;
        RECT 66.265 141.830 66.555 141.875 ;
        RECT 68.100 141.830 68.390 141.875 ;
        RECT 62.685 141.690 68.390 141.830 ;
        RECT 62.685 141.645 62.975 141.690 ;
        RECT 66.265 141.645 66.555 141.690 ;
        RECT 68.100 141.645 68.390 141.690 ;
        RECT 68.550 141.630 68.870 141.890 ;
        RECT 69.930 141.630 70.250 141.890 ;
        RECT 71.785 141.830 72.075 141.875 ;
        RECT 71.170 141.690 72.075 141.830 ;
        RECT 61.305 141.490 61.895 141.535 ;
        RECT 64.545 141.490 65.195 141.535 ;
        RECT 58.890 141.350 65.195 141.490 ;
        RECT 58.890 141.290 59.210 141.350 ;
        RECT 61.305 141.305 61.595 141.350 ;
        RECT 64.545 141.305 65.195 141.350 ;
        RECT 69.470 141.490 69.790 141.550 ;
        RECT 70.390 141.490 70.710 141.550 ;
        RECT 71.170 141.490 71.310 141.690 ;
        RECT 71.785 141.645 72.075 141.690 ;
        RECT 108.570 141.630 108.890 141.890 ;
        RECT 109.965 141.830 110.255 141.875 ;
        RECT 110.870 141.830 111.190 141.890 ;
        RECT 109.965 141.690 111.190 141.830 ;
        RECT 109.965 141.645 110.255 141.690 ;
        RECT 110.870 141.630 111.190 141.690 ;
        RECT 117.770 141.630 118.090 141.890 ;
        RECT 120.085 141.830 120.375 141.875 ;
        RECT 120.530 141.830 120.850 141.890 ;
        RECT 120.085 141.690 120.850 141.830 ;
        RECT 120.085 141.645 120.375 141.690 ;
        RECT 120.530 141.630 120.850 141.690 ;
        RECT 69.470 141.350 71.310 141.490 ;
        RECT 69.470 141.290 69.790 141.350 ;
        RECT 70.390 141.290 70.710 141.350 ;
        RECT 51.530 141.010 54.520 141.150 ;
        RECT 51.530 140.950 51.850 141.010 ;
        RECT 72.230 140.950 72.550 141.210 ;
        RECT 110.885 141.150 111.175 141.195 ;
        RECT 113.630 141.150 113.950 141.210 ;
        RECT 110.885 141.010 113.950 141.150 ;
        RECT 110.885 140.965 111.175 141.010 ;
        RECT 113.630 140.950 113.950 141.010 ;
        RECT 117.310 140.950 117.630 141.210 ;
        RECT 120.530 140.950 120.850 141.210 ;
        RECT 35.890 139.930 36.210 140.190 ;
        RECT 38.665 139.945 38.955 140.175 ;
        RECT 48.770 140.130 49.090 140.190 ;
        RECT 39.660 139.990 49.090 140.130 ;
        RECT 18.410 139.835 18.730 139.850 ;
        RECT 18.360 139.790 18.730 139.835 ;
        RECT 21.620 139.790 21.910 139.835 ;
        RECT 18.360 139.650 21.910 139.790 ;
        RECT 18.360 139.605 18.730 139.650 ;
        RECT 21.620 139.605 21.910 139.650 ;
        RECT 22.540 139.790 22.830 139.835 ;
        RECT 24.400 139.790 24.690 139.835 ;
        RECT 22.540 139.650 24.690 139.790 ;
        RECT 22.540 139.605 22.830 139.650 ;
        RECT 24.400 139.605 24.690 139.650 ;
        RECT 25.770 139.790 26.090 139.850 ;
        RECT 38.740 139.790 38.880 139.945 ;
        RECT 25.770 139.650 38.880 139.790 ;
        RECT 18.410 139.590 18.730 139.605 ;
        RECT 20.220 139.450 20.510 139.495 ;
        RECT 22.540 139.450 22.755 139.605 ;
        RECT 25.770 139.590 26.090 139.650 ;
        RECT 39.660 139.495 39.800 139.990 ;
        RECT 48.770 139.930 49.090 139.990 ;
        RECT 49.245 140.130 49.535 140.175 ;
        RECT 50.610 140.130 50.930 140.190 ;
        RECT 49.245 139.990 50.930 140.130 ;
        RECT 49.245 139.945 49.535 139.990 ;
        RECT 50.610 139.930 50.930 139.990 ;
        RECT 51.070 140.130 51.390 140.190 ;
        RECT 59.365 140.130 59.655 140.175 ;
        RECT 63.950 140.130 64.270 140.190 ;
        RECT 70.850 140.130 71.170 140.190 ;
        RECT 51.070 139.990 59.655 140.130 ;
        RECT 51.070 139.930 51.390 139.990 ;
        RECT 59.365 139.945 59.655 139.990 ;
        RECT 59.900 139.990 64.270 140.130 ;
        RECT 40.965 139.790 41.255 139.835 ;
        RECT 41.410 139.790 41.730 139.850 ;
        RECT 40.965 139.650 41.730 139.790 ;
        RECT 40.965 139.605 41.255 139.650 ;
        RECT 41.410 139.590 41.730 139.650 ;
        RECT 46.945 139.790 47.235 139.835 ;
        RECT 49.705 139.790 49.995 139.835 ;
        RECT 59.900 139.790 60.040 139.990 ;
        RECT 63.950 139.930 64.270 139.990 ;
        RECT 65.420 139.990 71.170 140.130 ;
        RECT 64.410 139.790 64.730 139.850 ;
        RECT 46.945 139.650 49.995 139.790 ;
        RECT 46.945 139.605 47.235 139.650 ;
        RECT 49.705 139.605 49.995 139.650 ;
        RECT 50.700 139.650 60.040 139.790 ;
        RECT 61.740 139.650 64.730 139.790 ;
        RECT 20.220 139.310 22.755 139.450 ;
        RECT 20.220 139.265 20.510 139.310 ;
        RECT 34.065 139.265 34.355 139.495 ;
        RECT 34.985 139.265 35.275 139.495 ;
        RECT 39.585 139.265 39.875 139.495 ;
        RECT 45.550 139.450 45.870 139.510 ;
        RECT 48.325 139.450 48.615 139.495 ;
        RECT 45.550 139.310 48.615 139.450 ;
        RECT 23.470 138.910 23.790 139.170 ;
        RECT 25.325 139.110 25.615 139.155 ;
        RECT 26.230 139.110 26.550 139.170 ;
        RECT 25.325 138.970 26.550 139.110 ;
        RECT 25.325 138.925 25.615 138.970 ;
        RECT 26.230 138.910 26.550 138.970 ;
        RECT 20.220 138.770 20.510 138.815 ;
        RECT 23.000 138.770 23.290 138.815 ;
        RECT 24.860 138.770 25.150 138.815 ;
        RECT 20.220 138.630 25.150 138.770 ;
        RECT 20.220 138.585 20.510 138.630 ;
        RECT 23.000 138.585 23.290 138.630 ;
        RECT 24.860 138.585 25.150 138.630 ;
        RECT 30.830 138.770 31.150 138.830 ;
        RECT 34.140 138.770 34.280 139.265 ;
        RECT 30.830 138.630 34.280 138.770 ;
        RECT 35.060 138.770 35.200 139.265 ;
        RECT 45.550 139.250 45.870 139.310 ;
        RECT 48.325 139.265 48.615 139.310 ;
        RECT 48.770 139.450 49.090 139.510 ;
        RECT 50.700 139.450 50.840 139.650 ;
        RECT 48.770 139.310 50.840 139.450 ;
        RECT 48.770 139.250 49.090 139.310 ;
        RECT 51.085 139.265 51.375 139.495 ;
        RECT 40.030 138.910 40.350 139.170 ;
        RECT 46.010 139.110 46.330 139.170 ;
        RECT 47.405 139.110 47.695 139.155 ;
        RECT 46.010 138.970 47.695 139.110 ;
        RECT 46.010 138.910 46.330 138.970 ;
        RECT 47.405 138.925 47.695 138.970 ;
        RECT 49.690 139.110 50.010 139.170 ;
        RECT 51.160 139.110 51.300 139.265 ;
        RECT 51.530 139.250 51.850 139.510 ;
        RECT 52.005 139.450 52.295 139.495 ;
        RECT 52.450 139.450 52.770 139.510 ;
        RECT 52.005 139.310 52.770 139.450 ;
        RECT 52.005 139.265 52.295 139.310 ;
        RECT 52.450 139.250 52.770 139.310 ;
        RECT 52.925 139.265 53.215 139.495 ;
        RECT 55.225 139.265 55.515 139.495 ;
        RECT 49.690 138.970 51.300 139.110 ;
        RECT 49.690 138.910 50.010 138.970 ;
        RECT 41.410 138.770 41.730 138.830 ;
        RECT 35.060 138.630 41.730 138.770 ;
        RECT 30.830 138.570 31.150 138.630 ;
        RECT 41.410 138.570 41.730 138.630 ;
        RECT 48.770 138.770 49.090 138.830 ;
        RECT 53.000 138.770 53.140 139.265 ;
        RECT 55.300 139.110 55.440 139.265 ;
        RECT 55.670 139.250 55.990 139.510 ;
        RECT 61.740 139.495 61.880 139.650 ;
        RECT 64.410 139.590 64.730 139.650 ;
        RECT 64.870 139.590 65.190 139.850 ;
        RECT 60.745 139.265 61.035 139.495 ;
        RECT 61.205 139.265 61.495 139.495 ;
        RECT 61.665 139.265 61.955 139.495 ;
        RECT 62.585 139.450 62.875 139.495 ;
        RECT 64.960 139.450 65.100 139.590 ;
        RECT 65.420 139.510 65.560 139.990 ;
        RECT 70.850 139.930 71.170 139.990 ;
        RECT 86.030 139.930 86.350 140.190 ;
        RECT 88.345 139.945 88.635 140.175 ;
        RECT 99.370 140.130 99.690 140.190 ;
        RECT 110.870 140.130 111.190 140.190 ;
        RECT 99.370 139.990 111.190 140.130 ;
        RECT 68.090 139.790 68.410 139.850 ;
        RECT 65.880 139.650 68.410 139.790 ;
        RECT 62.585 139.310 65.100 139.450 ;
        RECT 62.585 139.265 62.875 139.310 ;
        RECT 56.130 139.110 56.450 139.170 ;
        RECT 55.300 138.970 56.450 139.110 ;
        RECT 56.130 138.910 56.450 138.970 ;
        RECT 55.210 138.770 55.530 138.830 ;
        RECT 48.770 138.630 55.530 138.770 ;
        RECT 60.820 138.770 60.960 139.265 ;
        RECT 61.280 139.110 61.420 139.265 ;
        RECT 65.330 139.250 65.650 139.510 ;
        RECT 65.880 139.495 66.020 139.650 ;
        RECT 68.090 139.590 68.410 139.650 ;
        RECT 68.570 139.790 68.860 139.835 ;
        RECT 70.430 139.790 70.720 139.835 ;
        RECT 68.570 139.650 70.720 139.790 ;
        RECT 68.570 139.605 68.860 139.650 ;
        RECT 70.430 139.605 70.720 139.650 ;
        RECT 71.350 139.790 71.640 139.835 ;
        RECT 72.230 139.790 72.550 139.850 ;
        RECT 74.610 139.790 74.900 139.835 ;
        RECT 86.120 139.790 86.260 139.930 ;
        RECT 71.350 139.650 74.900 139.790 ;
        RECT 71.350 139.605 71.640 139.650 ;
        RECT 65.805 139.265 66.095 139.495 ;
        RECT 64.870 139.110 65.190 139.170 ;
        RECT 65.880 139.110 66.020 139.265 ;
        RECT 66.250 139.250 66.570 139.510 ;
        RECT 67.170 139.250 67.490 139.510 ;
        RECT 70.505 139.450 70.720 139.605 ;
        RECT 72.230 139.590 72.550 139.650 ;
        RECT 74.610 139.605 74.900 139.650 ;
        RECT 82.440 139.650 86.260 139.790 ;
        RECT 72.750 139.450 73.040 139.495 ;
        RECT 70.505 139.310 73.040 139.450 ;
        RECT 72.750 139.265 73.040 139.310 ;
        RECT 81.430 139.250 81.750 139.510 ;
        RECT 81.890 139.250 82.210 139.510 ;
        RECT 82.440 139.495 82.580 139.650 ;
        RECT 83.270 139.495 83.590 139.510 ;
        RECT 82.365 139.265 82.655 139.495 ;
        RECT 83.255 139.450 83.590 139.495 ;
        RECT 83.075 139.310 83.590 139.450 ;
        RECT 83.255 139.265 83.590 139.310 ;
        RECT 86.505 139.265 86.795 139.495 ;
        RECT 88.420 139.450 88.560 139.945 ;
        RECT 99.370 139.930 99.690 139.990 ;
        RECT 100.290 139.790 100.610 139.850 ;
        RECT 105.810 139.790 106.130 139.850 ;
        RECT 106.285 139.790 106.575 139.835 ;
        RECT 100.290 139.650 105.120 139.790 ;
        RECT 100.290 139.590 100.610 139.650 ;
        RECT 89.725 139.450 90.015 139.495 ;
        RECT 88.420 139.310 90.015 139.450 ;
        RECT 89.725 139.265 90.015 139.310 ;
        RECT 83.270 139.250 83.590 139.265 ;
        RECT 61.280 138.970 66.020 139.110 ;
        RECT 67.645 139.110 67.935 139.155 ;
        RECT 68.550 139.110 68.870 139.170 ;
        RECT 67.645 138.970 68.870 139.110 ;
        RECT 64.870 138.910 65.190 138.970 ;
        RECT 67.645 138.925 67.935 138.970 ;
        RECT 68.550 138.910 68.870 138.970 ;
        RECT 69.470 138.910 69.790 139.170 ;
        RECT 70.850 139.110 71.170 139.170 ;
        RECT 70.850 138.970 83.040 139.110 ;
        RECT 70.850 138.910 71.170 138.970 ;
        RECT 65.330 138.770 65.650 138.830 ;
        RECT 60.820 138.630 65.650 138.770 ;
        RECT 48.770 138.570 49.090 138.630 ;
        RECT 55.210 138.570 55.530 138.630 ;
        RECT 65.330 138.570 65.650 138.630 ;
        RECT 68.110 138.770 68.400 138.815 ;
        RECT 69.970 138.770 70.260 138.815 ;
        RECT 72.750 138.770 73.040 138.815 ;
        RECT 68.110 138.630 73.040 138.770 ;
        RECT 82.900 138.770 83.040 138.970 ;
        RECT 85.110 138.910 85.430 139.170 ;
        RECT 86.580 139.110 86.720 139.265 ;
        RECT 101.210 139.250 101.530 139.510 ;
        RECT 101.670 139.250 101.990 139.510 ;
        RECT 104.980 139.450 105.120 139.650 ;
        RECT 105.810 139.650 106.575 139.790 ;
        RECT 105.810 139.590 106.130 139.650 ;
        RECT 106.285 139.605 106.575 139.650 ;
        RECT 108.200 139.495 108.340 139.990 ;
        RECT 110.870 139.930 111.190 139.990 ;
        RECT 111.330 139.930 111.650 140.190 ;
        RECT 120.990 140.130 121.310 140.190 ;
        RECT 118.780 139.990 121.310 140.130 ;
        RECT 111.420 139.790 111.560 139.930 ;
        RECT 112.250 139.790 112.570 139.850 ;
        RECT 113.185 139.790 113.475 139.835 ;
        RECT 110.500 139.650 112.020 139.790 ;
        RECT 107.665 139.450 107.955 139.495 ;
        RECT 104.980 139.310 107.955 139.450 ;
        RECT 107.665 139.265 107.955 139.310 ;
        RECT 108.125 139.265 108.415 139.495 ;
        RECT 90.630 139.110 90.950 139.170 ;
        RECT 86.580 138.970 90.950 139.110 ;
        RECT 101.300 139.110 101.440 139.250 ;
        RECT 107.740 139.110 107.880 139.265 ;
        RECT 108.570 139.250 108.890 139.510 ;
        RECT 109.030 139.450 109.350 139.510 ;
        RECT 109.505 139.450 109.795 139.495 ;
        RECT 109.965 139.450 110.255 139.495 ;
        RECT 109.030 139.310 110.255 139.450 ;
        RECT 109.030 139.250 109.350 139.310 ;
        RECT 109.505 139.265 109.795 139.310 ;
        RECT 109.965 139.265 110.255 139.310 ;
        RECT 110.500 139.110 110.640 139.650 ;
        RECT 110.885 139.265 111.175 139.495 ;
        RECT 101.300 138.970 101.900 139.110 ;
        RECT 107.740 138.970 110.640 139.110 ;
        RECT 110.960 139.110 111.100 139.265 ;
        RECT 111.330 139.250 111.650 139.510 ;
        RECT 111.880 139.495 112.020 139.650 ;
        RECT 112.250 139.650 113.475 139.790 ;
        RECT 112.250 139.590 112.570 139.650 ;
        RECT 113.185 139.605 113.475 139.650 ;
        RECT 111.805 139.265 112.095 139.495 ;
        RECT 115.485 139.265 115.775 139.495 ;
        RECT 115.560 139.110 115.700 139.265 ;
        RECT 115.930 139.250 116.250 139.510 ;
        RECT 118.780 139.110 118.920 139.990 ;
        RECT 120.990 139.930 121.310 139.990 ;
        RECT 119.100 139.790 119.390 139.835 ;
        RECT 120.530 139.790 120.850 139.850 ;
        RECT 122.360 139.790 122.650 139.835 ;
        RECT 119.100 139.650 122.650 139.790 ;
        RECT 119.100 139.605 119.390 139.650 ;
        RECT 120.530 139.590 120.850 139.650 ;
        RECT 122.360 139.605 122.650 139.650 ;
        RECT 123.280 139.790 123.570 139.835 ;
        RECT 125.140 139.790 125.430 139.835 ;
        RECT 123.280 139.650 125.430 139.790 ;
        RECT 123.280 139.605 123.570 139.650 ;
        RECT 125.140 139.605 125.430 139.650 ;
        RECT 120.960 139.450 121.250 139.495 ;
        RECT 123.280 139.450 123.495 139.605 ;
        RECT 120.960 139.310 123.495 139.450 ;
        RECT 120.960 139.265 121.250 139.310 ;
        RECT 110.960 138.970 111.560 139.110 ;
        RECT 115.560 138.970 118.920 139.110 ;
        RECT 90.630 138.910 90.950 138.970 ;
        RECT 100.290 138.770 100.610 138.830 ;
        RECT 82.900 138.630 100.610 138.770 ;
        RECT 68.110 138.585 68.400 138.630 ;
        RECT 69.970 138.585 70.260 138.630 ;
        RECT 72.750 138.585 73.040 138.630 ;
        RECT 100.290 138.570 100.610 138.630 ;
        RECT 16.355 138.430 16.645 138.475 ;
        RECT 19.330 138.430 19.650 138.490 ;
        RECT 16.355 138.290 19.650 138.430 ;
        RECT 16.355 138.245 16.645 138.290 ;
        RECT 19.330 138.230 19.650 138.290 ;
        RECT 39.570 138.230 39.890 138.490 ;
        RECT 45.550 138.430 45.870 138.490 ;
        RECT 46.945 138.430 47.235 138.475 ;
        RECT 45.550 138.290 47.235 138.430 ;
        RECT 45.550 138.230 45.870 138.290 ;
        RECT 46.945 138.245 47.235 138.290 ;
        RECT 64.410 138.430 64.730 138.490 ;
        RECT 70.850 138.430 71.170 138.490 ;
        RECT 76.615 138.430 76.905 138.475 ;
        RECT 64.410 138.290 76.905 138.430 ;
        RECT 64.410 138.230 64.730 138.290 ;
        RECT 70.850 138.230 71.170 138.290 ;
        RECT 76.615 138.245 76.905 138.290 ;
        RECT 79.590 138.430 79.910 138.490 ;
        RECT 80.065 138.430 80.355 138.475 ;
        RECT 79.590 138.290 80.355 138.430 ;
        RECT 79.590 138.230 79.910 138.290 ;
        RECT 80.065 138.245 80.355 138.290 ;
        RECT 90.645 138.430 90.935 138.475 ;
        RECT 91.090 138.430 91.410 138.490 ;
        RECT 90.645 138.290 91.410 138.430 ;
        RECT 90.645 138.245 90.935 138.290 ;
        RECT 91.090 138.230 91.410 138.290 ;
        RECT 94.310 138.430 94.630 138.490 ;
        RECT 101.760 138.430 101.900 138.970 ;
        RECT 111.420 138.830 111.560 138.970 ;
        RECT 124.210 138.910 124.530 139.170 ;
        RECT 126.050 138.910 126.370 139.170 ;
        RECT 111.330 138.770 111.650 138.830 ;
        RECT 117.310 138.815 117.630 138.830 ;
        RECT 117.095 138.770 117.630 138.815 ;
        RECT 111.330 138.630 117.630 138.770 ;
        RECT 111.330 138.570 111.650 138.630 ;
        RECT 117.095 138.585 117.630 138.630 ;
        RECT 120.960 138.770 121.250 138.815 ;
        RECT 123.740 138.770 124.030 138.815 ;
        RECT 125.600 138.770 125.890 138.815 ;
        RECT 120.960 138.630 125.890 138.770 ;
        RECT 120.960 138.585 121.250 138.630 ;
        RECT 123.740 138.585 124.030 138.630 ;
        RECT 125.600 138.585 125.890 138.630 ;
        RECT 117.310 138.570 117.630 138.585 ;
        RECT 116.390 138.430 116.710 138.490 ;
        RECT 94.310 138.290 116.710 138.430 ;
        RECT 94.310 138.230 94.630 138.290 ;
        RECT 116.390 138.230 116.710 138.290 ;
        RECT 22.565 137.410 22.855 137.455 ;
        RECT 23.470 137.410 23.790 137.470 ;
        RECT 22.565 137.270 23.790 137.410 ;
        RECT 22.565 137.225 22.855 137.270 ;
        RECT 23.470 137.210 23.790 137.270 ;
        RECT 37.270 137.210 37.590 137.470 ;
        RECT 39.570 137.210 39.890 137.470 ;
        RECT 44.170 137.410 44.490 137.470 ;
        RECT 44.645 137.410 44.935 137.455 ;
        RECT 65.330 137.410 65.650 137.470 ;
        RECT 44.170 137.270 44.935 137.410 ;
        RECT 44.170 137.210 44.490 137.270 ;
        RECT 44.645 137.225 44.935 137.270 ;
        RECT 63.580 137.270 65.650 137.410 ;
        RECT 39.110 137.070 39.430 137.130 ;
        RECT 35.980 136.930 39.430 137.070 ;
        RECT 29.925 136.730 30.215 136.775 ;
        RECT 34.050 136.730 34.370 136.790 ;
        RECT 29.925 136.590 34.370 136.730 ;
        RECT 29.925 136.545 30.215 136.590 ;
        RECT 34.050 136.530 34.370 136.590 ;
        RECT 21.170 136.390 21.490 136.450 ;
        RECT 21.645 136.390 21.935 136.435 ;
        RECT 21.170 136.250 21.935 136.390 ;
        RECT 21.170 136.190 21.490 136.250 ;
        RECT 21.645 136.205 21.935 136.250 ;
        RECT 23.025 136.390 23.315 136.435 ;
        RECT 23.470 136.390 23.790 136.450 ;
        RECT 35.980 136.435 36.120 136.930 ;
        RECT 39.110 136.870 39.430 136.930 ;
        RECT 56.605 136.885 56.895 137.115 ;
        RECT 36.350 136.530 36.670 136.790 ;
        RECT 45.565 136.730 45.855 136.775 ;
        RECT 46.470 136.730 46.790 136.790 ;
        RECT 37.360 136.590 45.320 136.730 ;
        RECT 37.360 136.435 37.500 136.590 ;
        RECT 23.025 136.250 23.790 136.390 ;
        RECT 23.025 136.205 23.315 136.250 ;
        RECT 17.030 136.050 17.350 136.110 ;
        RECT 23.100 136.050 23.240 136.205 ;
        RECT 23.470 136.190 23.790 136.250 ;
        RECT 35.905 136.205 36.195 136.435 ;
        RECT 37.285 136.205 37.575 136.435 ;
        RECT 37.745 136.205 38.035 136.435 ;
        RECT 38.665 136.390 38.955 136.435 ;
        RECT 41.410 136.390 41.730 136.450 ;
        RECT 38.665 136.250 41.730 136.390 ;
        RECT 38.665 136.205 38.955 136.250 ;
        RECT 37.820 136.050 37.960 136.205 ;
        RECT 41.410 136.190 41.730 136.250 ;
        RECT 44.630 136.190 44.950 136.450 ;
        RECT 45.180 136.390 45.320 136.590 ;
        RECT 45.565 136.590 46.790 136.730 ;
        RECT 45.565 136.545 45.855 136.590 ;
        RECT 46.470 136.530 46.790 136.590 ;
        RECT 53.845 136.730 54.135 136.775 ;
        RECT 54.290 136.730 54.610 136.790 ;
        RECT 53.845 136.590 54.610 136.730 ;
        RECT 53.845 136.545 54.135 136.590 ;
        RECT 54.290 136.530 54.610 136.590 ;
        RECT 47.850 136.390 48.170 136.450 ;
        RECT 45.180 136.250 48.170 136.390 ;
        RECT 47.850 136.190 48.170 136.250 ;
        RECT 52.450 136.390 52.770 136.450 ;
        RECT 54.765 136.390 55.055 136.435 ;
        RECT 52.450 136.250 55.055 136.390 ;
        RECT 56.680 136.390 56.820 136.885 ;
        RECT 63.580 136.730 63.720 137.270 ;
        RECT 65.330 137.210 65.650 137.270 ;
        RECT 67.185 137.410 67.475 137.455 ;
        RECT 69.470 137.410 69.790 137.470 ;
        RECT 67.185 137.270 69.790 137.410 ;
        RECT 67.185 137.225 67.475 137.270 ;
        RECT 69.470 137.210 69.790 137.270 ;
        RECT 78.670 137.210 78.990 137.470 ;
        RECT 83.975 137.410 84.265 137.455 ;
        RECT 86.030 137.410 86.350 137.470 ;
        RECT 97.990 137.410 98.310 137.470 ;
        RECT 107.650 137.410 107.970 137.470 ;
        RECT 109.030 137.410 109.350 137.470 ;
        RECT 83.975 137.270 86.350 137.410 ;
        RECT 83.975 137.225 84.265 137.270 ;
        RECT 86.030 137.210 86.350 137.270 ;
        RECT 87.500 137.270 109.350 137.410 ;
        RECT 63.950 136.870 64.270 137.130 ;
        RECT 65.790 137.070 66.110 137.130 ;
        RECT 87.500 137.070 87.640 137.270 ;
        RECT 97.990 137.210 98.310 137.270 ;
        RECT 107.650 137.210 107.970 137.270 ;
        RECT 109.030 137.210 109.350 137.270 ;
        RECT 124.210 137.210 124.530 137.470 ;
        RECT 65.790 136.930 87.640 137.070 ;
        RECT 87.840 137.070 88.130 137.115 ;
        RECT 90.620 137.070 90.910 137.115 ;
        RECT 92.480 137.070 92.770 137.115 ;
        RECT 87.840 136.930 92.770 137.070 ;
        RECT 65.790 136.870 66.110 136.930 ;
        RECT 87.840 136.885 88.130 136.930 ;
        RECT 90.620 136.885 90.910 136.930 ;
        RECT 92.480 136.885 92.770 136.930 ;
        RECT 106.745 136.885 107.035 137.115 ;
        RECT 62.660 136.590 63.720 136.730 ;
        RECT 64.040 136.730 64.180 136.870 ;
        RECT 70.850 136.730 71.170 136.790 ;
        RECT 73.165 136.730 73.455 136.775 ;
        RECT 64.040 136.590 68.320 136.730 ;
        RECT 62.660 136.435 62.800 136.590 ;
        RECT 57.525 136.390 57.815 136.435 ;
        RECT 56.680 136.250 57.815 136.390 ;
        RECT 52.450 136.190 52.770 136.250 ;
        RECT 54.765 136.205 55.055 136.250 ;
        RECT 57.525 136.205 57.815 136.250 ;
        RECT 62.585 136.205 62.875 136.435 ;
        RECT 63.045 136.205 63.335 136.435 ;
        RECT 63.505 136.390 63.795 136.435 ;
        RECT 63.950 136.390 64.270 136.450 ;
        RECT 63.505 136.250 64.270 136.390 ;
        RECT 63.505 136.205 63.795 136.250 ;
        RECT 17.030 135.910 23.240 136.050 ;
        RECT 30.460 135.910 37.960 136.050 ;
        RECT 40.030 136.050 40.350 136.110 ;
        RECT 40.030 135.910 45.780 136.050 ;
        RECT 17.030 135.850 17.350 135.910 ;
        RECT 30.460 135.770 30.600 135.910 ;
        RECT 40.030 135.850 40.350 135.910 ;
        RECT 23.485 135.710 23.775 135.755 ;
        RECT 23.930 135.710 24.250 135.770 ;
        RECT 23.485 135.570 24.250 135.710 ;
        RECT 23.485 135.525 23.775 135.570 ;
        RECT 23.930 135.510 24.250 135.570 ;
        RECT 30.370 135.510 30.690 135.770 ;
        RECT 30.830 135.510 31.150 135.770 ;
        RECT 32.670 135.510 32.990 135.770 ;
        RECT 34.985 135.710 35.275 135.755 ;
        RECT 35.430 135.710 35.750 135.770 ;
        RECT 34.985 135.570 35.750 135.710 ;
        RECT 34.985 135.525 35.275 135.570 ;
        RECT 35.430 135.510 35.750 135.570 ;
        RECT 42.330 135.710 42.650 135.770 ;
        RECT 43.725 135.710 44.015 135.755 ;
        RECT 42.330 135.570 44.015 135.710 ;
        RECT 45.640 135.710 45.780 135.910 ;
        RECT 46.010 135.850 46.330 136.110 ;
        RECT 61.205 136.050 61.495 136.095 ;
        RECT 50.700 135.910 61.495 136.050 ;
        RECT 63.120 136.050 63.260 136.205 ;
        RECT 63.950 136.190 64.270 136.250 ;
        RECT 64.425 136.390 64.715 136.435 ;
        RECT 65.790 136.390 66.110 136.450 ;
        RECT 68.180 136.435 68.320 136.590 ;
        RECT 70.850 136.590 73.455 136.730 ;
        RECT 70.850 136.530 71.170 136.590 ;
        RECT 73.165 136.545 73.455 136.590 ;
        RECT 79.130 136.530 79.450 136.790 ;
        RECT 85.110 136.730 85.430 136.790 ;
        RECT 85.110 136.590 90.860 136.730 ;
        RECT 85.110 136.530 85.430 136.590 ;
        RECT 64.425 136.250 66.110 136.390 ;
        RECT 64.425 136.205 64.715 136.250 ;
        RECT 65.790 136.190 66.110 136.250 ;
        RECT 68.105 136.205 68.395 136.435 ;
        RECT 69.010 136.190 69.330 136.450 ;
        RECT 69.945 136.390 70.235 136.435 ;
        RECT 70.405 136.390 70.695 136.435 ;
        RECT 69.945 136.250 70.695 136.390 ;
        RECT 69.945 136.205 70.235 136.250 ;
        RECT 70.405 136.205 70.695 136.250 ;
        RECT 76.830 136.390 77.150 136.450 ;
        RECT 78.225 136.390 78.515 136.435 ;
        RECT 76.830 136.250 78.515 136.390 ;
        RECT 76.830 136.190 77.150 136.250 ;
        RECT 78.225 136.205 78.515 136.250 ;
        RECT 79.590 136.190 79.910 136.450 ;
        RECT 81.430 136.190 81.750 136.450 ;
        RECT 81.890 136.190 82.210 136.450 ;
        RECT 82.365 136.205 82.655 136.435 ;
        RECT 64.870 136.050 65.190 136.110 ;
        RECT 63.120 135.910 65.190 136.050 ;
        RECT 50.700 135.710 50.840 135.910 ;
        RECT 61.205 135.865 61.495 135.910 ;
        RECT 64.870 135.850 65.190 135.910 ;
        RECT 68.565 136.050 68.855 136.095 ;
        RECT 74.070 136.050 74.390 136.110 ;
        RECT 68.565 135.910 74.390 136.050 ;
        RECT 68.565 135.865 68.855 135.910 ;
        RECT 74.070 135.850 74.390 135.910 ;
        RECT 45.640 135.570 50.840 135.710 ;
        RECT 42.330 135.510 42.650 135.570 ;
        RECT 43.725 135.525 44.015 135.570 ;
        RECT 54.290 135.510 54.610 135.770 ;
        RECT 58.445 135.710 58.735 135.755 ;
        RECT 60.270 135.710 60.590 135.770 ;
        RECT 58.445 135.570 60.590 135.710 ;
        RECT 58.445 135.525 58.735 135.570 ;
        RECT 60.270 135.510 60.590 135.570 ;
        RECT 77.305 135.710 77.595 135.755 ;
        RECT 77.750 135.710 78.070 135.770 ;
        RECT 77.305 135.570 78.070 135.710 ;
        RECT 77.305 135.525 77.595 135.570 ;
        RECT 77.750 135.510 78.070 135.570 ;
        RECT 79.130 135.710 79.450 135.770 ;
        RECT 80.065 135.710 80.355 135.755 ;
        RECT 79.130 135.570 80.355 135.710 ;
        RECT 82.440 135.710 82.580 136.205 ;
        RECT 83.270 136.190 83.590 136.450 ;
        RECT 87.840 136.390 88.130 136.435 ;
        RECT 90.720 136.390 90.860 136.590 ;
        RECT 91.090 136.530 91.410 136.790 ;
        RECT 92.945 136.730 93.235 136.775 ;
        RECT 93.850 136.730 94.170 136.790 ;
        RECT 92.945 136.590 94.170 136.730 ;
        RECT 92.945 136.545 93.235 136.590 ;
        RECT 93.850 136.530 94.170 136.590 ;
        RECT 94.325 136.730 94.615 136.775 ;
        RECT 103.510 136.730 103.830 136.790 ;
        RECT 94.325 136.590 103.830 136.730 ;
        RECT 94.325 136.545 94.615 136.590 ;
        RECT 94.400 136.390 94.540 136.545 ;
        RECT 103.510 136.530 103.830 136.590 ;
        RECT 87.840 136.250 90.375 136.390 ;
        RECT 90.720 136.250 94.540 136.390 ;
        RECT 87.840 136.205 88.130 136.250 ;
        RECT 85.980 136.050 86.270 136.095 ;
        RECT 87.410 136.050 87.730 136.110 ;
        RECT 90.160 136.095 90.375 136.250 ;
        RECT 95.245 136.205 95.535 136.435 ;
        RECT 89.240 136.050 89.530 136.095 ;
        RECT 85.980 135.910 89.530 136.050 ;
        RECT 85.980 135.865 86.270 135.910 ;
        RECT 87.410 135.850 87.730 135.910 ;
        RECT 89.240 135.865 89.530 135.910 ;
        RECT 90.160 136.050 90.450 136.095 ;
        RECT 92.020 136.050 92.310 136.095 ;
        RECT 90.160 135.910 92.310 136.050 ;
        RECT 95.320 136.050 95.460 136.205 ;
        RECT 97.990 136.190 98.310 136.450 ;
        RECT 98.925 136.205 99.215 136.435 ;
        RECT 98.450 136.050 98.770 136.110 ;
        RECT 99.000 136.050 99.140 136.205 ;
        RECT 99.370 136.190 99.690 136.450 ;
        RECT 99.845 136.390 100.135 136.435 ;
        RECT 100.290 136.390 100.610 136.450 ;
        RECT 99.845 136.250 100.610 136.390 ;
        RECT 106.820 136.390 106.960 136.885 ;
        RECT 113.170 136.870 113.490 137.130 ;
        RECT 117.740 137.070 118.030 137.115 ;
        RECT 120.520 137.070 120.810 137.115 ;
        RECT 122.380 137.070 122.670 137.115 ;
        RECT 117.740 136.930 122.670 137.070 ;
        RECT 117.740 136.885 118.030 136.930 ;
        RECT 120.520 136.885 120.810 136.930 ;
        RECT 122.380 136.885 122.670 136.930 ;
        RECT 109.030 136.730 109.350 136.790 ;
        RECT 109.965 136.730 110.255 136.775 ;
        RECT 112.710 136.730 113.030 136.790 ;
        RECT 122.845 136.730 123.135 136.775 ;
        RECT 126.050 136.730 126.370 136.790 ;
        RECT 109.030 136.590 113.030 136.730 ;
        RECT 109.030 136.530 109.350 136.590 ;
        RECT 109.965 136.545 110.255 136.590 ;
        RECT 112.710 136.530 113.030 136.590 ;
        RECT 117.400 136.590 126.370 136.730 ;
        RECT 106.820 136.370 107.420 136.390 ;
        RECT 108.005 136.370 108.295 136.415 ;
        RECT 106.820 136.250 108.295 136.370 ;
        RECT 99.845 136.205 100.135 136.250 ;
        RECT 100.290 136.190 100.610 136.250 ;
        RECT 107.280 136.230 108.295 136.250 ;
        RECT 108.005 136.185 108.295 136.230 ;
        RECT 111.330 136.190 111.650 136.450 ;
        RECT 111.790 136.390 112.110 136.450 ;
        RECT 117.400 136.390 117.540 136.590 ;
        RECT 122.845 136.545 123.135 136.590 ;
        RECT 126.050 136.530 126.370 136.590 ;
        RECT 111.790 136.250 117.540 136.390 ;
        RECT 117.740 136.390 118.030 136.435 ;
        RECT 117.740 136.250 120.275 136.390 ;
        RECT 111.790 136.190 112.110 136.250 ;
        RECT 117.740 136.205 118.030 136.250 ;
        RECT 104.445 136.050 104.735 136.095 ;
        RECT 95.320 135.910 104.735 136.050 ;
        RECT 90.160 135.865 90.450 135.910 ;
        RECT 92.020 135.865 92.310 135.910 ;
        RECT 98.450 135.850 98.770 135.910 ;
        RECT 104.445 135.865 104.735 135.910 ;
        RECT 104.905 136.050 105.195 136.095 ;
        RECT 108.570 136.050 108.890 136.110 ;
        RECT 115.930 136.095 116.250 136.110 ;
        RECT 120.060 136.095 120.275 136.250 ;
        RECT 120.990 136.190 121.310 136.450 ;
        RECT 123.305 136.390 123.595 136.435 ;
        RECT 124.670 136.390 124.990 136.450 ;
        RECT 123.305 136.250 124.990 136.390 ;
        RECT 123.305 136.205 123.595 136.250 ;
        RECT 124.670 136.190 124.990 136.250 ;
        RECT 110.885 136.050 111.175 136.095 ;
        RECT 113.875 136.050 114.165 136.095 ;
        RECT 104.905 135.910 107.880 136.050 ;
        RECT 104.905 135.865 105.195 135.910 ;
        RECT 90.630 135.710 90.950 135.770 ;
        RECT 94.785 135.710 95.075 135.755 ;
        RECT 82.440 135.570 95.075 135.710 ;
        RECT 79.130 135.510 79.450 135.570 ;
        RECT 80.065 135.525 80.355 135.570 ;
        RECT 90.630 135.510 90.950 135.570 ;
        RECT 94.785 135.525 95.075 135.570 ;
        RECT 95.230 135.710 95.550 135.770 ;
        RECT 97.085 135.710 97.375 135.755 ;
        RECT 95.230 135.570 97.375 135.710 ;
        RECT 95.230 135.510 95.550 135.570 ;
        RECT 97.085 135.525 97.375 135.570 ;
        RECT 101.210 135.510 101.530 135.770 ;
        RECT 106.270 135.710 106.590 135.770 ;
        RECT 107.205 135.710 107.495 135.755 ;
        RECT 106.270 135.570 107.495 135.710 ;
        RECT 107.740 135.710 107.880 135.910 ;
        RECT 108.570 135.910 114.165 136.050 ;
        RECT 108.570 135.850 108.890 135.910 ;
        RECT 110.885 135.865 111.175 135.910 ;
        RECT 113.875 135.865 114.165 135.910 ;
        RECT 115.880 136.050 116.250 136.095 ;
        RECT 119.140 136.050 119.430 136.095 ;
        RECT 115.880 135.910 119.430 136.050 ;
        RECT 115.880 135.865 116.250 135.910 ;
        RECT 119.140 135.865 119.430 135.910 ;
        RECT 120.060 136.050 120.350 136.095 ;
        RECT 121.920 136.050 122.210 136.095 ;
        RECT 120.060 135.910 122.210 136.050 ;
        RECT 120.060 135.865 120.350 135.910 ;
        RECT 121.920 135.865 122.210 135.910 ;
        RECT 115.930 135.850 116.250 135.865 ;
        RECT 108.660 135.710 108.800 135.850 ;
        RECT 107.740 135.570 108.800 135.710 ;
        RECT 106.270 135.510 106.590 135.570 ;
        RECT 107.205 135.525 107.495 135.570 ;
        RECT 16.585 134.690 16.875 134.735 ;
        RECT 18.410 134.690 18.730 134.750 ;
        RECT 16.585 134.550 18.730 134.690 ;
        RECT 16.585 134.505 16.875 134.550 ;
        RECT 18.410 134.490 18.730 134.550 ;
        RECT 19.330 134.490 19.650 134.750 ;
        RECT 21.170 134.490 21.490 134.750 ;
        RECT 30.830 134.690 31.150 134.750 ;
        RECT 22.870 134.550 31.150 134.690 ;
        RECT 18.885 134.350 19.175 134.395 ;
        RECT 21.875 134.350 22.165 134.395 ;
        RECT 22.870 134.350 23.010 134.550 ;
        RECT 30.830 134.490 31.150 134.550 ;
        RECT 31.305 134.505 31.595 134.735 ;
        RECT 44.645 134.690 44.935 134.735 ;
        RECT 46.010 134.690 46.330 134.750 ;
        RECT 44.645 134.550 46.330 134.690 ;
        RECT 44.645 134.505 44.935 134.550 ;
        RECT 23.930 134.395 24.250 134.410 ;
        RECT 18.885 134.210 23.010 134.350 ;
        RECT 23.880 134.350 24.250 134.395 ;
        RECT 27.140 134.350 27.430 134.395 ;
        RECT 23.880 134.210 27.430 134.350 ;
        RECT 18.885 134.165 19.175 134.210 ;
        RECT 21.875 134.165 22.165 134.210 ;
        RECT 23.880 134.165 24.250 134.210 ;
        RECT 27.140 134.165 27.430 134.210 ;
        RECT 28.060 134.350 28.350 134.395 ;
        RECT 29.920 134.350 30.210 134.395 ;
        RECT 28.060 134.210 30.210 134.350 ;
        RECT 28.060 134.165 28.350 134.210 ;
        RECT 29.920 134.165 30.210 134.210 ;
        RECT 23.930 134.150 24.250 134.165 ;
        RECT 17.030 133.810 17.350 134.070 ;
        RECT 25.740 134.010 26.030 134.055 ;
        RECT 28.060 134.010 28.275 134.165 ;
        RECT 25.740 133.870 28.275 134.010 ;
        RECT 29.005 134.010 29.295 134.055 ;
        RECT 31.380 134.010 31.520 134.505 ;
        RECT 46.010 134.490 46.330 134.550 ;
        RECT 47.850 134.690 48.170 134.750 ;
        RECT 63.505 134.690 63.795 134.735 ;
        RECT 47.850 134.550 63.795 134.690 ;
        RECT 47.850 134.490 48.170 134.550 ;
        RECT 63.505 134.505 63.795 134.550 ;
        RECT 65.330 134.490 65.650 134.750 ;
        RECT 65.790 134.490 66.110 134.750 ;
        RECT 87.410 134.690 87.730 134.750 ;
        RECT 87.885 134.690 88.175 134.735 ;
        RECT 87.410 134.550 88.175 134.690 ;
        RECT 87.410 134.490 87.730 134.550 ;
        RECT 87.885 134.505 88.175 134.550 ;
        RECT 89.495 134.690 89.785 134.735 ;
        RECT 90.170 134.690 90.490 134.750 ;
        RECT 89.495 134.550 90.490 134.690 ;
        RECT 89.495 134.505 89.785 134.550 ;
        RECT 90.170 134.490 90.490 134.550 ;
        RECT 92.010 134.690 92.330 134.750 ;
        RECT 94.310 134.690 94.630 134.750 ;
        RECT 92.010 134.550 94.630 134.690 ;
        RECT 92.010 134.490 92.330 134.550 ;
        RECT 94.310 134.490 94.630 134.550 ;
        RECT 120.085 134.690 120.375 134.735 ;
        RECT 120.990 134.690 121.310 134.750 ;
        RECT 120.085 134.550 121.310 134.690 ;
        RECT 120.085 134.505 120.375 134.550 ;
        RECT 120.990 134.490 121.310 134.550 ;
        RECT 31.750 134.350 32.070 134.410 ;
        RECT 34.985 134.350 35.275 134.395 ;
        RECT 31.750 134.210 35.275 134.350 ;
        RECT 31.750 134.150 32.070 134.210 ;
        RECT 34.985 134.165 35.275 134.210 ;
        RECT 38.190 134.350 38.510 134.410 ;
        RECT 38.190 134.210 39.340 134.350 ;
        RECT 38.190 134.150 38.510 134.210 ;
        RECT 29.005 133.870 31.520 134.010 ;
        RECT 32.225 134.010 32.515 134.055 ;
        RECT 32.670 134.010 32.990 134.070 ;
        RECT 36.350 134.010 36.670 134.070 ;
        RECT 32.225 133.870 32.990 134.010 ;
        RECT 25.740 133.825 26.030 133.870 ;
        RECT 29.005 133.825 29.295 133.870 ;
        RECT 32.225 133.825 32.515 133.870 ;
        RECT 32.670 133.810 32.990 133.870 ;
        RECT 33.680 133.870 36.670 134.010 ;
        RECT 18.425 133.670 18.715 133.715 ;
        RECT 20.710 133.670 21.030 133.730 ;
        RECT 18.425 133.530 21.030 133.670 ;
        RECT 18.425 133.485 18.715 133.530 ;
        RECT 20.710 133.470 21.030 133.530 ;
        RECT 26.230 133.670 26.550 133.730 ;
        RECT 30.845 133.670 31.135 133.715 ;
        RECT 33.680 133.670 33.820 133.870 ;
        RECT 36.350 133.810 36.670 133.870 ;
        RECT 38.650 133.810 38.970 134.070 ;
        RECT 39.200 134.010 39.340 134.210 ;
        RECT 40.030 134.150 40.350 134.410 ;
        RECT 41.885 134.350 42.175 134.395 ;
        RECT 48.325 134.350 48.615 134.395 ;
        RECT 53.370 134.350 53.690 134.410 ;
        RECT 41.885 134.210 48.615 134.350 ;
        RECT 41.885 134.165 42.175 134.210 ;
        RECT 48.325 134.165 48.615 134.210 ;
        RECT 49.320 134.210 53.690 134.350 ;
        RECT 42.805 134.010 43.095 134.055 ;
        RECT 39.200 133.870 43.095 134.010 ;
        RECT 42.805 133.825 43.095 133.870 ;
        RECT 43.265 134.010 43.555 134.055 ;
        RECT 43.710 134.010 44.030 134.070 ;
        RECT 43.265 133.870 44.030 134.010 ;
        RECT 43.265 133.825 43.555 133.870 ;
        RECT 43.710 133.810 44.030 133.870 ;
        RECT 46.025 133.825 46.315 134.055 ;
        RECT 46.485 133.825 46.775 134.055 ;
        RECT 46.945 133.825 47.235 134.055 ;
        RECT 47.865 134.010 48.155 134.055 ;
        RECT 48.770 134.010 49.090 134.070 ;
        RECT 47.865 133.870 49.090 134.010 ;
        RECT 47.865 133.825 48.155 133.870 ;
        RECT 26.230 133.530 33.820 133.670 ;
        RECT 26.230 133.470 26.550 133.530 ;
        RECT 30.845 133.485 31.135 133.530 ;
        RECT 34.050 133.470 34.370 133.730 ;
        RECT 34.525 133.670 34.815 133.715 ;
        RECT 34.970 133.670 35.290 133.730 ;
        RECT 34.525 133.530 35.290 133.670 ;
        RECT 34.525 133.485 34.815 133.530 ;
        RECT 34.970 133.470 35.290 133.530 ;
        RECT 39.585 133.670 39.875 133.715 ;
        RECT 40.490 133.670 40.810 133.730 ;
        RECT 39.585 133.530 40.810 133.670 ;
        RECT 39.585 133.485 39.875 133.530 ;
        RECT 40.490 133.470 40.810 133.530 ;
        RECT 25.740 133.330 26.030 133.375 ;
        RECT 28.520 133.330 28.810 133.375 ;
        RECT 30.380 133.330 30.670 133.375 ;
        RECT 25.740 133.190 30.670 133.330 ;
        RECT 25.740 133.145 26.030 133.190 ;
        RECT 28.520 133.145 28.810 133.190 ;
        RECT 30.380 133.145 30.670 133.190 ;
        RECT 36.825 133.330 37.115 133.375 ;
        RECT 40.950 133.330 41.270 133.390 ;
        RECT 36.825 133.190 41.270 133.330 ;
        RECT 36.825 133.145 37.115 133.190 ;
        RECT 40.950 133.130 41.270 133.190 ;
        RECT 30.830 132.990 31.150 133.050 ;
        RECT 37.745 132.990 38.035 133.035 ;
        RECT 30.830 132.850 38.035 132.990 ;
        RECT 30.830 132.790 31.150 132.850 ;
        RECT 37.745 132.805 38.035 132.850 ;
        RECT 39.110 132.790 39.430 133.050 ;
        RECT 43.250 132.790 43.570 133.050 ;
        RECT 44.185 132.990 44.475 133.035 ;
        RECT 44.630 132.990 44.950 133.050 ;
        RECT 44.185 132.850 44.950 132.990 ;
        RECT 46.100 132.990 46.240 133.825 ;
        RECT 46.560 133.330 46.700 133.825 ;
        RECT 47.020 133.670 47.160 133.825 ;
        RECT 48.770 133.810 49.090 133.870 ;
        RECT 49.320 133.670 49.460 134.210 ;
        RECT 53.370 134.150 53.690 134.210 ;
        RECT 54.240 134.350 54.530 134.395 ;
        RECT 55.670 134.350 55.990 134.410 ;
        RECT 57.500 134.350 57.790 134.395 ;
        RECT 54.240 134.210 57.790 134.350 ;
        RECT 54.240 134.165 54.530 134.210 ;
        RECT 55.670 134.150 55.990 134.210 ;
        RECT 57.500 134.165 57.790 134.210 ;
        RECT 58.420 134.350 58.710 134.395 ;
        RECT 60.280 134.350 60.570 134.395 ;
        RECT 65.420 134.350 65.560 134.490 ;
        RECT 58.420 134.210 60.570 134.350 ;
        RECT 58.420 134.165 58.710 134.210 ;
        RECT 60.280 134.165 60.570 134.210 ;
        RECT 64.960 134.210 65.560 134.350 ;
        RECT 65.880 134.350 66.020 134.490 ;
        RECT 65.880 134.210 66.940 134.350 ;
        RECT 49.690 133.810 50.010 134.070 ;
        RECT 50.165 133.825 50.455 134.055 ;
        RECT 50.625 133.825 50.915 134.055 ;
        RECT 51.545 134.010 51.835 134.055 ;
        RECT 55.210 134.010 55.530 134.070 ;
        RECT 51.545 133.870 55.530 134.010 ;
        RECT 51.545 133.825 51.835 133.870 ;
        RECT 47.020 133.530 49.460 133.670 ;
        RECT 50.240 133.330 50.380 133.825 ;
        RECT 50.700 133.670 50.840 133.825 ;
        RECT 55.210 133.810 55.530 133.870 ;
        RECT 56.100 134.010 56.390 134.055 ;
        RECT 58.420 134.010 58.635 134.165 ;
        RECT 64.960 134.055 65.100 134.210 ;
        RECT 56.100 133.870 58.635 134.010 ;
        RECT 56.100 133.825 56.390 133.870 ;
        RECT 64.885 133.825 65.175 134.055 ;
        RECT 65.330 133.810 65.650 134.070 ;
        RECT 65.790 133.810 66.110 134.070 ;
        RECT 66.800 134.055 66.940 134.210 ;
        RECT 79.130 134.150 79.450 134.410 ;
        RECT 90.630 134.350 90.950 134.410 ;
        RECT 91.500 134.350 91.790 134.395 ;
        RECT 94.760 134.350 95.050 134.395 ;
        RECT 90.630 134.210 95.050 134.350 ;
        RECT 90.630 134.150 90.950 134.210 ;
        RECT 91.500 134.165 91.790 134.210 ;
        RECT 94.760 134.165 95.050 134.210 ;
        RECT 95.680 134.350 95.970 134.395 ;
        RECT 97.540 134.350 97.830 134.395 ;
        RECT 95.680 134.210 97.830 134.350 ;
        RECT 95.680 134.165 95.970 134.210 ;
        RECT 97.540 134.165 97.830 134.210 ;
        RECT 101.160 134.350 101.450 134.395 ;
        RECT 101.670 134.350 101.990 134.410 ;
        RECT 104.420 134.350 104.710 134.395 ;
        RECT 101.160 134.210 104.710 134.350 ;
        RECT 101.160 134.165 101.450 134.210 ;
        RECT 66.725 133.825 67.015 134.055 ;
        RECT 80.525 134.010 80.815 134.055 ;
        RECT 82.810 134.010 83.130 134.070 ;
        RECT 80.525 133.870 83.130 134.010 ;
        RECT 80.525 133.825 80.815 133.870 ;
        RECT 82.810 133.810 83.130 133.870 ;
        RECT 87.870 134.010 88.190 134.070 ;
        RECT 88.345 134.010 88.635 134.055 ;
        RECT 92.010 134.010 92.330 134.070 ;
        RECT 87.870 133.870 92.330 134.010 ;
        RECT 87.870 133.810 88.190 133.870 ;
        RECT 88.345 133.825 88.635 133.870 ;
        RECT 92.010 133.810 92.330 133.870 ;
        RECT 93.360 134.010 93.650 134.055 ;
        RECT 95.680 134.010 95.895 134.165 ;
        RECT 101.670 134.150 101.990 134.210 ;
        RECT 104.420 134.165 104.710 134.210 ;
        RECT 105.340 134.350 105.630 134.395 ;
        RECT 107.200 134.350 107.490 134.395 ;
        RECT 105.340 134.210 107.490 134.350 ;
        RECT 105.340 134.165 105.630 134.210 ;
        RECT 107.200 134.165 107.490 134.210 ;
        RECT 108.585 134.350 108.875 134.395 ;
        RECT 112.250 134.350 112.570 134.410 ;
        RECT 108.585 134.210 112.570 134.350 ;
        RECT 108.585 134.165 108.875 134.210 ;
        RECT 93.360 133.870 95.895 134.010 ;
        RECT 93.360 133.825 93.650 133.870 ;
        RECT 96.610 133.810 96.930 134.070 ;
        RECT 103.020 134.010 103.310 134.055 ;
        RECT 105.340 134.010 105.555 134.165 ;
        RECT 112.250 134.150 112.570 134.210 ;
        RECT 103.020 133.870 105.555 134.010 ;
        RECT 103.020 133.825 103.310 133.870 ;
        RECT 106.270 133.810 106.590 134.070 ;
        RECT 109.490 133.810 109.810 134.070 ;
        RECT 109.965 134.010 110.255 134.055 ;
        RECT 110.410 134.010 110.730 134.070 ;
        RECT 109.965 133.870 110.730 134.010 ;
        RECT 109.965 133.825 110.255 133.870 ;
        RECT 110.410 133.810 110.730 133.870 ;
        RECT 113.170 134.010 113.490 134.070 ;
        RECT 119.165 134.010 119.455 134.055 ;
        RECT 113.170 133.870 119.455 134.010 ;
        RECT 113.170 133.810 113.490 133.870 ;
        RECT 119.165 133.825 119.455 133.870 ;
        RECT 59.365 133.670 59.655 133.715 ;
        RECT 60.270 133.670 60.590 133.730 ;
        RECT 50.700 133.530 51.730 133.670 ;
        RECT 51.070 133.330 51.390 133.390 ;
        RECT 46.560 133.190 51.390 133.330 ;
        RECT 51.070 133.130 51.390 133.190 ;
        RECT 49.690 132.990 50.010 133.050 ;
        RECT 46.100 132.850 50.010 132.990 ;
        RECT 51.590 132.990 51.730 133.530 ;
        RECT 59.365 133.530 60.590 133.670 ;
        RECT 59.365 133.485 59.655 133.530 ;
        RECT 60.270 133.470 60.590 133.530 ;
        RECT 61.205 133.670 61.495 133.715 ;
        RECT 68.550 133.670 68.870 133.730 ;
        RECT 61.205 133.530 68.870 133.670 ;
        RECT 61.205 133.485 61.495 133.530 ;
        RECT 68.550 133.470 68.870 133.530 ;
        RECT 80.065 133.670 80.355 133.715 ;
        RECT 82.350 133.670 82.670 133.730 ;
        RECT 80.065 133.530 82.670 133.670 ;
        RECT 80.065 133.485 80.355 133.530 ;
        RECT 82.350 133.470 82.670 133.530 ;
        RECT 93.850 133.670 94.170 133.730 ;
        RECT 98.465 133.670 98.755 133.715 ;
        RECT 98.910 133.670 99.230 133.730 ;
        RECT 93.850 133.530 99.230 133.670 ;
        RECT 93.850 133.470 94.170 133.530 ;
        RECT 98.465 133.485 98.755 133.530 ;
        RECT 98.910 133.470 99.230 133.530 ;
        RECT 105.350 133.670 105.670 133.730 ;
        RECT 108.125 133.670 108.415 133.715 ;
        RECT 111.790 133.670 112.110 133.730 ;
        RECT 105.350 133.530 112.110 133.670 ;
        RECT 105.350 133.470 105.670 133.530 ;
        RECT 108.125 133.485 108.415 133.530 ;
        RECT 111.790 133.470 112.110 133.530 ;
        RECT 56.100 133.330 56.390 133.375 ;
        RECT 58.880 133.330 59.170 133.375 ;
        RECT 60.740 133.330 61.030 133.375 ;
        RECT 83.270 133.330 83.590 133.390 ;
        RECT 56.100 133.190 61.030 133.330 ;
        RECT 56.100 133.145 56.390 133.190 ;
        RECT 58.880 133.145 59.170 133.190 ;
        RECT 60.740 133.145 61.030 133.190 ;
        RECT 80.600 133.190 83.590 133.330 ;
        RECT 52.235 132.990 52.525 133.035 ;
        RECT 54.290 132.990 54.610 133.050 ;
        RECT 56.590 132.990 56.910 133.050 ;
        RECT 80.600 133.035 80.740 133.190 ;
        RECT 83.270 133.130 83.590 133.190 ;
        RECT 93.360 133.330 93.650 133.375 ;
        RECT 96.140 133.330 96.430 133.375 ;
        RECT 98.000 133.330 98.290 133.375 ;
        RECT 93.360 133.190 98.290 133.330 ;
        RECT 93.360 133.145 93.650 133.190 ;
        RECT 96.140 133.145 96.430 133.190 ;
        RECT 98.000 133.145 98.290 133.190 ;
        RECT 103.020 133.330 103.310 133.375 ;
        RECT 105.800 133.330 106.090 133.375 ;
        RECT 107.660 133.330 107.950 133.375 ;
        RECT 103.020 133.190 107.950 133.330 ;
        RECT 103.020 133.145 103.310 133.190 ;
        RECT 105.800 133.145 106.090 133.190 ;
        RECT 107.660 133.145 107.950 133.190 ;
        RECT 51.590 132.850 56.910 132.990 ;
        RECT 44.185 132.805 44.475 132.850 ;
        RECT 44.630 132.790 44.950 132.850 ;
        RECT 49.690 132.790 50.010 132.850 ;
        RECT 52.235 132.805 52.525 132.850 ;
        RECT 54.290 132.790 54.610 132.850 ;
        RECT 56.590 132.790 56.910 132.850 ;
        RECT 80.525 132.805 80.815 133.035 ;
        RECT 81.430 132.790 81.750 133.050 ;
        RECT 98.450 132.990 98.770 133.050 ;
        RECT 99.155 132.990 99.445 133.035 ;
        RECT 98.450 132.850 99.445 132.990 ;
        RECT 98.450 132.790 98.770 132.850 ;
        RECT 99.155 132.805 99.445 132.850 ;
        RECT 109.030 132.790 109.350 133.050 ;
        RECT 110.870 132.790 111.190 133.050 ;
        RECT 30.370 132.015 30.690 132.030 ;
        RECT 30.370 131.785 30.905 132.015 ;
        RECT 41.410 131.970 41.730 132.030 ;
        RECT 34.140 131.830 40.720 131.970 ;
        RECT 30.370 131.770 30.690 131.785 ;
        RECT 20.710 131.090 21.030 131.350 ;
        RECT 34.140 131.290 34.280 131.830 ;
        RECT 34.480 131.630 34.770 131.675 ;
        RECT 37.260 131.630 37.550 131.675 ;
        RECT 39.120 131.630 39.410 131.675 ;
        RECT 34.480 131.490 39.410 131.630 ;
        RECT 34.480 131.445 34.770 131.490 ;
        RECT 37.260 131.445 37.550 131.490 ;
        RECT 39.120 131.445 39.410 131.490 ;
        RECT 40.045 131.445 40.335 131.675 ;
        RECT 40.580 131.630 40.720 131.830 ;
        RECT 41.410 131.830 45.780 131.970 ;
        RECT 41.410 131.770 41.730 131.830 ;
        RECT 45.640 131.630 45.780 131.830 ;
        RECT 46.930 131.770 47.250 132.030 ;
        RECT 78.670 131.770 78.990 132.030 ;
        RECT 88.345 131.970 88.635 132.015 ;
        RECT 90.630 131.970 90.950 132.030 ;
        RECT 88.345 131.830 90.950 131.970 ;
        RECT 88.345 131.785 88.635 131.830 ;
        RECT 90.630 131.770 90.950 131.830 ;
        RECT 96.165 131.970 96.455 132.015 ;
        RECT 96.610 131.970 96.930 132.030 ;
        RECT 96.165 131.830 96.930 131.970 ;
        RECT 96.165 131.785 96.455 131.830 ;
        RECT 96.610 131.770 96.930 131.830 ;
        RECT 100.290 131.770 100.610 132.030 ;
        RECT 104.430 131.770 104.750 132.030 ;
        RECT 109.950 131.970 110.270 132.030 ;
        RECT 110.425 131.970 110.715 132.015 ;
        RECT 109.950 131.830 110.715 131.970 ;
        RECT 109.950 131.770 110.270 131.830 ;
        RECT 110.425 131.785 110.715 131.830 ;
        RECT 69.945 131.630 70.235 131.675 ;
        RECT 99.370 131.630 99.690 131.690 ;
        RECT 40.580 131.490 45.320 131.630 ;
        RECT 45.640 131.490 99.690 131.630 ;
        RECT 21.720 131.150 34.280 131.290 ;
        RECT 36.810 131.290 37.130 131.350 ;
        RECT 37.745 131.290 38.035 131.335 ;
        RECT 40.120 131.290 40.260 131.445 ;
        RECT 45.180 131.335 45.320 131.490 ;
        RECT 69.945 131.445 70.235 131.490 ;
        RECT 99.370 131.430 99.690 131.490 ;
        RECT 36.810 131.150 37.500 131.290 ;
        RECT 19.330 130.950 19.650 131.010 ;
        RECT 21.720 130.995 21.860 131.150 ;
        RECT 36.810 131.090 37.130 131.150 ;
        RECT 21.645 130.950 21.935 130.995 ;
        RECT 19.330 130.810 21.935 130.950 ;
        RECT 19.330 130.750 19.650 130.810 ;
        RECT 21.645 130.765 21.935 130.810 ;
        RECT 34.480 130.950 34.770 130.995 ;
        RECT 37.360 130.950 37.500 131.150 ;
        RECT 37.745 131.150 40.260 131.290 ;
        RECT 37.745 131.105 38.035 131.150 ;
        RECT 45.105 131.105 45.395 131.335 ;
        RECT 66.265 131.290 66.555 131.335 ;
        RECT 69.010 131.290 69.330 131.350 ;
        RECT 66.265 131.150 69.330 131.290 ;
        RECT 66.265 131.105 66.555 131.150 ;
        RECT 69.010 131.090 69.330 131.150 ;
        RECT 73.625 131.290 73.915 131.335 ;
        RECT 74.070 131.290 74.390 131.350 ;
        RECT 73.625 131.150 74.390 131.290 ;
        RECT 73.625 131.105 73.915 131.150 ;
        RECT 74.070 131.090 74.390 131.150 ;
        RECT 79.130 131.290 79.450 131.350 ;
        RECT 89.725 131.290 90.015 131.335 ;
        RECT 79.130 131.150 90.015 131.290 ;
        RECT 79.130 131.090 79.450 131.150 ;
        RECT 89.725 131.105 90.015 131.150 ;
        RECT 99.830 131.090 100.150 131.350 ;
        RECT 103.050 131.290 103.370 131.350 ;
        RECT 104.445 131.290 104.735 131.335 ;
        RECT 103.050 131.150 104.735 131.290 ;
        RECT 103.050 131.090 103.370 131.150 ;
        RECT 104.445 131.105 104.735 131.150 ;
        RECT 39.585 130.950 39.875 130.995 ;
        RECT 40.490 130.950 40.810 131.010 ;
        RECT 34.480 130.810 37.015 130.950 ;
        RECT 37.360 130.810 40.810 130.950 ;
        RECT 34.480 130.765 34.770 130.810 ;
        RECT 22.105 130.610 22.395 130.655 ;
        RECT 24.390 130.610 24.710 130.670 ;
        RECT 32.620 130.610 32.910 130.655 ;
        RECT 34.050 130.610 34.370 130.670 ;
        RECT 36.800 130.655 37.015 130.810 ;
        RECT 39.585 130.765 39.875 130.810 ;
        RECT 40.490 130.750 40.810 130.810 ;
        RECT 40.950 130.750 41.270 131.010 ;
        RECT 42.805 130.765 43.095 130.995 ;
        RECT 43.725 130.950 44.015 130.995 ;
        RECT 46.025 130.950 46.315 130.995 ;
        RECT 46.930 130.950 47.250 131.010 ;
        RECT 43.725 130.810 47.250 130.950 ;
        RECT 43.725 130.765 44.015 130.810 ;
        RECT 46.025 130.765 46.315 130.810 ;
        RECT 35.880 130.610 36.170 130.655 ;
        RECT 22.105 130.470 27.840 130.610 ;
        RECT 22.105 130.425 22.395 130.470 ;
        RECT 24.390 130.410 24.710 130.470 ;
        RECT 27.700 130.330 27.840 130.470 ;
        RECT 32.620 130.470 36.170 130.610 ;
        RECT 32.620 130.425 32.910 130.470 ;
        RECT 34.050 130.410 34.370 130.470 ;
        RECT 35.880 130.425 36.170 130.470 ;
        RECT 36.800 130.610 37.090 130.655 ;
        RECT 38.660 130.610 38.950 130.655 ;
        RECT 36.800 130.470 38.950 130.610 ;
        RECT 36.800 130.425 37.090 130.470 ;
        RECT 38.660 130.425 38.950 130.470 ;
        RECT 23.010 130.270 23.330 130.330 ;
        RECT 23.945 130.270 24.235 130.315 ;
        RECT 23.010 130.130 24.235 130.270 ;
        RECT 23.010 130.070 23.330 130.130 ;
        RECT 23.945 130.085 24.235 130.130 ;
        RECT 27.610 130.270 27.930 130.330 ;
        RECT 42.880 130.270 43.020 130.765 ;
        RECT 46.930 130.750 47.250 130.810 ;
        RECT 70.865 130.950 71.155 130.995 ;
        RECT 72.690 130.950 73.010 131.010 ;
        RECT 74.545 130.950 74.835 130.995 ;
        RECT 79.605 130.950 79.895 130.995 ;
        RECT 70.865 130.810 74.835 130.950 ;
        RECT 70.865 130.765 71.155 130.810 ;
        RECT 72.690 130.750 73.010 130.810 ;
        RECT 74.545 130.765 74.835 130.810 ;
        RECT 75.080 130.810 79.895 130.950 ;
        RECT 44.645 130.610 44.935 130.655 ;
        RECT 48.310 130.610 48.630 130.670 ;
        RECT 44.645 130.470 48.630 130.610 ;
        RECT 44.645 130.425 44.935 130.470 ;
        RECT 48.310 130.410 48.630 130.470 ;
        RECT 64.870 130.610 65.190 130.670 ;
        RECT 65.790 130.610 66.110 130.670 ;
        RECT 67.185 130.610 67.475 130.655 ;
        RECT 64.870 130.470 67.475 130.610 ;
        RECT 64.870 130.410 65.190 130.470 ;
        RECT 65.790 130.410 66.110 130.470 ;
        RECT 67.185 130.425 67.475 130.470 ;
        RECT 75.080 130.330 75.220 130.810 ;
        RECT 79.605 130.765 79.895 130.810 ;
        RECT 80.065 130.765 80.355 130.995 ;
        RECT 78.670 130.610 78.990 130.670 ;
        RECT 80.140 130.610 80.280 130.765 ;
        RECT 87.870 130.750 88.190 131.010 ;
        RECT 93.865 130.950 94.155 130.995 ;
        RECT 93.020 130.810 94.155 130.950 ;
        RECT 78.670 130.470 80.280 130.610 ;
        RECT 78.670 130.410 78.990 130.470 ;
        RECT 27.610 130.130 43.020 130.270 ;
        RECT 66.250 130.270 66.570 130.330 ;
        RECT 66.725 130.270 67.015 130.315 ;
        RECT 66.250 130.130 67.015 130.270 ;
        RECT 27.610 130.070 27.930 130.130 ;
        RECT 66.250 130.070 66.570 130.130 ;
        RECT 66.725 130.085 67.015 130.130 ;
        RECT 69.025 130.270 69.315 130.315 ;
        RECT 69.930 130.270 70.250 130.330 ;
        RECT 69.025 130.130 70.250 130.270 ;
        RECT 69.025 130.085 69.315 130.130 ;
        RECT 69.930 130.070 70.250 130.130 ;
        RECT 71.785 130.270 72.075 130.315 ;
        RECT 73.150 130.270 73.470 130.330 ;
        RECT 71.785 130.130 73.470 130.270 ;
        RECT 71.785 130.085 72.075 130.130 ;
        RECT 73.150 130.070 73.470 130.130 ;
        RECT 74.990 130.070 75.310 130.330 ;
        RECT 80.970 130.270 81.290 130.330 ;
        RECT 90.645 130.270 90.935 130.315 ;
        RECT 80.970 130.130 90.935 130.270 ;
        RECT 80.970 130.070 81.290 130.130 ;
        RECT 90.645 130.085 90.935 130.130 ;
        RECT 91.105 130.270 91.395 130.315 ;
        RECT 91.550 130.270 91.870 130.330 ;
        RECT 93.020 130.315 93.160 130.810 ;
        RECT 93.865 130.765 94.155 130.810 ;
        RECT 95.230 130.750 95.550 131.010 ;
        RECT 97.530 130.950 97.850 131.010 ;
        RECT 98.925 130.950 99.215 130.995 ;
        RECT 97.530 130.810 99.215 130.950 ;
        RECT 97.530 130.750 97.850 130.810 ;
        RECT 98.925 130.765 99.215 130.810 ;
        RECT 100.305 130.950 100.595 130.995 ;
        RECT 101.210 130.950 101.530 131.010 ;
        RECT 100.305 130.810 101.530 130.950 ;
        RECT 100.305 130.765 100.595 130.810 ;
        RECT 101.210 130.750 101.530 130.810 ;
        RECT 104.890 130.950 105.210 131.010 ;
        RECT 105.365 130.950 105.655 130.995 ;
        RECT 104.890 130.810 105.655 130.950 ;
        RECT 104.890 130.750 105.210 130.810 ;
        RECT 105.365 130.765 105.655 130.810 ;
        RECT 109.950 130.950 110.270 131.010 ;
        RECT 111.345 130.950 111.635 130.995 ;
        RECT 109.950 130.810 111.635 130.950 ;
        RECT 109.950 130.750 110.270 130.810 ;
        RECT 111.345 130.765 111.635 130.810 ;
        RECT 112.250 130.750 112.570 131.010 ;
        RECT 103.985 130.610 104.275 130.655 ;
        RECT 105.810 130.610 106.130 130.670 ;
        RECT 103.985 130.470 106.130 130.610 ;
        RECT 103.985 130.425 104.275 130.470 ;
        RECT 105.810 130.410 106.130 130.470 ;
        RECT 91.105 130.130 91.870 130.270 ;
        RECT 91.105 130.085 91.395 130.130 ;
        RECT 91.550 130.070 91.870 130.130 ;
        RECT 92.945 130.085 93.235 130.315 ;
        RECT 94.785 130.270 95.075 130.315 ;
        RECT 97.070 130.270 97.390 130.330 ;
        RECT 94.785 130.130 97.390 130.270 ;
        RECT 94.785 130.085 95.075 130.130 ;
        RECT 97.070 130.070 97.390 130.130 ;
        RECT 97.990 130.070 98.310 130.330 ;
        RECT 106.285 130.270 106.575 130.315 ;
        RECT 107.190 130.270 107.510 130.330 ;
        RECT 106.285 130.130 107.510 130.270 ;
        RECT 106.285 130.085 106.575 130.130 ;
        RECT 107.190 130.070 107.510 130.130 ;
        RECT 17.275 129.250 17.565 129.295 ;
        RECT 24.390 129.250 24.710 129.310 ;
        RECT 17.275 129.110 24.710 129.250 ;
        RECT 17.275 129.065 17.565 129.110 ;
        RECT 24.390 129.050 24.710 129.110 ;
        RECT 34.050 129.050 34.370 129.310 ;
        RECT 36.825 129.250 37.115 129.295 ;
        RECT 37.270 129.250 37.590 129.310 ;
        RECT 36.825 129.110 37.590 129.250 ;
        RECT 36.825 129.065 37.115 129.110 ;
        RECT 37.270 129.050 37.590 129.110 ;
        RECT 47.390 129.250 47.710 129.310 ;
        RECT 48.325 129.250 48.615 129.295 ;
        RECT 47.390 129.110 48.615 129.250 ;
        RECT 47.390 129.050 47.710 129.110 ;
        RECT 48.325 129.065 48.615 129.110 ;
        RECT 53.370 129.250 53.690 129.310 ;
        RECT 56.130 129.250 56.450 129.310 ;
        RECT 53.370 129.110 56.450 129.250 ;
        RECT 53.370 129.050 53.690 129.110 ;
        RECT 56.130 129.050 56.450 129.110 ;
        RECT 56.590 129.050 56.910 129.310 ;
        RECT 58.445 129.065 58.735 129.295 ;
        RECT 65.115 129.250 65.405 129.295 ;
        RECT 66.250 129.250 66.570 129.310 ;
        RECT 74.990 129.250 75.310 129.310 ;
        RECT 65.115 129.110 66.570 129.250 ;
        RECT 65.115 129.065 65.405 129.110 ;
        RECT 19.280 128.910 19.570 128.955 ;
        RECT 20.710 128.910 21.030 128.970 ;
        RECT 22.540 128.910 22.830 128.955 ;
        RECT 19.280 128.770 22.830 128.910 ;
        RECT 19.280 128.725 19.570 128.770 ;
        RECT 20.710 128.710 21.030 128.770 ;
        RECT 22.540 128.725 22.830 128.770 ;
        RECT 23.460 128.910 23.750 128.955 ;
        RECT 25.320 128.910 25.610 128.955 ;
        RECT 23.460 128.770 25.610 128.910 ;
        RECT 23.460 128.725 23.750 128.770 ;
        RECT 25.320 128.725 25.610 128.770 ;
        RECT 21.140 128.570 21.430 128.615 ;
        RECT 23.460 128.570 23.675 128.725 ;
        RECT 21.140 128.430 23.675 128.570 ;
        RECT 21.140 128.385 21.430 128.430 ;
        RECT 26.230 128.370 26.550 128.630 ;
        RECT 31.290 128.570 31.610 128.630 ;
        RECT 33.605 128.570 33.895 128.615 ;
        RECT 31.290 128.430 33.895 128.570 ;
        RECT 31.290 128.370 31.610 128.430 ;
        RECT 33.605 128.385 33.895 128.430 ;
        RECT 35.905 128.570 36.195 128.615 ;
        RECT 38.190 128.570 38.510 128.630 ;
        RECT 41.410 128.570 41.730 128.630 ;
        RECT 35.905 128.430 41.730 128.570 ;
        RECT 35.905 128.385 36.195 128.430 ;
        RECT 38.190 128.370 38.510 128.430 ;
        RECT 41.410 128.370 41.730 128.430 ;
        RECT 46.930 128.570 47.250 128.630 ;
        RECT 47.405 128.570 47.695 128.615 ;
        RECT 58.520 128.570 58.660 129.065 ;
        RECT 66.250 129.050 66.570 129.110 ;
        RECT 66.800 129.110 75.310 129.250 ;
        RECT 58.905 128.570 59.195 128.615 ;
        RECT 46.930 128.430 56.360 128.570 ;
        RECT 58.520 128.430 59.195 128.570 ;
        RECT 46.930 128.370 47.250 128.430 ;
        RECT 47.405 128.385 47.695 128.430 ;
        RECT 24.390 128.030 24.710 128.290 ;
        RECT 34.970 128.030 35.290 128.290 ;
        RECT 46.485 128.045 46.775 128.275 ;
        RECT 54.750 128.230 55.070 128.290 ;
        RECT 55.225 128.230 55.515 128.275 ;
        RECT 54.750 128.090 55.515 128.230 ;
        RECT 56.220 128.230 56.360 128.430 ;
        RECT 58.905 128.385 59.195 128.430 ;
        RECT 66.800 128.230 66.940 129.110 ;
        RECT 74.990 129.050 75.310 129.110 ;
        RECT 76.370 129.050 76.690 129.310 ;
        RECT 78.685 129.250 78.975 129.295 ;
        RECT 80.050 129.250 80.370 129.310 ;
        RECT 78.685 129.110 80.370 129.250 ;
        RECT 78.685 129.065 78.975 129.110 ;
        RECT 80.050 129.050 80.370 129.110 ;
        RECT 80.970 129.050 81.290 129.310 ;
        RECT 83.270 129.050 83.590 129.310 ;
        RECT 100.290 129.250 100.610 129.310 ;
        RECT 101.225 129.250 101.515 129.295 ;
        RECT 100.290 129.110 101.515 129.250 ;
        RECT 100.290 129.050 100.610 129.110 ;
        RECT 101.225 129.065 101.515 129.110 ;
        RECT 104.430 129.050 104.750 129.310 ;
        RECT 106.730 129.050 107.050 129.310 ;
        RECT 109.030 129.050 109.350 129.310 ;
        RECT 114.090 129.250 114.410 129.310 ;
        RECT 115.025 129.250 115.315 129.295 ;
        RECT 114.090 129.110 115.315 129.250 ;
        RECT 114.090 129.050 114.410 129.110 ;
        RECT 115.025 129.065 115.315 129.110 ;
        RECT 67.120 128.910 67.410 128.955 ;
        RECT 69.470 128.910 69.790 128.970 ;
        RECT 70.380 128.910 70.670 128.955 ;
        RECT 67.120 128.770 70.670 128.910 ;
        RECT 67.120 128.725 67.410 128.770 ;
        RECT 69.470 128.710 69.790 128.770 ;
        RECT 70.380 128.725 70.670 128.770 ;
        RECT 71.300 128.910 71.590 128.955 ;
        RECT 73.160 128.910 73.450 128.955 ;
        RECT 71.300 128.770 73.450 128.910 ;
        RECT 71.300 128.725 71.590 128.770 ;
        RECT 73.160 128.725 73.450 128.770 ;
        RECT 76.830 128.910 77.150 128.970 ;
        RECT 81.060 128.910 81.200 129.050 ;
        RECT 76.830 128.770 81.200 128.910 ;
        RECT 91.090 128.910 91.410 128.970 ;
        RECT 91.960 128.910 92.250 128.955 ;
        RECT 95.220 128.910 95.510 128.955 ;
        RECT 91.090 128.770 95.510 128.910 ;
        RECT 68.980 128.570 69.270 128.615 ;
        RECT 71.300 128.570 71.515 128.725 ;
        RECT 76.830 128.710 77.150 128.770 ;
        RECT 91.090 128.710 91.410 128.770 ;
        RECT 91.960 128.725 92.250 128.770 ;
        RECT 95.220 128.725 95.510 128.770 ;
        RECT 96.140 128.910 96.430 128.955 ;
        RECT 98.000 128.910 98.290 128.955 ;
        RECT 96.140 128.770 98.290 128.910 ;
        RECT 96.140 128.725 96.430 128.770 ;
        RECT 98.000 128.725 98.290 128.770 ;
        RECT 68.980 128.430 71.515 128.570 ;
        RECT 71.770 128.570 72.090 128.630 ;
        RECT 72.245 128.570 72.535 128.615 ;
        RECT 71.770 128.430 72.535 128.570 ;
        RECT 68.980 128.385 69.270 128.430 ;
        RECT 71.770 128.370 72.090 128.430 ;
        RECT 72.245 128.385 72.535 128.430 ;
        RECT 74.990 128.570 75.310 128.630 ;
        RECT 75.465 128.570 75.755 128.615 ;
        RECT 77.765 128.570 78.055 128.615 ;
        RECT 74.990 128.430 78.055 128.570 ;
        RECT 74.990 128.370 75.310 128.430 ;
        RECT 75.465 128.385 75.755 128.430 ;
        RECT 77.765 128.385 78.055 128.430 ;
        RECT 78.210 128.570 78.530 128.630 ;
        RECT 80.525 128.570 80.815 128.615 ;
        RECT 78.210 128.430 80.815 128.570 ;
        RECT 56.220 128.090 66.940 128.230 ;
        RECT 68.550 128.230 68.870 128.290 ;
        RECT 74.085 128.230 74.375 128.275 ;
        RECT 68.550 128.090 74.375 128.230 ;
        RECT 21.140 127.890 21.430 127.935 ;
        RECT 23.920 127.890 24.210 127.935 ;
        RECT 25.780 127.890 26.070 127.935 ;
        RECT 21.140 127.750 26.070 127.890 ;
        RECT 21.140 127.705 21.430 127.750 ;
        RECT 23.920 127.705 24.210 127.750 ;
        RECT 25.780 127.705 26.070 127.750 ;
        RECT 28.070 127.890 28.390 127.950 ;
        RECT 46.560 127.890 46.700 128.045 ;
        RECT 54.750 128.030 55.070 128.090 ;
        RECT 55.225 128.045 55.515 128.090 ;
        RECT 68.550 128.030 68.870 128.090 ;
        RECT 74.085 128.045 74.375 128.090 ;
        RECT 74.545 128.230 74.835 128.275 ;
        RECT 74.545 128.090 76.600 128.230 ;
        RECT 74.545 128.045 74.835 128.090 ;
        RECT 28.070 127.750 46.700 127.890 ;
        RECT 68.980 127.890 69.270 127.935 ;
        RECT 71.760 127.890 72.050 127.935 ;
        RECT 73.620 127.890 73.910 127.935 ;
        RECT 68.980 127.750 73.910 127.890 ;
        RECT 28.070 127.690 28.390 127.750 ;
        RECT 68.980 127.705 69.270 127.750 ;
        RECT 71.760 127.705 72.050 127.750 ;
        RECT 73.620 127.705 73.910 127.750 ;
        RECT 59.825 127.550 60.115 127.595 ;
        RECT 60.270 127.550 60.590 127.610 ;
        RECT 59.825 127.410 60.590 127.550 ;
        RECT 76.460 127.550 76.600 128.090 ;
        RECT 76.830 128.030 77.150 128.290 ;
        RECT 77.840 128.230 77.980 128.385 ;
        RECT 78.210 128.370 78.530 128.430 ;
        RECT 80.525 128.385 80.815 128.430 ;
        RECT 84.205 128.385 84.495 128.615 ;
        RECT 93.820 128.570 94.110 128.615 ;
        RECT 96.140 128.570 96.355 128.725 ;
        RECT 99.370 128.710 99.690 128.970 ;
        RECT 111.790 128.910 112.110 128.970 ;
        RECT 113.645 128.910 113.935 128.955 ;
        RECT 111.790 128.770 113.935 128.910 ;
        RECT 111.790 128.710 112.110 128.770 ;
        RECT 113.645 128.725 113.935 128.770 ;
        RECT 93.820 128.430 96.355 128.570 ;
        RECT 93.820 128.385 94.110 128.430 ;
        RECT 77.840 128.090 78.440 128.230 ;
        RECT 78.300 127.890 78.440 128.090 ;
        RECT 79.590 128.030 79.910 128.290 ;
        RECT 84.280 127.890 84.420 128.385 ;
        RECT 97.070 128.370 97.390 128.630 ;
        RECT 98.910 128.370 99.230 128.630 ;
        RECT 99.460 128.570 99.600 128.710 ;
        RECT 100.305 128.570 100.595 128.615 ;
        RECT 105.365 128.570 105.655 128.615 ;
        RECT 107.665 128.570 107.955 128.615 ;
        RECT 109.950 128.570 110.270 128.630 ;
        RECT 99.460 128.430 110.270 128.570 ;
        RECT 100.305 128.385 100.595 128.430 ;
        RECT 105.365 128.385 105.655 128.430 ;
        RECT 107.665 128.385 107.955 128.430 ;
        RECT 109.950 128.370 110.270 128.430 ;
        RECT 110.410 128.370 110.730 128.630 ;
        RECT 115.945 128.570 116.235 128.615 ;
        RECT 110.960 128.430 116.235 128.570 ;
        RECT 85.110 128.030 85.430 128.290 ;
        RECT 97.530 128.230 97.850 128.290 ;
        RECT 99.385 128.230 99.675 128.275 ;
        RECT 97.530 128.090 99.675 128.230 ;
        RECT 97.530 128.030 97.850 128.090 ;
        RECT 99.385 128.045 99.675 128.090 ;
        RECT 104.890 128.230 105.210 128.290 ;
        RECT 106.285 128.230 106.575 128.275 ;
        RECT 104.890 128.090 106.575 128.230 ;
        RECT 104.890 128.030 105.210 128.090 ;
        RECT 106.285 128.045 106.575 128.090 ;
        RECT 108.585 128.230 108.875 128.275 ;
        RECT 109.030 128.230 109.350 128.290 ;
        RECT 108.585 128.090 109.350 128.230 ;
        RECT 110.040 128.230 110.180 128.370 ;
        RECT 110.960 128.230 111.100 128.430 ;
        RECT 115.945 128.385 116.235 128.430 ;
        RECT 116.390 128.370 116.710 128.630 ;
        RECT 116.850 128.570 117.170 128.630 ;
        RECT 118.245 128.570 118.535 128.615 ;
        RECT 116.850 128.430 118.535 128.570 ;
        RECT 116.850 128.370 117.170 128.430 ;
        RECT 118.245 128.385 118.535 128.430 ;
        RECT 120.085 128.385 120.375 128.615 ;
        RECT 110.040 128.090 111.100 128.230 ;
        RECT 115.010 128.230 115.330 128.290 ;
        RECT 120.160 128.230 120.300 128.385 ;
        RECT 115.010 128.090 120.300 128.230 ;
        RECT 108.585 128.045 108.875 128.090 ;
        RECT 78.300 127.750 84.420 127.890 ;
        RECT 93.820 127.890 94.110 127.935 ;
        RECT 96.600 127.890 96.890 127.935 ;
        RECT 98.460 127.890 98.750 127.935 ;
        RECT 93.820 127.750 98.750 127.890 ;
        RECT 93.820 127.705 94.110 127.750 ;
        RECT 96.600 127.705 96.890 127.750 ;
        RECT 98.460 127.705 98.750 127.750 ;
        RECT 78.210 127.550 78.530 127.610 ;
        RECT 76.460 127.410 78.530 127.550 ;
        RECT 59.825 127.365 60.115 127.410 ;
        RECT 60.270 127.350 60.590 127.410 ;
        RECT 78.210 127.350 78.530 127.410 ;
        RECT 82.825 127.550 83.115 127.595 ;
        RECT 83.270 127.550 83.590 127.610 ;
        RECT 82.825 127.410 83.590 127.550 ;
        RECT 82.825 127.365 83.115 127.410 ;
        RECT 83.270 127.350 83.590 127.410 ;
        RECT 89.955 127.550 90.245 127.595 ;
        RECT 91.550 127.550 91.870 127.610 ;
        RECT 108.660 127.550 108.800 128.045 ;
        RECT 109.030 128.030 109.350 128.090 ;
        RECT 115.010 128.030 115.330 128.090 ;
        RECT 89.955 127.410 108.800 127.550 ;
        RECT 89.955 127.365 90.245 127.410 ;
        RECT 91.550 127.350 91.870 127.410 ;
        RECT 118.690 127.350 119.010 127.610 ;
        RECT 120.990 127.350 121.310 127.610 ;
        RECT 23.945 126.530 24.235 126.575 ;
        RECT 24.390 126.530 24.710 126.590 ;
        RECT 23.945 126.390 24.710 126.530 ;
        RECT 23.945 126.345 24.235 126.390 ;
        RECT 24.390 126.330 24.710 126.390 ;
        RECT 69.025 126.530 69.315 126.575 ;
        RECT 69.470 126.530 69.790 126.590 ;
        RECT 69.025 126.390 69.790 126.530 ;
        RECT 69.025 126.345 69.315 126.390 ;
        RECT 69.470 126.330 69.790 126.390 ;
        RECT 70.850 126.330 71.170 126.590 ;
        RECT 76.830 126.575 77.150 126.590 ;
        RECT 76.615 126.345 77.150 126.575 ;
        RECT 76.830 126.330 77.150 126.345 ;
        RECT 115.010 126.330 115.330 126.590 ;
        RECT 21.170 126.190 21.490 126.250 ;
        RECT 54.750 126.190 55.070 126.250 ;
        RECT 74.545 126.190 74.835 126.235 ;
        RECT 79.590 126.190 79.910 126.250 ;
        RECT 21.170 126.050 23.010 126.190 ;
        RECT 21.170 125.990 21.490 126.050 ;
        RECT 22.870 125.850 23.010 126.050 ;
        RECT 54.750 126.050 61.420 126.190 ;
        RECT 54.750 125.990 55.070 126.050 ;
        RECT 29.465 125.850 29.755 125.895 ;
        RECT 34.065 125.850 34.355 125.895 ;
        RECT 34.510 125.850 34.830 125.910 ;
        RECT 37.730 125.850 38.050 125.910 ;
        RECT 22.870 125.710 38.050 125.850 ;
        RECT 29.465 125.665 29.755 125.710 ;
        RECT 34.065 125.665 34.355 125.710 ;
        RECT 34.510 125.650 34.830 125.710 ;
        RECT 37.730 125.650 38.050 125.710 ;
        RECT 42.790 125.650 43.110 125.910 ;
        RECT 56.130 125.850 56.450 125.910 ;
        RECT 61.280 125.895 61.420 126.050 ;
        RECT 74.545 126.050 79.910 126.190 ;
        RECT 74.545 126.005 74.835 126.050 ;
        RECT 79.590 125.990 79.910 126.050 ;
        RECT 80.480 126.190 80.770 126.235 ;
        RECT 83.260 126.190 83.550 126.235 ;
        RECT 85.120 126.190 85.410 126.235 ;
        RECT 80.480 126.050 85.410 126.190 ;
        RECT 80.480 126.005 80.770 126.050 ;
        RECT 83.260 126.005 83.550 126.050 ;
        RECT 85.120 126.005 85.410 126.050 ;
        RECT 119.580 126.190 119.870 126.235 ;
        RECT 122.360 126.190 122.650 126.235 ;
        RECT 124.220 126.190 124.510 126.235 ;
        RECT 119.580 126.050 124.510 126.190 ;
        RECT 119.580 126.005 119.870 126.050 ;
        RECT 122.360 126.005 122.650 126.050 ;
        RECT 124.220 126.005 124.510 126.050 ;
        RECT 61.205 125.850 61.495 125.895 ;
        RECT 64.410 125.850 64.730 125.910 ;
        RECT 43.800 125.710 46.240 125.850 ;
        RECT 20.710 125.510 21.030 125.570 ;
        RECT 21.185 125.510 21.475 125.555 ;
        RECT 20.710 125.370 21.475 125.510 ;
        RECT 20.710 125.310 21.030 125.370 ;
        RECT 21.185 125.325 21.475 125.370 ;
        RECT 21.630 125.310 21.950 125.570 ;
        RECT 23.010 125.310 23.330 125.570 ;
        RECT 27.150 125.510 27.470 125.570 ;
        RECT 28.070 125.510 28.390 125.570 ;
        RECT 27.150 125.370 28.390 125.510 ;
        RECT 27.150 125.310 27.470 125.370 ;
        RECT 28.070 125.310 28.390 125.370 ;
        RECT 37.285 125.325 37.575 125.555 ;
        RECT 27.610 125.170 27.930 125.230 ;
        RECT 28.545 125.170 28.835 125.215 ;
        RECT 37.360 125.170 37.500 125.325 ;
        RECT 38.190 125.310 38.510 125.570 ;
        RECT 39.110 125.310 39.430 125.570 ;
        RECT 39.570 125.510 39.890 125.570 ;
        RECT 43.800 125.555 43.940 125.710 ;
        RECT 40.505 125.510 40.795 125.555 ;
        RECT 39.570 125.370 40.795 125.510 ;
        RECT 39.570 125.310 39.890 125.370 ;
        RECT 40.505 125.325 40.795 125.370 ;
        RECT 41.425 125.510 41.715 125.555 ;
        RECT 43.725 125.510 44.015 125.555 ;
        RECT 41.425 125.370 44.015 125.510 ;
        RECT 41.425 125.325 41.715 125.370 ;
        RECT 43.725 125.325 44.015 125.370 ;
        RECT 44.645 125.510 44.935 125.555 ;
        RECT 45.550 125.510 45.870 125.570 ;
        RECT 46.100 125.555 46.240 125.710 ;
        RECT 56.130 125.710 60.960 125.850 ;
        RECT 56.130 125.650 56.450 125.710 ;
        RECT 44.645 125.370 45.870 125.510 ;
        RECT 44.645 125.325 44.935 125.370 ;
        RECT 45.550 125.310 45.870 125.370 ;
        RECT 46.025 125.510 46.315 125.555 ;
        RECT 46.470 125.510 46.790 125.570 ;
        RECT 46.025 125.370 46.790 125.510 ;
        RECT 46.025 125.325 46.315 125.370 ;
        RECT 46.470 125.310 46.790 125.370 ;
        RECT 46.945 125.510 47.235 125.555 ;
        RECT 47.850 125.510 48.170 125.570 ;
        RECT 46.945 125.370 48.170 125.510 ;
        RECT 46.945 125.325 47.235 125.370 ;
        RECT 47.850 125.310 48.170 125.370 ;
        RECT 49.245 125.510 49.535 125.555 ;
        RECT 60.820 125.510 60.960 125.710 ;
        RECT 61.205 125.710 64.730 125.850 ;
        RECT 61.205 125.665 61.495 125.710 ;
        RECT 64.410 125.650 64.730 125.710 ;
        RECT 105.810 125.850 106.130 125.910 ;
        RECT 107.665 125.850 107.955 125.895 ;
        RECT 111.805 125.850 112.095 125.895 ;
        RECT 105.810 125.710 112.095 125.850 ;
        RECT 105.810 125.650 106.130 125.710 ;
        RECT 107.665 125.665 107.955 125.710 ;
        RECT 111.805 125.665 112.095 125.710 ;
        RECT 120.990 125.850 121.310 125.910 ;
        RECT 122.845 125.850 123.135 125.895 ;
        RECT 120.990 125.710 123.135 125.850 ;
        RECT 120.990 125.650 121.310 125.710 ;
        RECT 122.845 125.665 123.135 125.710 ;
        RECT 62.125 125.510 62.415 125.555 ;
        RECT 49.245 125.370 60.500 125.510 ;
        RECT 60.820 125.370 62.415 125.510 ;
        RECT 49.245 125.325 49.535 125.370 ;
        RECT 27.610 125.030 28.835 125.170 ;
        RECT 27.610 124.970 27.930 125.030 ;
        RECT 28.545 124.985 28.835 125.030 ;
        RECT 34.600 125.030 37.500 125.170 ;
        RECT 43.250 125.170 43.570 125.230 ;
        RECT 45.105 125.170 45.395 125.215 ;
        RECT 43.250 125.030 45.395 125.170 ;
        RECT 34.600 124.890 34.740 125.030 ;
        RECT 43.250 124.970 43.570 125.030 ;
        RECT 45.105 124.985 45.395 125.030 ;
        RECT 51.070 124.970 51.390 125.230 ;
        RECT 60.360 125.170 60.500 125.370 ;
        RECT 62.125 125.325 62.415 125.370 ;
        RECT 69.485 125.325 69.775 125.555 ;
        RECT 62.570 125.170 62.890 125.230 ;
        RECT 60.360 125.030 62.890 125.170 ;
        RECT 69.560 125.170 69.700 125.325 ;
        RECT 69.930 125.310 70.250 125.570 ;
        RECT 80.480 125.510 80.770 125.555 ;
        RECT 80.480 125.370 83.015 125.510 ;
        RECT 80.480 125.325 80.770 125.370 ;
        RECT 70.390 125.170 70.710 125.230 ;
        RECT 69.560 125.030 70.710 125.170 ;
        RECT 62.570 124.970 62.890 125.030 ;
        RECT 70.390 124.970 70.710 125.030 ;
        RECT 73.150 124.970 73.470 125.230 ;
        RECT 81.890 125.215 82.210 125.230 ;
        RECT 78.620 125.170 78.910 125.215 ;
        RECT 81.880 125.170 82.210 125.215 ;
        RECT 78.620 125.030 82.210 125.170 ;
        RECT 78.620 124.985 78.910 125.030 ;
        RECT 81.880 124.985 82.210 125.030 ;
        RECT 82.800 125.215 83.015 125.370 ;
        RECT 83.730 125.310 84.050 125.570 ;
        RECT 85.585 125.510 85.875 125.555 ;
        RECT 96.625 125.510 96.915 125.555 ;
        RECT 98.450 125.510 98.770 125.570 ;
        RECT 85.585 125.370 98.770 125.510 ;
        RECT 85.585 125.325 85.875 125.370 ;
        RECT 96.625 125.325 96.915 125.370 ;
        RECT 98.450 125.310 98.770 125.370 ;
        RECT 109.030 125.510 109.350 125.570 ;
        RECT 112.725 125.510 113.015 125.555 ;
        RECT 109.030 125.370 113.015 125.510 ;
        RECT 109.030 125.310 109.350 125.370 ;
        RECT 112.725 125.325 113.015 125.370 ;
        RECT 119.580 125.510 119.870 125.555 ;
        RECT 119.580 125.370 122.115 125.510 ;
        RECT 119.580 125.325 119.870 125.370 ;
        RECT 82.800 125.170 83.090 125.215 ;
        RECT 84.660 125.170 84.950 125.215 ;
        RECT 82.800 125.030 84.950 125.170 ;
        RECT 82.800 124.985 83.090 125.030 ;
        RECT 84.660 124.985 84.950 125.030 ;
        RECT 108.585 125.170 108.875 125.215 ;
        RECT 113.185 125.170 113.475 125.215 ;
        RECT 115.715 125.170 116.005 125.215 ;
        RECT 116.390 125.170 116.710 125.230 ;
        RECT 108.585 125.030 116.710 125.170 ;
        RECT 108.585 124.985 108.875 125.030 ;
        RECT 113.185 124.985 113.475 125.030 ;
        RECT 115.715 124.985 116.005 125.030 ;
        RECT 81.890 124.970 82.210 124.985 ;
        RECT 116.390 124.970 116.710 125.030 ;
        RECT 117.720 125.170 118.010 125.215 ;
        RECT 118.690 125.170 119.010 125.230 ;
        RECT 121.900 125.215 122.115 125.370 ;
        RECT 124.670 125.310 124.990 125.570 ;
        RECT 120.980 125.170 121.270 125.215 ;
        RECT 117.720 125.030 121.270 125.170 ;
        RECT 117.720 124.985 118.010 125.030 ;
        RECT 118.690 124.970 119.010 125.030 ;
        RECT 120.980 124.985 121.270 125.030 ;
        RECT 121.900 125.170 122.190 125.215 ;
        RECT 123.760 125.170 124.050 125.215 ;
        RECT 121.900 125.030 124.050 125.170 ;
        RECT 121.900 124.985 122.190 125.030 ;
        RECT 123.760 124.985 124.050 125.030 ;
        RECT 26.245 124.830 26.535 124.875 ;
        RECT 26.690 124.830 27.010 124.890 ;
        RECT 26.245 124.690 27.010 124.830 ;
        RECT 26.245 124.645 26.535 124.690 ;
        RECT 26.690 124.630 27.010 124.690 ;
        RECT 34.510 124.630 34.830 124.890 ;
        RECT 34.970 124.630 35.290 124.890 ;
        RECT 36.825 124.830 37.115 124.875 ;
        RECT 37.270 124.830 37.590 124.890 ;
        RECT 36.825 124.690 37.590 124.830 ;
        RECT 36.825 124.645 37.115 124.690 ;
        RECT 37.270 124.630 37.590 124.690 ;
        RECT 42.345 124.830 42.635 124.875 ;
        RECT 44.170 124.830 44.490 124.890 ;
        RECT 42.345 124.690 44.490 124.830 ;
        RECT 42.345 124.645 42.635 124.690 ;
        RECT 44.170 124.630 44.490 124.690 ;
        RECT 46.470 124.830 46.790 124.890 ;
        RECT 47.865 124.830 48.155 124.875 ;
        RECT 46.470 124.690 48.155 124.830 ;
        RECT 46.470 124.630 46.790 124.690 ;
        RECT 47.865 124.645 48.155 124.690 ;
        RECT 57.510 124.630 57.830 124.890 ;
        RECT 61.665 124.830 61.955 124.875 ;
        RECT 63.490 124.830 63.810 124.890 ;
        RECT 61.665 124.690 63.810 124.830 ;
        RECT 61.665 124.645 61.955 124.690 ;
        RECT 63.490 124.630 63.810 124.690 ;
        RECT 63.965 124.830 64.255 124.875 ;
        RECT 69.930 124.830 70.250 124.890 ;
        RECT 63.965 124.690 70.250 124.830 ;
        RECT 63.965 124.645 64.255 124.690 ;
        RECT 69.930 124.630 70.250 124.690 ;
        RECT 109.030 124.630 109.350 124.890 ;
        RECT 110.885 124.830 111.175 124.875 ;
        RECT 120.530 124.830 120.850 124.890 ;
        RECT 110.885 124.690 120.850 124.830 ;
        RECT 110.885 124.645 111.175 124.690 ;
        RECT 120.530 124.630 120.850 124.690 ;
        RECT 53.155 123.810 53.445 123.855 ;
        RECT 56.130 123.810 56.450 123.870 ;
        RECT 53.155 123.670 56.450 123.810 ;
        RECT 53.155 123.625 53.445 123.670 ;
        RECT 56.130 123.610 56.450 123.670 ;
        RECT 63.950 123.810 64.270 123.870 ;
        RECT 65.345 123.810 65.635 123.855 ;
        RECT 63.950 123.670 65.635 123.810 ;
        RECT 63.950 123.610 64.270 123.670 ;
        RECT 65.345 123.625 65.635 123.670 ;
        RECT 81.890 123.610 82.210 123.870 ;
        RECT 83.730 123.810 84.050 123.870 ;
        RECT 84.205 123.810 84.495 123.855 ;
        RECT 83.730 123.670 84.495 123.810 ;
        RECT 83.730 123.610 84.050 123.670 ;
        RECT 84.205 123.625 84.495 123.670 ;
        RECT 111.790 123.610 112.110 123.870 ;
        RECT 26.230 123.470 26.550 123.530 ;
        RECT 28.085 123.470 28.375 123.515 ;
        RECT 26.230 123.330 28.375 123.470 ;
        RECT 26.230 123.270 26.550 123.330 ;
        RECT 28.085 123.285 28.375 123.330 ;
        RECT 36.810 123.270 37.130 123.530 ;
        RECT 55.160 123.470 55.450 123.515 ;
        RECT 56.590 123.470 56.910 123.530 ;
        RECT 58.420 123.470 58.710 123.515 ;
        RECT 55.160 123.330 58.710 123.470 ;
        RECT 55.160 123.285 55.450 123.330 ;
        RECT 56.590 123.270 56.910 123.330 ;
        RECT 58.420 123.285 58.710 123.330 ;
        RECT 59.340 123.470 59.630 123.515 ;
        RECT 61.200 123.470 61.490 123.515 ;
        RECT 59.340 123.330 61.490 123.470 ;
        RECT 59.340 123.285 59.630 123.330 ;
        RECT 61.200 123.285 61.490 123.330 ;
        RECT 17.045 123.130 17.335 123.175 ;
        RECT 18.870 123.130 19.190 123.190 ;
        RECT 17.045 122.990 19.190 123.130 ;
        RECT 17.045 122.945 17.335 122.990 ;
        RECT 18.870 122.930 19.190 122.990 ;
        RECT 34.510 123.130 34.830 123.190 ;
        RECT 39.585 123.130 39.875 123.175 ;
        RECT 34.510 122.990 39.875 123.130 ;
        RECT 34.510 122.930 34.830 122.990 ;
        RECT 39.585 122.945 39.875 122.990 ;
        RECT 57.020 123.130 57.310 123.175 ;
        RECT 59.340 123.130 59.555 123.285 ;
        RECT 89.250 123.270 89.570 123.530 ;
        RECT 105.350 123.270 105.670 123.530 ;
        RECT 117.720 123.470 118.010 123.515 ;
        RECT 119.150 123.470 119.470 123.530 ;
        RECT 120.980 123.470 121.270 123.515 ;
        RECT 117.720 123.330 121.270 123.470 ;
        RECT 117.720 123.285 118.010 123.330 ;
        RECT 119.150 123.270 119.470 123.330 ;
        RECT 120.980 123.285 121.270 123.330 ;
        RECT 121.900 123.470 122.190 123.515 ;
        RECT 123.760 123.470 124.050 123.515 ;
        RECT 121.900 123.330 124.050 123.470 ;
        RECT 121.900 123.285 122.190 123.330 ;
        RECT 123.760 123.285 124.050 123.330 ;
        RECT 57.020 122.990 59.555 123.130 ;
        RECT 57.020 122.945 57.310 122.990 ;
        RECT 60.270 122.930 60.590 123.190 ;
        RECT 73.610 123.130 73.930 123.190 ;
        RECT 82.350 123.130 82.670 123.190 ;
        RECT 73.610 122.990 82.670 123.130 ;
        RECT 73.610 122.930 73.930 122.990 ;
        RECT 82.350 122.930 82.670 122.990 ;
        RECT 83.270 122.930 83.590 123.190 ;
        RECT 119.580 123.130 119.870 123.175 ;
        RECT 121.900 123.130 122.115 123.285 ;
        RECT 119.580 122.990 122.115 123.130 ;
        RECT 122.845 123.130 123.135 123.175 ;
        RECT 124.210 123.130 124.530 123.190 ;
        RECT 122.845 122.990 124.530 123.130 ;
        RECT 119.580 122.945 119.870 122.990 ;
        RECT 122.845 122.945 123.135 122.990 ;
        RECT 124.210 122.930 124.530 122.990 ;
        RECT 37.730 122.790 38.050 122.850 ;
        RECT 38.205 122.790 38.495 122.835 ;
        RECT 37.730 122.650 38.495 122.790 ;
        RECT 37.730 122.590 38.050 122.650 ;
        RECT 38.205 122.605 38.495 122.650 ;
        RECT 39.110 122.590 39.430 122.850 ;
        RECT 57.510 122.790 57.830 122.850 ;
        RECT 62.125 122.790 62.415 122.835 ;
        RECT 57.510 122.650 62.415 122.790 ;
        RECT 57.510 122.590 57.830 122.650 ;
        RECT 62.125 122.605 62.415 122.650 ;
        RECT 64.410 122.590 64.730 122.850 ;
        RECT 64.870 122.590 65.190 122.850 ;
        RECT 98.005 122.790 98.295 122.835 ;
        RECT 98.450 122.790 98.770 122.850 ;
        RECT 98.005 122.650 98.770 122.790 ;
        RECT 98.005 122.605 98.295 122.650 ;
        RECT 98.450 122.590 98.770 122.650 ;
        RECT 111.790 122.790 112.110 122.850 ;
        RECT 118.230 122.790 118.550 122.850 ;
        RECT 124.670 122.790 124.990 122.850 ;
        RECT 111.790 122.650 124.990 122.790 ;
        RECT 111.790 122.590 112.110 122.650 ;
        RECT 118.230 122.590 118.550 122.650 ;
        RECT 124.670 122.590 124.990 122.650 ;
        RECT 31.290 122.450 31.610 122.510 ;
        RECT 45.550 122.450 45.870 122.510 ;
        RECT 50.150 122.450 50.470 122.510 ;
        RECT 31.290 122.310 50.470 122.450 ;
        RECT 31.290 122.250 31.610 122.310 ;
        RECT 45.550 122.250 45.870 122.310 ;
        RECT 50.150 122.250 50.470 122.310 ;
        RECT 57.020 122.450 57.310 122.495 ;
        RECT 59.800 122.450 60.090 122.495 ;
        RECT 61.660 122.450 61.950 122.495 ;
        RECT 57.020 122.310 61.950 122.450 ;
        RECT 57.020 122.265 57.310 122.310 ;
        RECT 59.800 122.265 60.090 122.310 ;
        RECT 61.660 122.265 61.950 122.310 ;
        RECT 62.570 122.450 62.890 122.510 ;
        RECT 73.150 122.450 73.470 122.510 ;
        RECT 62.570 122.310 73.470 122.450 ;
        RECT 62.570 122.250 62.890 122.310 ;
        RECT 73.150 122.250 73.470 122.310 ;
        RECT 119.580 122.450 119.870 122.495 ;
        RECT 122.360 122.450 122.650 122.495 ;
        RECT 124.220 122.450 124.510 122.495 ;
        RECT 119.580 122.310 124.510 122.450 ;
        RECT 119.580 122.265 119.870 122.310 ;
        RECT 122.360 122.265 122.650 122.310 ;
        RECT 124.220 122.265 124.510 122.310 ;
        RECT 23.930 122.110 24.250 122.170 ;
        RECT 24.405 122.110 24.695 122.155 ;
        RECT 23.930 121.970 24.695 122.110 ;
        RECT 23.930 121.910 24.250 121.970 ;
        RECT 24.405 121.925 24.695 121.970 ;
        RECT 41.410 121.910 41.730 122.170 ;
        RECT 67.185 122.110 67.475 122.155 ;
        RECT 68.090 122.110 68.410 122.170 ;
        RECT 67.185 121.970 68.410 122.110 ;
        RECT 67.185 121.925 67.475 121.970 ;
        RECT 68.090 121.910 68.410 121.970 ;
        RECT 109.030 122.110 109.350 122.170 ;
        RECT 112.710 122.110 113.030 122.170 ;
        RECT 115.715 122.110 116.005 122.155 ;
        RECT 109.030 121.970 116.005 122.110 ;
        RECT 109.030 121.910 109.350 121.970 ;
        RECT 112.710 121.910 113.030 121.970 ;
        RECT 115.715 121.925 116.005 121.970 ;
        RECT 32.455 121.090 32.745 121.135 ;
        RECT 34.510 121.090 34.830 121.150 ;
        RECT 32.455 120.950 34.830 121.090 ;
        RECT 32.455 120.905 32.745 120.950 ;
        RECT 34.510 120.890 34.830 120.950 ;
        RECT 37.730 121.090 38.050 121.150 ;
        RECT 59.595 121.090 59.885 121.135 ;
        RECT 63.950 121.090 64.270 121.150 ;
        RECT 37.730 120.950 42.560 121.090 ;
        RECT 37.730 120.890 38.050 120.950 ;
        RECT 21.630 120.750 21.950 120.810 ;
        RECT 22.550 120.750 22.870 120.810 ;
        RECT 23.470 120.750 23.790 120.810 ;
        RECT 31.750 120.750 32.070 120.810 ;
        RECT 21.630 120.610 32.070 120.750 ;
        RECT 21.630 120.550 21.950 120.610 ;
        RECT 22.550 120.550 22.870 120.610 ;
        RECT 23.470 120.550 23.790 120.610 ;
        RECT 21.170 120.210 21.490 120.470 ;
        RECT 27.150 120.410 27.470 120.470 ;
        RECT 21.720 120.270 27.470 120.410 ;
        RECT 21.170 119.390 21.490 119.450 ;
        RECT 21.720 119.435 21.860 120.270 ;
        RECT 27.150 120.210 27.470 120.270 ;
        RECT 26.690 119.870 27.010 120.130 ;
        RECT 29.540 120.115 29.680 120.610 ;
        RECT 31.750 120.550 32.070 120.610 ;
        RECT 36.320 120.750 36.610 120.795 ;
        RECT 39.100 120.750 39.390 120.795 ;
        RECT 40.960 120.750 41.250 120.795 ;
        RECT 36.320 120.610 41.250 120.750 ;
        RECT 36.320 120.565 36.610 120.610 ;
        RECT 39.100 120.565 39.390 120.610 ;
        RECT 40.960 120.565 41.250 120.610 ;
        RECT 40.490 120.410 40.810 120.470 ;
        RECT 42.420 120.455 42.560 120.950 ;
        RECT 59.595 120.950 64.270 121.090 ;
        RECT 59.595 120.905 59.885 120.950 ;
        RECT 63.950 120.890 64.270 120.950 ;
        RECT 91.090 120.890 91.410 121.150 ;
        RECT 91.640 120.950 103.740 121.090 ;
        RECT 63.460 120.750 63.750 120.795 ;
        RECT 66.240 120.750 66.530 120.795 ;
        RECT 68.100 120.750 68.390 120.795 ;
        RECT 63.460 120.610 68.390 120.750 ;
        RECT 63.460 120.565 63.750 120.610 ;
        RECT 66.240 120.565 66.530 120.610 ;
        RECT 68.100 120.565 68.390 120.610 ;
        RECT 69.025 120.565 69.315 120.795 ;
        RECT 41.425 120.410 41.715 120.455 ;
        RECT 30.460 120.270 40.260 120.410 ;
        RECT 29.465 119.885 29.755 120.115 ;
        RECT 30.460 119.730 30.600 120.270 ;
        RECT 30.845 120.070 31.135 120.115 ;
        RECT 31.750 120.070 32.070 120.130 ;
        RECT 30.845 119.930 32.070 120.070 ;
        RECT 30.845 119.885 31.135 119.930 ;
        RECT 31.750 119.870 32.070 119.930 ;
        RECT 36.320 120.070 36.610 120.115 ;
        RECT 36.320 119.930 38.855 120.070 ;
        RECT 36.320 119.885 36.610 119.930 ;
        RECT 38.640 119.775 38.855 119.930 ;
        RECT 39.570 119.870 39.890 120.130 ;
        RECT 40.120 120.070 40.260 120.270 ;
        RECT 40.490 120.270 41.715 120.410 ;
        RECT 40.490 120.210 40.810 120.270 ;
        RECT 41.425 120.225 41.715 120.270 ;
        RECT 42.345 120.410 42.635 120.455 ;
        RECT 46.470 120.410 46.790 120.470 ;
        RECT 42.345 120.270 46.790 120.410 ;
        RECT 42.345 120.225 42.635 120.270 ;
        RECT 46.470 120.210 46.790 120.270 ;
        RECT 66.725 120.410 67.015 120.455 ;
        RECT 69.100 120.410 69.240 120.565 ;
        RECT 66.725 120.270 69.240 120.410 ;
        RECT 77.765 120.410 78.055 120.455 ;
        RECT 79.590 120.410 79.910 120.470 ;
        RECT 83.730 120.410 84.050 120.470 ;
        RECT 77.765 120.270 84.050 120.410 ;
        RECT 66.725 120.225 67.015 120.270 ;
        RECT 77.765 120.225 78.055 120.270 ;
        RECT 79.590 120.210 79.910 120.270 ;
        RECT 83.730 120.210 84.050 120.270 ;
        RECT 42.790 120.070 43.110 120.130 ;
        RECT 47.405 120.070 47.695 120.115 ;
        RECT 40.120 119.930 47.695 120.070 ;
        RECT 42.790 119.870 43.110 119.930 ;
        RECT 47.405 119.885 47.695 119.930 ;
        RECT 50.150 120.070 50.470 120.130 ;
        RECT 50.625 120.070 50.915 120.115 ;
        RECT 54.305 120.070 54.595 120.115 ;
        RECT 50.150 119.930 54.595 120.070 ;
        RECT 50.150 119.870 50.470 119.930 ;
        RECT 50.625 119.885 50.915 119.930 ;
        RECT 54.305 119.885 54.595 119.930 ;
        RECT 55.685 120.070 55.975 120.115 ;
        RECT 60.270 120.070 60.590 120.130 ;
        RECT 55.685 119.930 60.590 120.070 ;
        RECT 55.685 119.885 55.975 119.930 ;
        RECT 60.270 119.870 60.590 119.930 ;
        RECT 63.460 120.070 63.750 120.115 ;
        RECT 63.460 119.930 65.995 120.070 ;
        RECT 63.460 119.885 63.750 119.930 ;
        RECT 22.180 119.590 30.600 119.730 ;
        RECT 31.305 119.730 31.595 119.775 ;
        RECT 34.460 119.730 34.750 119.775 ;
        RECT 37.720 119.730 38.010 119.775 ;
        RECT 31.305 119.590 38.010 119.730 ;
        RECT 22.180 119.450 22.320 119.590 ;
        RECT 31.305 119.545 31.595 119.590 ;
        RECT 34.460 119.545 34.750 119.590 ;
        RECT 37.720 119.545 38.010 119.590 ;
        RECT 38.640 119.730 38.930 119.775 ;
        RECT 40.500 119.730 40.790 119.775 ;
        RECT 38.640 119.590 40.790 119.730 ;
        RECT 38.640 119.545 38.930 119.590 ;
        RECT 40.500 119.545 40.790 119.590 ;
        RECT 43.265 119.730 43.555 119.775 ;
        RECT 47.850 119.730 48.170 119.790 ;
        RECT 43.265 119.590 48.170 119.730 ;
        RECT 43.265 119.545 43.555 119.590 ;
        RECT 47.850 119.530 48.170 119.590 ;
        RECT 57.510 119.730 57.830 119.790 ;
        RECT 58.905 119.730 59.195 119.775 ;
        RECT 57.510 119.590 59.195 119.730 ;
        RECT 57.510 119.530 57.830 119.590 ;
        RECT 58.905 119.545 59.195 119.590 ;
        RECT 61.600 119.730 61.890 119.775 ;
        RECT 62.110 119.730 62.430 119.790 ;
        RECT 65.780 119.775 65.995 119.930 ;
        RECT 68.565 119.885 68.855 120.115 ;
        RECT 64.860 119.730 65.150 119.775 ;
        RECT 61.600 119.590 65.150 119.730 ;
        RECT 61.600 119.545 61.890 119.590 ;
        RECT 21.645 119.390 21.935 119.435 ;
        RECT 21.170 119.250 21.935 119.390 ;
        RECT 21.170 119.190 21.490 119.250 ;
        RECT 21.645 119.205 21.935 119.250 ;
        RECT 22.090 119.190 22.410 119.450 ;
        RECT 23.010 119.390 23.330 119.450 ;
        RECT 23.945 119.390 24.235 119.435 ;
        RECT 23.010 119.250 24.235 119.390 ;
        RECT 23.010 119.190 23.330 119.250 ;
        RECT 23.945 119.205 24.235 119.250 ;
        RECT 25.310 119.390 25.630 119.450 ;
        RECT 25.785 119.390 26.075 119.435 ;
        RECT 25.310 119.250 26.075 119.390 ;
        RECT 25.310 119.190 25.630 119.250 ;
        RECT 25.785 119.205 26.075 119.250 ;
        RECT 29.925 119.390 30.215 119.435 ;
        RECT 30.370 119.390 30.690 119.450 ;
        RECT 29.925 119.250 30.690 119.390 ;
        RECT 29.925 119.205 30.215 119.250 ;
        RECT 30.370 119.190 30.690 119.250 ;
        RECT 39.110 119.390 39.430 119.450 ;
        RECT 43.725 119.390 44.015 119.435 ;
        RECT 39.110 119.250 44.015 119.390 ;
        RECT 39.110 119.190 39.430 119.250 ;
        RECT 43.725 119.205 44.015 119.250 ;
        RECT 45.565 119.390 45.855 119.435 ;
        RECT 48.770 119.390 49.090 119.450 ;
        RECT 45.565 119.250 49.090 119.390 ;
        RECT 45.565 119.205 45.855 119.250 ;
        RECT 48.770 119.190 49.090 119.250 ;
        RECT 49.690 119.190 50.010 119.450 ;
        RECT 51.070 119.190 51.390 119.450 ;
        RECT 58.980 119.390 59.120 119.545 ;
        RECT 62.110 119.530 62.430 119.590 ;
        RECT 64.860 119.545 65.150 119.590 ;
        RECT 65.780 119.730 66.070 119.775 ;
        RECT 67.640 119.730 67.930 119.775 ;
        RECT 65.780 119.590 67.930 119.730 ;
        RECT 65.780 119.545 66.070 119.590 ;
        RECT 67.640 119.545 67.930 119.590 ;
        RECT 68.640 119.450 68.780 119.885 ;
        RECT 69.930 119.870 70.250 120.130 ;
        RECT 73.610 120.070 73.930 120.130 ;
        RECT 74.545 120.070 74.835 120.115 ;
        RECT 73.610 119.930 74.835 120.070 ;
        RECT 73.610 119.870 73.930 119.930 ;
        RECT 74.545 119.885 74.835 119.930 ;
        RECT 78.225 120.070 78.515 120.115 ;
        RECT 78.670 120.070 78.990 120.130 ;
        RECT 81.905 120.070 82.195 120.115 ;
        RECT 78.225 119.930 78.990 120.070 ;
        RECT 78.225 119.885 78.515 119.930 ;
        RECT 78.670 119.870 78.990 119.930 ;
        RECT 80.600 119.930 82.195 120.070 ;
        RECT 68.550 119.390 68.870 119.450 ;
        RECT 58.980 119.250 68.870 119.390 ;
        RECT 68.550 119.190 68.870 119.250 ;
        RECT 75.005 119.390 75.295 119.435 ;
        RECT 75.450 119.390 75.770 119.450 ;
        RECT 75.005 119.250 75.770 119.390 ;
        RECT 75.005 119.205 75.295 119.250 ;
        RECT 75.450 119.190 75.770 119.250 ;
        RECT 78.210 119.390 78.530 119.450 ;
        RECT 80.600 119.435 80.740 119.930 ;
        RECT 81.905 119.885 82.195 119.930 ;
        RECT 82.350 120.070 82.670 120.130 ;
        RECT 83.285 120.070 83.575 120.115 ;
        RECT 82.350 119.930 83.575 120.070 ;
        RECT 82.350 119.870 82.670 119.930 ;
        RECT 83.285 119.885 83.575 119.930 ;
        RECT 83.360 119.730 83.500 119.885 ;
        RECT 84.190 119.870 84.510 120.130 ;
        RECT 89.265 119.885 89.555 120.115 ;
        RECT 90.645 120.070 90.935 120.115 ;
        RECT 91.640 120.070 91.780 120.950 ;
        RECT 96.120 120.750 96.410 120.795 ;
        RECT 98.900 120.750 99.190 120.795 ;
        RECT 100.760 120.750 101.050 120.795 ;
        RECT 96.120 120.610 101.050 120.750 ;
        RECT 96.120 120.565 96.410 120.610 ;
        RECT 98.900 120.565 99.190 120.610 ;
        RECT 100.760 120.565 101.050 120.610 ;
        RECT 102.145 120.565 102.435 120.795 ;
        RECT 103.600 120.750 103.740 120.950 ;
        RECT 119.150 120.890 119.470 121.150 ;
        RECT 121.465 121.090 121.755 121.135 ;
        RECT 124.210 121.090 124.530 121.150 ;
        RECT 121.465 120.950 124.530 121.090 ;
        RECT 121.465 120.905 121.755 120.950 ;
        RECT 124.210 120.890 124.530 120.950 ;
        RECT 113.140 120.750 113.430 120.795 ;
        RECT 115.920 120.750 116.210 120.795 ;
        RECT 117.780 120.750 118.070 120.795 ;
        RECT 103.600 120.610 106.500 120.750 ;
        RECT 92.255 120.410 92.545 120.455 ;
        RECT 97.530 120.410 97.850 120.470 ;
        RECT 92.255 120.270 97.850 120.410 ;
        RECT 92.255 120.225 92.545 120.270 ;
        RECT 97.530 120.210 97.850 120.270 ;
        RECT 99.385 120.410 99.675 120.455 ;
        RECT 102.220 120.410 102.360 120.565 ;
        RECT 99.385 120.270 102.360 120.410 ;
        RECT 99.385 120.225 99.675 120.270 ;
        RECT 90.645 119.930 91.780 120.070 ;
        RECT 96.120 120.070 96.410 120.115 ;
        RECT 98.910 120.070 99.230 120.130 ;
        RECT 101.225 120.070 101.515 120.115 ;
        RECT 96.120 119.930 98.655 120.070 ;
        RECT 90.645 119.885 90.935 119.930 ;
        RECT 96.120 119.885 96.410 119.930 ;
        RECT 87.410 119.730 87.730 119.790 ;
        RECT 89.340 119.730 89.480 119.885 ;
        RECT 98.440 119.775 98.655 119.930 ;
        RECT 98.910 119.930 101.515 120.070 ;
        RECT 98.910 119.870 99.230 119.930 ;
        RECT 101.225 119.885 101.515 119.930 ;
        RECT 103.050 119.870 103.370 120.130 ;
        RECT 103.600 120.115 103.740 120.610 ;
        RECT 105.810 120.210 106.130 120.470 ;
        RECT 106.360 120.410 106.500 120.610 ;
        RECT 113.140 120.610 118.070 120.750 ;
        RECT 113.140 120.565 113.430 120.610 ;
        RECT 115.920 120.565 116.210 120.610 ;
        RECT 117.780 120.565 118.070 120.610 ;
        RECT 106.360 120.270 117.080 120.410 ;
        RECT 116.940 120.130 117.080 120.270 ;
        RECT 118.230 120.210 118.550 120.470 ;
        RECT 103.525 119.885 103.815 120.115 ;
        RECT 104.890 120.070 105.210 120.130 ;
        RECT 106.745 120.070 107.035 120.115 ;
        RECT 104.890 119.930 107.035 120.070 ;
        RECT 104.890 119.870 105.210 119.930 ;
        RECT 106.745 119.885 107.035 119.930 ;
        RECT 113.140 120.070 113.430 120.115 ;
        RECT 113.140 119.930 115.675 120.070 ;
        RECT 113.140 119.885 113.430 119.930 ;
        RECT 83.360 119.590 89.480 119.730 ;
        RECT 89.725 119.730 90.015 119.775 ;
        RECT 94.260 119.730 94.550 119.775 ;
        RECT 97.520 119.730 97.810 119.775 ;
        RECT 89.725 119.590 97.810 119.730 ;
        RECT 87.410 119.530 87.730 119.590 ;
        RECT 89.725 119.545 90.015 119.590 ;
        RECT 94.260 119.545 94.550 119.590 ;
        RECT 97.520 119.545 97.810 119.590 ;
        RECT 98.440 119.730 98.730 119.775 ;
        RECT 100.300 119.730 100.590 119.775 ;
        RECT 109.275 119.730 109.565 119.775 ;
        RECT 110.410 119.730 110.730 119.790 ;
        RECT 98.440 119.590 100.590 119.730 ;
        RECT 98.440 119.545 98.730 119.590 ;
        RECT 100.300 119.545 100.590 119.590 ;
        RECT 106.360 119.590 110.730 119.730 ;
        RECT 106.360 119.450 106.500 119.590 ;
        RECT 109.275 119.545 109.565 119.590 ;
        RECT 110.410 119.530 110.730 119.590 ;
        RECT 111.280 119.730 111.570 119.775 ;
        RECT 113.630 119.730 113.950 119.790 ;
        RECT 115.460 119.775 115.675 119.930 ;
        RECT 116.390 119.870 116.710 120.130 ;
        RECT 116.850 120.070 117.170 120.130 ;
        RECT 118.705 120.070 118.995 120.115 ;
        RECT 116.850 119.930 118.995 120.070 ;
        RECT 116.850 119.870 117.170 119.930 ;
        RECT 118.705 119.885 118.995 119.930 ;
        RECT 120.530 119.870 120.850 120.130 ;
        RECT 114.540 119.730 114.830 119.775 ;
        RECT 111.280 119.590 114.830 119.730 ;
        RECT 111.280 119.545 111.570 119.590 ;
        RECT 113.630 119.530 113.950 119.590 ;
        RECT 114.540 119.545 114.830 119.590 ;
        RECT 115.460 119.730 115.750 119.775 ;
        RECT 117.320 119.730 117.610 119.775 ;
        RECT 115.460 119.590 117.610 119.730 ;
        RECT 115.460 119.545 115.750 119.590 ;
        RECT 117.320 119.545 117.610 119.590 ;
        RECT 78.685 119.390 78.975 119.435 ;
        RECT 78.210 119.250 78.975 119.390 ;
        RECT 78.210 119.190 78.530 119.250 ;
        RECT 78.685 119.205 78.975 119.250 ;
        RECT 80.525 119.205 80.815 119.435 ;
        RECT 80.970 119.190 81.290 119.450 ;
        RECT 82.810 119.190 83.130 119.450 ;
        RECT 84.650 119.390 84.970 119.450 ;
        RECT 85.125 119.390 85.415 119.435 ;
        RECT 84.650 119.250 85.415 119.390 ;
        RECT 84.650 119.190 84.970 119.250 ;
        RECT 85.125 119.205 85.415 119.250 ;
        RECT 103.970 119.190 104.290 119.450 ;
        RECT 106.270 119.190 106.590 119.450 ;
        RECT 108.585 119.390 108.875 119.435 ;
        RECT 109.950 119.390 110.270 119.450 ;
        RECT 108.585 119.250 110.270 119.390 ;
        RECT 108.585 119.205 108.875 119.250 ;
        RECT 109.950 119.190 110.270 119.250 ;
        RECT 18.195 118.370 18.485 118.415 ;
        RECT 21.170 118.370 21.490 118.430 ;
        RECT 18.195 118.230 21.490 118.370 ;
        RECT 18.195 118.185 18.485 118.230 ;
        RECT 21.170 118.170 21.490 118.230 ;
        RECT 27.855 118.370 28.145 118.415 ;
        RECT 34.970 118.370 35.290 118.430 ;
        RECT 27.855 118.230 35.290 118.370 ;
        RECT 27.855 118.185 28.145 118.230 ;
        RECT 34.970 118.170 35.290 118.230 ;
        RECT 37.975 118.370 38.265 118.415 ;
        RECT 39.110 118.370 39.430 118.430 ;
        RECT 47.850 118.415 48.170 118.430 ;
        RECT 37.975 118.230 39.430 118.370 ;
        RECT 37.975 118.185 38.265 118.230 ;
        RECT 39.110 118.170 39.430 118.230 ;
        RECT 47.635 118.185 48.170 118.415 ;
        RECT 47.850 118.170 48.170 118.185 ;
        RECT 56.590 118.370 56.910 118.430 ;
        RECT 57.525 118.370 57.815 118.415 ;
        RECT 56.590 118.230 57.815 118.370 ;
        RECT 56.590 118.170 56.910 118.230 ;
        RECT 57.525 118.185 57.815 118.230 ;
        RECT 62.110 118.170 62.430 118.430 ;
        RECT 63.735 118.370 64.025 118.415 ;
        RECT 64.870 118.370 65.190 118.430 ;
        RECT 63.735 118.230 65.190 118.370 ;
        RECT 63.735 118.185 64.025 118.230 ;
        RECT 64.870 118.170 65.190 118.230 ;
        RECT 73.395 118.370 73.685 118.415 ;
        RECT 78.210 118.370 78.530 118.430 ;
        RECT 73.395 118.230 78.530 118.370 ;
        RECT 73.395 118.185 73.685 118.230 ;
        RECT 78.210 118.170 78.530 118.230 ;
        RECT 82.825 118.370 83.115 118.415 ;
        RECT 84.190 118.370 84.510 118.430 ;
        RECT 82.825 118.230 84.510 118.370 ;
        RECT 82.825 118.185 83.115 118.230 ;
        RECT 84.190 118.170 84.510 118.230 ;
        RECT 85.110 118.370 85.430 118.430 ;
        RECT 89.710 118.415 90.030 118.430 ;
        RECT 89.495 118.370 90.030 118.415 ;
        RECT 85.110 118.230 90.030 118.370 ;
        RECT 85.110 118.170 85.430 118.230 ;
        RECT 89.495 118.185 90.030 118.230 ;
        RECT 89.710 118.170 90.030 118.185 ;
        RECT 98.910 118.370 99.230 118.430 ;
        RECT 101.455 118.370 101.745 118.415 ;
        RECT 104.890 118.370 105.210 118.430 ;
        RECT 98.910 118.230 105.210 118.370 ;
        RECT 98.910 118.170 99.230 118.230 ;
        RECT 101.455 118.185 101.745 118.230 ;
        RECT 104.890 118.170 105.210 118.230 ;
        RECT 113.185 118.370 113.475 118.415 ;
        RECT 113.630 118.370 113.950 118.430 ;
        RECT 113.185 118.230 113.950 118.370 ;
        RECT 113.185 118.185 113.475 118.230 ;
        RECT 113.630 118.170 113.950 118.230 ;
        RECT 116.390 118.170 116.710 118.430 ;
        RECT 20.200 118.030 20.490 118.075 ;
        RECT 21.630 118.030 21.950 118.090 ;
        RECT 23.460 118.030 23.750 118.075 ;
        RECT 20.200 117.890 23.750 118.030 ;
        RECT 20.200 117.845 20.490 117.890 ;
        RECT 21.630 117.830 21.950 117.890 ;
        RECT 23.460 117.845 23.750 117.890 ;
        RECT 24.380 118.030 24.670 118.075 ;
        RECT 26.240 118.030 26.530 118.075 ;
        RECT 24.380 117.890 26.530 118.030 ;
        RECT 24.380 117.845 24.670 117.890 ;
        RECT 26.240 117.845 26.530 117.890 ;
        RECT 29.860 118.030 30.150 118.075 ;
        RECT 30.370 118.030 30.690 118.090 ;
        RECT 43.250 118.075 43.570 118.090 ;
        RECT 33.120 118.030 33.410 118.075 ;
        RECT 29.860 117.890 33.410 118.030 ;
        RECT 29.860 117.845 30.150 117.890 ;
        RECT 22.060 117.690 22.350 117.735 ;
        RECT 24.380 117.690 24.595 117.845 ;
        RECT 30.370 117.830 30.690 117.890 ;
        RECT 33.120 117.845 33.410 117.890 ;
        RECT 34.040 118.030 34.330 118.075 ;
        RECT 35.900 118.030 36.190 118.075 ;
        RECT 34.040 117.890 36.190 118.030 ;
        RECT 34.040 117.845 34.330 117.890 ;
        RECT 35.900 117.845 36.190 117.890 ;
        RECT 39.980 118.030 40.270 118.075 ;
        RECT 43.240 118.030 43.570 118.075 ;
        RECT 39.980 117.890 43.570 118.030 ;
        RECT 39.980 117.845 40.270 117.890 ;
        RECT 43.240 117.845 43.570 117.890 ;
        RECT 22.060 117.550 24.595 117.690 ;
        RECT 22.060 117.505 22.350 117.550 ;
        RECT 25.310 117.490 25.630 117.750 ;
        RECT 26.690 117.690 27.010 117.750 ;
        RECT 27.165 117.690 27.455 117.735 ;
        RECT 26.690 117.550 27.455 117.690 ;
        RECT 26.690 117.490 27.010 117.550 ;
        RECT 27.165 117.505 27.455 117.550 ;
        RECT 31.720 117.690 32.010 117.735 ;
        RECT 34.040 117.690 34.255 117.845 ;
        RECT 43.250 117.830 43.570 117.845 ;
        RECT 44.160 118.030 44.450 118.075 ;
        RECT 46.020 118.030 46.310 118.075 ;
        RECT 44.160 117.890 46.310 118.030 ;
        RECT 44.160 117.845 44.450 117.890 ;
        RECT 46.020 117.845 46.310 117.890 ;
        RECT 49.640 118.030 49.930 118.075 ;
        RECT 51.070 118.030 51.390 118.090 ;
        RECT 52.900 118.030 53.190 118.075 ;
        RECT 49.640 117.890 53.190 118.030 ;
        RECT 49.640 117.845 49.930 117.890 ;
        RECT 31.720 117.550 34.255 117.690 ;
        RECT 36.825 117.690 37.115 117.735 ;
        RECT 38.190 117.690 38.510 117.750 ;
        RECT 40.490 117.690 40.810 117.750 ;
        RECT 36.825 117.550 40.810 117.690 ;
        RECT 31.720 117.505 32.010 117.550 ;
        RECT 36.825 117.505 37.115 117.550 ;
        RECT 38.190 117.490 38.510 117.550 ;
        RECT 40.490 117.490 40.810 117.550 ;
        RECT 41.840 117.690 42.130 117.735 ;
        RECT 44.160 117.690 44.375 117.845 ;
        RECT 51.070 117.830 51.390 117.890 ;
        RECT 52.900 117.845 53.190 117.890 ;
        RECT 53.820 118.030 54.110 118.075 ;
        RECT 55.680 118.030 55.970 118.075 ;
        RECT 53.820 117.890 55.970 118.030 ;
        RECT 53.820 117.845 54.110 117.890 ;
        RECT 55.680 117.845 55.970 117.890 ;
        RECT 65.740 118.030 66.030 118.075 ;
        RECT 66.250 118.030 66.570 118.090 ;
        RECT 75.450 118.075 75.770 118.090 ;
        RECT 69.000 118.030 69.290 118.075 ;
        RECT 65.740 117.890 69.290 118.030 ;
        RECT 65.740 117.845 66.030 117.890 ;
        RECT 41.840 117.550 44.375 117.690 ;
        RECT 41.840 117.505 42.130 117.550 ;
        RECT 45.090 117.490 45.410 117.750 ;
        RECT 51.500 117.690 51.790 117.735 ;
        RECT 53.820 117.690 54.035 117.845 ;
        RECT 66.250 117.830 66.570 117.890 ;
        RECT 69.000 117.845 69.290 117.890 ;
        RECT 69.920 118.030 70.210 118.075 ;
        RECT 71.780 118.030 72.070 118.075 ;
        RECT 69.920 117.890 72.070 118.030 ;
        RECT 69.920 117.845 70.210 117.890 ;
        RECT 71.780 117.845 72.070 117.890 ;
        RECT 75.400 118.030 75.770 118.075 ;
        RECT 78.660 118.030 78.950 118.075 ;
        RECT 75.400 117.890 78.950 118.030 ;
        RECT 75.400 117.845 75.770 117.890 ;
        RECT 78.660 117.845 78.950 117.890 ;
        RECT 79.580 118.030 79.870 118.075 ;
        RECT 81.440 118.030 81.730 118.075 ;
        RECT 84.665 118.030 84.955 118.075 ;
        RECT 79.580 117.890 81.730 118.030 ;
        RECT 79.580 117.845 79.870 117.890 ;
        RECT 81.440 117.845 81.730 117.890 ;
        RECT 81.980 117.890 84.955 118.030 ;
        RECT 51.500 117.550 54.035 117.690 ;
        RECT 57.985 117.690 58.275 117.735 ;
        RECT 60.270 117.690 60.590 117.750 ;
        RECT 61.665 117.690 61.955 117.735 ;
        RECT 63.950 117.690 64.270 117.750 ;
        RECT 57.985 117.550 64.270 117.690 ;
        RECT 51.500 117.505 51.790 117.550 ;
        RECT 57.985 117.505 58.275 117.550 ;
        RECT 60.270 117.490 60.590 117.550 ;
        RECT 61.665 117.505 61.955 117.550 ;
        RECT 63.950 117.490 64.270 117.550 ;
        RECT 67.600 117.690 67.890 117.735 ;
        RECT 69.920 117.690 70.135 117.845 ;
        RECT 75.450 117.830 75.770 117.845 ;
        RECT 67.600 117.550 70.135 117.690 ;
        RECT 67.600 117.505 67.890 117.550 ;
        RECT 70.850 117.490 71.170 117.750 ;
        RECT 77.260 117.690 77.550 117.735 ;
        RECT 79.580 117.690 79.795 117.845 ;
        RECT 77.260 117.550 79.795 117.690 ;
        RECT 80.525 117.690 80.815 117.735 ;
        RECT 80.970 117.690 81.290 117.750 ;
        RECT 81.980 117.690 82.120 117.890 ;
        RECT 84.665 117.845 84.955 117.890 ;
        RECT 87.885 118.030 88.175 118.075 ;
        RECT 91.500 118.030 91.790 118.075 ;
        RECT 94.760 118.030 95.050 118.075 ;
        RECT 87.885 117.890 95.050 118.030 ;
        RECT 87.885 117.845 88.175 117.890 ;
        RECT 91.500 117.845 91.790 117.890 ;
        RECT 94.760 117.845 95.050 117.890 ;
        RECT 95.680 118.030 95.970 118.075 ;
        RECT 97.540 118.030 97.830 118.075 ;
        RECT 95.680 117.890 97.830 118.030 ;
        RECT 95.680 117.845 95.970 117.890 ;
        RECT 97.540 117.845 97.830 117.890 ;
        RECT 103.460 118.030 103.750 118.075 ;
        RECT 103.970 118.030 104.290 118.090 ;
        RECT 106.720 118.030 107.010 118.075 ;
        RECT 103.460 117.890 107.010 118.030 ;
        RECT 103.460 117.845 103.750 117.890 ;
        RECT 80.525 117.550 81.290 117.690 ;
        RECT 77.260 117.505 77.550 117.550 ;
        RECT 80.525 117.505 80.815 117.550 ;
        RECT 80.970 117.490 81.290 117.550 ;
        RECT 81.520 117.550 82.120 117.690 ;
        RECT 82.365 117.690 82.655 117.735 ;
        RECT 85.110 117.690 85.430 117.750 ;
        RECT 82.365 117.550 85.430 117.690 ;
        RECT 34.985 117.350 35.275 117.395 ;
        RECT 35.890 117.350 36.210 117.410 ;
        RECT 34.985 117.210 36.210 117.350 ;
        RECT 40.580 117.350 40.720 117.490 ;
        RECT 46.945 117.350 47.235 117.395 ;
        RECT 40.580 117.210 47.235 117.350 ;
        RECT 34.985 117.165 35.275 117.210 ;
        RECT 35.890 117.150 36.210 117.210 ;
        RECT 46.945 117.165 47.235 117.210 ;
        RECT 54.750 117.150 55.070 117.410 ;
        RECT 56.605 117.350 56.895 117.395 ;
        RECT 57.050 117.350 57.370 117.410 ;
        RECT 56.605 117.210 57.370 117.350 ;
        RECT 56.605 117.165 56.895 117.210 ;
        RECT 57.050 117.150 57.370 117.210 ;
        RECT 68.550 117.350 68.870 117.410 ;
        RECT 72.705 117.350 72.995 117.395 ;
        RECT 73.610 117.350 73.930 117.410 ;
        RECT 68.550 117.210 73.930 117.350 ;
        RECT 68.550 117.150 68.870 117.210 ;
        RECT 72.705 117.165 72.995 117.210 ;
        RECT 73.610 117.150 73.930 117.210 ;
        RECT 78.670 117.350 78.990 117.410 ;
        RECT 81.520 117.350 81.660 117.550 ;
        RECT 82.365 117.505 82.655 117.550 ;
        RECT 85.110 117.490 85.430 117.550 ;
        RECT 87.410 117.490 87.730 117.750 ;
        RECT 93.360 117.690 93.650 117.735 ;
        RECT 95.680 117.690 95.895 117.845 ;
        RECT 103.970 117.830 104.290 117.890 ;
        RECT 106.720 117.845 107.010 117.890 ;
        RECT 107.640 118.030 107.930 118.075 ;
        RECT 109.500 118.030 109.790 118.075 ;
        RECT 107.640 117.890 109.790 118.030 ;
        RECT 107.640 117.845 107.930 117.890 ;
        RECT 109.500 117.845 109.790 117.890 ;
        RECT 109.950 118.030 110.270 118.090 ;
        RECT 116.850 118.030 117.170 118.090 ;
        RECT 109.950 117.890 112.020 118.030 ;
        RECT 93.360 117.550 95.895 117.690 ;
        RECT 93.360 117.505 93.650 117.550 ;
        RECT 98.450 117.490 98.770 117.750 ;
        RECT 99.830 117.490 100.150 117.750 ;
        RECT 105.320 117.690 105.610 117.735 ;
        RECT 107.640 117.690 107.855 117.845 ;
        RECT 109.950 117.830 110.270 117.890 ;
        RECT 105.320 117.550 107.855 117.690 ;
        RECT 110.425 117.690 110.715 117.735 ;
        RECT 111.330 117.690 111.650 117.750 ;
        RECT 111.880 117.735 112.020 117.890 ;
        RECT 113.720 117.890 117.170 118.030 ;
        RECT 113.720 117.735 113.860 117.890 ;
        RECT 116.850 117.830 117.170 117.890 ;
        RECT 110.425 117.550 111.650 117.690 ;
        RECT 105.320 117.505 105.610 117.550 ;
        RECT 110.425 117.505 110.715 117.550 ;
        RECT 111.330 117.490 111.650 117.550 ;
        RECT 111.805 117.505 112.095 117.735 ;
        RECT 113.645 117.505 113.935 117.735 ;
        RECT 115.470 117.490 115.790 117.750 ;
        RECT 117.310 117.490 117.630 117.750 ;
        RECT 78.670 117.210 81.660 117.350 ;
        RECT 83.730 117.350 84.050 117.410 ;
        RECT 85.585 117.350 85.875 117.395 ;
        RECT 83.730 117.210 85.875 117.350 ;
        RECT 78.670 117.150 78.990 117.210 ;
        RECT 83.730 117.150 84.050 117.210 ;
        RECT 85.585 117.165 85.875 117.210 ;
        RECT 96.625 117.350 96.915 117.395 ;
        RECT 108.585 117.350 108.875 117.395 ;
        RECT 126.065 117.350 126.355 117.395 ;
        RECT 127.890 117.350 128.210 117.410 ;
        RECT 96.625 117.210 99.140 117.350 ;
        RECT 96.625 117.165 96.915 117.210 ;
        RECT 99.000 117.055 99.140 117.210 ;
        RECT 108.585 117.210 111.100 117.350 ;
        RECT 108.585 117.165 108.875 117.210 ;
        RECT 110.960 117.055 111.100 117.210 ;
        RECT 126.065 117.210 128.210 117.350 ;
        RECT 126.065 117.165 126.355 117.210 ;
        RECT 127.890 117.150 128.210 117.210 ;
        RECT 22.060 117.010 22.350 117.055 ;
        RECT 24.840 117.010 25.130 117.055 ;
        RECT 26.700 117.010 26.990 117.055 ;
        RECT 22.060 116.870 26.990 117.010 ;
        RECT 22.060 116.825 22.350 116.870 ;
        RECT 24.840 116.825 25.130 116.870 ;
        RECT 26.700 116.825 26.990 116.870 ;
        RECT 31.720 117.010 32.010 117.055 ;
        RECT 34.500 117.010 34.790 117.055 ;
        RECT 36.360 117.010 36.650 117.055 ;
        RECT 31.720 116.870 36.650 117.010 ;
        RECT 31.720 116.825 32.010 116.870 ;
        RECT 34.500 116.825 34.790 116.870 ;
        RECT 36.360 116.825 36.650 116.870 ;
        RECT 41.840 117.010 42.130 117.055 ;
        RECT 44.620 117.010 44.910 117.055 ;
        RECT 46.480 117.010 46.770 117.055 ;
        RECT 41.840 116.870 46.770 117.010 ;
        RECT 41.840 116.825 42.130 116.870 ;
        RECT 44.620 116.825 44.910 116.870 ;
        RECT 46.480 116.825 46.770 116.870 ;
        RECT 51.500 117.010 51.790 117.055 ;
        RECT 54.280 117.010 54.570 117.055 ;
        RECT 56.140 117.010 56.430 117.055 ;
        RECT 51.500 116.870 56.430 117.010 ;
        RECT 51.500 116.825 51.790 116.870 ;
        RECT 54.280 116.825 54.570 116.870 ;
        RECT 56.140 116.825 56.430 116.870 ;
        RECT 67.600 117.010 67.890 117.055 ;
        RECT 70.380 117.010 70.670 117.055 ;
        RECT 72.240 117.010 72.530 117.055 ;
        RECT 67.600 116.870 72.530 117.010 ;
        RECT 67.600 116.825 67.890 116.870 ;
        RECT 70.380 116.825 70.670 116.870 ;
        RECT 72.240 116.825 72.530 116.870 ;
        RECT 77.260 117.010 77.550 117.055 ;
        RECT 80.040 117.010 80.330 117.055 ;
        RECT 81.900 117.010 82.190 117.055 ;
        RECT 77.260 116.870 82.190 117.010 ;
        RECT 77.260 116.825 77.550 116.870 ;
        RECT 80.040 116.825 80.330 116.870 ;
        RECT 81.900 116.825 82.190 116.870 ;
        RECT 93.360 117.010 93.650 117.055 ;
        RECT 96.140 117.010 96.430 117.055 ;
        RECT 98.000 117.010 98.290 117.055 ;
        RECT 93.360 116.870 98.290 117.010 ;
        RECT 93.360 116.825 93.650 116.870 ;
        RECT 96.140 116.825 96.430 116.870 ;
        RECT 98.000 116.825 98.290 116.870 ;
        RECT 98.925 116.825 99.215 117.055 ;
        RECT 105.320 117.010 105.610 117.055 ;
        RECT 108.100 117.010 108.390 117.055 ;
        RECT 109.960 117.010 110.250 117.055 ;
        RECT 105.320 116.870 110.250 117.010 ;
        RECT 105.320 116.825 105.610 116.870 ;
        RECT 108.100 116.825 108.390 116.870 ;
        RECT 109.960 116.825 110.250 116.870 ;
        RECT 110.885 116.825 111.175 117.055 ;
        RECT 21.630 115.650 21.950 115.710 ;
        RECT 22.105 115.650 22.395 115.695 ;
        RECT 21.630 115.510 22.395 115.650 ;
        RECT 21.630 115.450 21.950 115.510 ;
        RECT 22.105 115.465 22.395 115.510 ;
        RECT 39.570 115.650 39.890 115.710 ;
        RECT 43.265 115.650 43.555 115.695 ;
        RECT 39.570 115.510 43.555 115.650 ;
        RECT 39.570 115.450 39.890 115.510 ;
        RECT 43.265 115.465 43.555 115.510 ;
        RECT 45.090 115.650 45.410 115.710 ;
        RECT 47.865 115.650 48.155 115.695 ;
        RECT 45.090 115.510 48.155 115.650 ;
        RECT 45.090 115.450 45.410 115.510 ;
        RECT 47.865 115.465 48.155 115.510 ;
        RECT 53.385 115.650 53.675 115.695 ;
        RECT 54.750 115.650 55.070 115.710 ;
        RECT 53.385 115.510 55.070 115.650 ;
        RECT 53.385 115.465 53.675 115.510 ;
        RECT 54.750 115.450 55.070 115.510 ;
        RECT 66.250 115.450 66.570 115.710 ;
        RECT 69.025 115.650 69.315 115.695 ;
        RECT 70.850 115.650 71.170 115.710 ;
        RECT 69.025 115.510 71.170 115.650 ;
        RECT 69.025 115.465 69.315 115.510 ;
        RECT 70.850 115.450 71.170 115.510 ;
        RECT 77.535 115.650 77.825 115.695 ;
        RECT 78.670 115.650 78.990 115.710 ;
        RECT 77.535 115.510 78.990 115.650 ;
        RECT 77.535 115.465 77.825 115.510 ;
        RECT 78.670 115.450 78.990 115.510 ;
        RECT 83.730 115.650 84.050 115.710 ;
        RECT 94.785 115.650 95.075 115.695 ;
        RECT 99.830 115.650 100.150 115.710 ;
        RECT 83.730 115.510 92.240 115.650 ;
        RECT 83.730 115.450 84.050 115.510 ;
        RECT 81.400 115.310 81.690 115.355 ;
        RECT 84.180 115.310 84.470 115.355 ;
        RECT 86.040 115.310 86.330 115.355 ;
        RECT 81.400 115.170 86.330 115.310 ;
        RECT 81.400 115.125 81.690 115.170 ;
        RECT 84.180 115.125 84.470 115.170 ;
        RECT 86.040 115.125 86.330 115.170 ;
        RECT 92.100 115.310 92.240 115.510 ;
        RECT 94.785 115.510 100.150 115.650 ;
        RECT 94.785 115.465 95.075 115.510 ;
        RECT 99.830 115.450 100.150 115.510 ;
        RECT 101.225 115.650 101.515 115.695 ;
        RECT 103.050 115.650 103.370 115.710 ;
        RECT 101.225 115.510 103.370 115.650 ;
        RECT 101.225 115.465 101.515 115.510 ;
        RECT 103.050 115.450 103.370 115.510 ;
        RECT 115.025 115.650 115.315 115.695 ;
        RECT 115.470 115.650 115.790 115.710 ;
        RECT 115.025 115.510 115.790 115.650 ;
        RECT 115.025 115.465 115.315 115.510 ;
        RECT 115.470 115.450 115.790 115.510 ;
        RECT 105.810 115.310 106.130 115.370 ;
        RECT 92.100 115.170 106.130 115.310 ;
        RECT 14.270 114.970 14.590 115.030 ;
        RECT 34.065 114.970 34.355 115.015 ;
        RECT 14.270 114.830 34.355 114.970 ;
        RECT 14.270 114.770 14.590 114.830 ;
        RECT 34.065 114.785 34.355 114.830 ;
        RECT 43.250 114.970 43.570 115.030 ;
        RECT 45.105 114.970 45.395 115.015 ;
        RECT 43.250 114.830 45.395 114.970 ;
        RECT 43.250 114.770 43.570 114.830 ;
        RECT 45.105 114.785 45.395 114.830 ;
        RECT 60.270 114.970 60.590 115.030 ;
        RECT 63.950 114.970 64.270 115.030 ;
        RECT 70.390 114.970 70.710 115.030 ;
        RECT 60.270 114.830 70.710 114.970 ;
        RECT 60.270 114.770 60.590 114.830 ;
        RECT 63.950 114.770 64.270 114.830 ;
        RECT 20.265 114.630 20.555 114.675 ;
        RECT 22.550 114.630 22.870 114.690 ;
        RECT 20.265 114.490 22.870 114.630 ;
        RECT 20.265 114.445 20.555 114.490 ;
        RECT 22.550 114.430 22.870 114.490 ;
        RECT 23.010 114.430 23.330 114.690 ;
        RECT 41.410 114.630 41.730 114.690 ;
        RECT 44.185 114.630 44.475 114.675 ;
        RECT 41.410 114.490 44.475 114.630 ;
        RECT 41.410 114.430 41.730 114.490 ;
        RECT 44.185 114.445 44.475 114.490 ;
        RECT 45.550 114.430 45.870 114.690 ;
        RECT 48.770 114.430 49.090 114.690 ;
        RECT 49.690 114.630 50.010 114.690 ;
        RECT 65.880 114.675 66.020 114.830 ;
        RECT 70.390 114.770 70.710 114.830 ;
        RECT 84.650 114.770 84.970 115.030 ;
        RECT 85.110 114.970 85.430 115.030 ;
        RECT 92.100 115.015 92.240 115.170 ;
        RECT 98.080 115.015 98.220 115.170 ;
        RECT 105.810 115.110 106.130 115.170 ;
        RECT 111.790 115.310 112.110 115.370 ;
        RECT 118.195 115.310 118.485 115.355 ;
        RECT 120.085 115.310 120.375 115.355 ;
        RECT 123.205 115.310 123.495 115.355 ;
        RECT 111.790 115.170 117.540 115.310 ;
        RECT 111.790 115.110 112.110 115.170 ;
        RECT 86.505 114.970 86.795 115.015 ;
        RECT 85.110 114.830 86.795 114.970 ;
        RECT 85.110 114.770 85.430 114.830 ;
        RECT 86.505 114.785 86.795 114.830 ;
        RECT 92.025 114.785 92.315 115.015 ;
        RECT 92.485 114.970 92.775 115.015 ;
        RECT 92.485 114.830 97.760 114.970 ;
        RECT 92.485 114.785 92.775 114.830 ;
        RECT 97.620 114.690 97.760 114.830 ;
        RECT 98.005 114.785 98.295 115.015 ;
        RECT 98.910 114.770 99.230 115.030 ;
        RECT 105.900 114.970 106.040 115.110 ;
        RECT 112.265 114.970 112.555 115.015 ;
        RECT 105.900 114.830 112.555 114.970 ;
        RECT 112.265 114.785 112.555 114.830 ;
        RECT 112.710 114.770 113.030 115.030 ;
        RECT 117.400 115.015 117.540 115.170 ;
        RECT 118.195 115.170 123.495 115.310 ;
        RECT 118.195 115.125 118.485 115.170 ;
        RECT 120.085 115.125 120.375 115.170 ;
        RECT 123.205 115.125 123.495 115.170 ;
        RECT 117.325 114.785 117.615 115.015 ;
        RECT 52.465 114.630 52.755 114.675 ;
        RECT 49.690 114.490 52.755 114.630 ;
        RECT 49.690 114.430 50.010 114.490 ;
        RECT 52.465 114.445 52.755 114.490 ;
        RECT 65.805 114.445 66.095 114.675 ;
        RECT 68.090 114.430 68.410 114.690 ;
        RECT 81.400 114.630 81.690 114.675 ;
        RECT 89.710 114.630 90.030 114.690 ;
        RECT 92.945 114.630 93.235 114.675 ;
        RECT 81.400 114.490 83.935 114.630 ;
        RECT 81.400 114.445 81.690 114.490 ;
        RECT 24.865 114.290 25.155 114.335 ;
        RECT 25.310 114.290 25.630 114.350 ;
        RECT 24.865 114.150 25.630 114.290 ;
        RECT 24.865 114.105 25.155 114.150 ;
        RECT 25.310 114.090 25.630 114.150 ;
        RECT 42.790 114.090 43.110 114.350 ;
        RECT 82.810 114.335 83.130 114.350 ;
        RECT 79.540 114.290 79.830 114.335 ;
        RECT 82.800 114.290 83.130 114.335 ;
        RECT 79.540 114.150 83.130 114.290 ;
        RECT 79.540 114.105 79.830 114.150 ;
        RECT 82.800 114.105 83.130 114.150 ;
        RECT 83.720 114.335 83.935 114.490 ;
        RECT 89.710 114.490 93.235 114.630 ;
        RECT 89.710 114.430 90.030 114.490 ;
        RECT 92.945 114.445 93.235 114.490 ;
        RECT 97.530 114.630 97.850 114.690 ;
        RECT 99.385 114.630 99.675 114.675 ;
        RECT 97.530 114.490 99.675 114.630 ;
        RECT 97.530 114.430 97.850 114.490 ;
        RECT 99.385 114.445 99.675 114.490 ;
        RECT 106.270 114.630 106.590 114.690 ;
        RECT 113.185 114.630 113.475 114.675 ;
        RECT 106.270 114.490 113.475 114.630 ;
        RECT 106.270 114.430 106.590 114.490 ;
        RECT 113.185 114.445 113.475 114.490 ;
        RECT 117.790 114.630 118.080 114.675 ;
        RECT 119.625 114.630 119.915 114.675 ;
        RECT 123.205 114.630 123.495 114.675 ;
        RECT 117.790 114.490 123.495 114.630 ;
        RECT 117.790 114.445 118.080 114.490 ;
        RECT 119.625 114.445 119.915 114.490 ;
        RECT 123.205 114.445 123.495 114.490 ;
        RECT 124.210 114.650 124.530 114.690 ;
        RECT 124.210 114.430 124.575 114.650 ;
        RECT 83.720 114.290 84.010 114.335 ;
        RECT 85.580 114.290 85.870 114.335 ;
        RECT 83.720 114.150 85.870 114.290 ;
        RECT 83.720 114.105 84.010 114.150 ;
        RECT 85.580 114.105 85.870 114.150 ;
        RECT 115.470 114.290 115.790 114.350 ;
        RECT 124.285 114.335 124.575 114.430 ;
        RECT 118.705 114.290 118.995 114.335 ;
        RECT 115.470 114.150 118.995 114.290 ;
        RECT 82.810 114.090 83.130 114.105 ;
        RECT 115.470 114.090 115.790 114.150 ;
        RECT 118.705 114.105 118.995 114.150 ;
        RECT 120.985 114.290 121.635 114.335 ;
        RECT 124.285 114.290 124.875 114.335 ;
        RECT 120.985 114.150 124.875 114.290 ;
        RECT 120.985 114.105 121.635 114.150 ;
        RECT 124.585 114.105 124.875 114.150 ;
        RECT 20.710 113.750 21.030 114.010 ;
        RECT 23.930 113.750 24.250 114.010 ;
        RECT 31.290 113.750 31.610 114.010 ;
        RECT 126.050 113.750 126.370 114.010 ;
        RECT 17.275 112.930 17.565 112.975 ;
        RECT 22.090 112.930 22.410 112.990 ;
        RECT 17.275 112.790 22.410 112.930 ;
        RECT 17.275 112.745 17.565 112.790 ;
        RECT 22.090 112.730 22.410 112.790 ;
        RECT 35.445 112.745 35.735 112.975 ;
        RECT 19.280 112.590 19.570 112.635 ;
        RECT 20.710 112.590 21.030 112.650 ;
        RECT 22.540 112.590 22.830 112.635 ;
        RECT 19.280 112.450 22.830 112.590 ;
        RECT 19.280 112.405 19.570 112.450 ;
        RECT 20.710 112.390 21.030 112.450 ;
        RECT 22.540 112.405 22.830 112.450 ;
        RECT 23.460 112.590 23.750 112.635 ;
        RECT 25.320 112.590 25.610 112.635 ;
        RECT 23.460 112.450 25.610 112.590 ;
        RECT 23.460 112.405 23.750 112.450 ;
        RECT 25.320 112.405 25.610 112.450 ;
        RECT 28.070 112.590 28.390 112.650 ;
        RECT 30.365 112.590 31.015 112.635 ;
        RECT 33.965 112.590 34.255 112.635 ;
        RECT 28.070 112.450 34.255 112.590 ;
        RECT 35.520 112.590 35.660 112.745 ;
        RECT 35.890 112.730 36.210 112.990 ;
        RECT 106.270 112.730 106.590 112.990 ;
        RECT 37.745 112.590 38.035 112.635 ;
        RECT 35.520 112.450 38.035 112.590 ;
        RECT 21.140 112.250 21.430 112.295 ;
        RECT 23.460 112.250 23.675 112.405 ;
        RECT 28.070 112.390 28.390 112.450 ;
        RECT 30.365 112.405 31.015 112.450 ;
        RECT 33.665 112.405 34.255 112.450 ;
        RECT 37.745 112.405 38.035 112.450 ;
        RECT 70.390 112.590 70.710 112.650 ;
        RECT 123.765 112.590 124.055 112.635 ;
        RECT 126.050 112.590 126.370 112.650 ;
        RECT 70.390 112.450 79.820 112.590 ;
        RECT 21.140 112.110 23.675 112.250 ;
        RECT 23.930 112.250 24.250 112.310 ;
        RECT 24.405 112.250 24.695 112.295 ;
        RECT 23.930 112.110 24.695 112.250 ;
        RECT 21.140 112.065 21.430 112.110 ;
        RECT 23.930 112.050 24.250 112.110 ;
        RECT 24.405 112.065 24.695 112.110 ;
        RECT 26.245 112.250 26.535 112.295 ;
        RECT 26.690 112.250 27.010 112.310 ;
        RECT 26.245 112.110 27.010 112.250 ;
        RECT 26.245 112.065 26.535 112.110 ;
        RECT 26.690 112.050 27.010 112.110 ;
        RECT 27.170 112.250 27.460 112.295 ;
        RECT 29.005 112.250 29.295 112.295 ;
        RECT 32.585 112.250 32.875 112.295 ;
        RECT 27.170 112.110 32.875 112.250 ;
        RECT 27.170 112.065 27.460 112.110 ;
        RECT 29.005 112.065 29.295 112.110 ;
        RECT 32.585 112.065 32.875 112.110 ;
        RECT 33.665 112.090 33.955 112.405 ;
        RECT 70.390 112.390 70.710 112.450 ;
        RECT 36.825 112.250 37.115 112.295 ;
        RECT 37.270 112.250 37.590 112.310 ;
        RECT 36.825 112.110 37.590 112.250 ;
        RECT 36.825 112.065 37.115 112.110 ;
        RECT 37.270 112.050 37.590 112.110 ;
        RECT 79.130 112.050 79.450 112.310 ;
        RECT 79.680 112.250 79.820 112.450 ;
        RECT 123.765 112.450 126.370 112.590 ;
        RECT 123.765 112.405 124.055 112.450 ;
        RECT 126.050 112.390 126.370 112.450 ;
        RECT 82.825 112.250 83.115 112.295 ;
        RECT 79.680 112.110 83.115 112.250 ;
        RECT 82.825 112.065 83.115 112.110 ;
        RECT 94.310 112.050 94.630 112.310 ;
        RECT 107.190 112.050 107.510 112.310 ;
        RECT 124.225 112.250 124.515 112.295 ;
        RECT 125.130 112.250 125.450 112.310 ;
        RECT 124.225 112.110 125.450 112.250 ;
        RECT 124.225 112.065 124.515 112.110 ;
        RECT 125.130 112.050 125.450 112.110 ;
        RECT 28.085 111.910 28.375 111.955 ;
        RECT 28.530 111.910 28.850 111.970 ;
        RECT 28.085 111.770 28.850 111.910 ;
        RECT 28.085 111.725 28.375 111.770 ;
        RECT 28.530 111.710 28.850 111.770 ;
        RECT 79.590 111.710 79.910 111.970 ;
        RECT 80.050 111.910 80.370 111.970 ;
        RECT 81.890 111.910 82.210 111.970 ;
        RECT 80.050 111.770 82.210 111.910 ;
        RECT 80.050 111.710 80.370 111.770 ;
        RECT 81.890 111.710 82.210 111.770 ;
        RECT 93.850 111.710 94.170 111.970 ;
        RECT 21.140 111.570 21.430 111.615 ;
        RECT 23.920 111.570 24.210 111.615 ;
        RECT 25.780 111.570 26.070 111.615 ;
        RECT 21.140 111.430 26.070 111.570 ;
        RECT 21.140 111.385 21.430 111.430 ;
        RECT 23.920 111.385 24.210 111.430 ;
        RECT 25.780 111.385 26.070 111.430 ;
        RECT 27.575 111.570 27.865 111.615 ;
        RECT 29.465 111.570 29.755 111.615 ;
        RECT 32.585 111.570 32.875 111.615 ;
        RECT 27.575 111.430 32.875 111.570 ;
        RECT 27.575 111.385 27.865 111.430 ;
        RECT 29.465 111.385 29.755 111.430 ;
        RECT 32.585 111.385 32.875 111.430 ;
        RECT 20.250 111.230 20.570 111.290 ;
        RECT 44.185 111.230 44.475 111.275 ;
        RECT 20.250 111.090 44.475 111.230 ;
        RECT 20.250 111.030 20.570 111.090 ;
        RECT 44.185 111.045 44.475 111.090 ;
        RECT 117.325 111.230 117.615 111.275 ;
        RECT 120.530 111.230 120.850 111.290 ;
        RECT 117.325 111.090 120.850 111.230 ;
        RECT 117.325 111.045 117.615 111.090 ;
        RECT 120.530 111.030 120.850 111.090 ;
        RECT 124.670 111.230 124.990 111.290 ;
        RECT 125.145 111.230 125.435 111.275 ;
        RECT 124.670 111.090 125.435 111.230 ;
        RECT 124.670 111.030 124.990 111.090 ;
        RECT 125.145 111.045 125.435 111.090 ;
        RECT 23.485 110.210 23.775 110.255 ;
        RECT 28.070 110.210 28.390 110.270 ;
        RECT 23.485 110.070 28.390 110.210 ;
        RECT 23.485 110.025 23.775 110.070 ;
        RECT 28.070 110.010 28.390 110.070 ;
        RECT 28.530 110.010 28.850 110.270 ;
        RECT 42.790 110.210 43.110 110.270 ;
        RECT 46.945 110.210 47.235 110.255 ;
        RECT 42.790 110.070 47.235 110.210 ;
        RECT 42.790 110.010 43.110 110.070 ;
        RECT 46.945 110.025 47.235 110.070 ;
        RECT 74.070 110.210 74.390 110.270 ;
        RECT 75.005 110.210 75.295 110.255 ;
        RECT 74.070 110.070 75.295 110.210 ;
        RECT 74.070 110.010 74.390 110.070 ;
        RECT 75.005 110.025 75.295 110.070 ;
        RECT 115.470 110.010 115.790 110.270 ;
        RECT 117.310 110.010 117.630 110.270 ;
        RECT 27.165 109.685 27.455 109.915 ;
        RECT 39.075 109.870 39.365 109.915 ;
        RECT 40.965 109.870 41.255 109.915 ;
        RECT 44.085 109.870 44.375 109.915 ;
        RECT 39.075 109.730 44.375 109.870 ;
        RECT 39.075 109.685 39.365 109.730 ;
        RECT 40.965 109.685 41.255 109.730 ;
        RECT 44.085 109.685 44.375 109.730 ;
        RECT 67.185 109.870 67.475 109.915 ;
        RECT 73.150 109.870 73.470 109.930 ;
        RECT 67.185 109.730 73.470 109.870 ;
        RECT 67.185 109.685 67.475 109.730 ;
        RECT 27.240 109.530 27.380 109.685 ;
        RECT 73.150 109.670 73.470 109.730 ;
        RECT 77.750 109.870 78.070 109.930 ;
        RECT 97.990 109.870 98.310 109.930 ;
        RECT 104.445 109.870 104.735 109.915 ;
        RECT 109.950 109.870 110.270 109.930 ;
        RECT 77.750 109.730 87.640 109.870 ;
        RECT 77.750 109.670 78.070 109.730 ;
        RECT 39.585 109.530 39.875 109.575 ;
        RECT 27.240 109.390 39.875 109.530 ;
        RECT 39.585 109.345 39.875 109.390 ;
        RECT 44.630 109.530 44.950 109.590 ;
        RECT 51.990 109.530 52.310 109.590 ;
        RECT 44.630 109.390 47.620 109.530 ;
        RECT 44.630 109.330 44.950 109.390 ;
        RECT 23.010 108.990 23.330 109.250 ;
        RECT 25.770 109.190 26.090 109.250 ;
        RECT 26.245 109.190 26.535 109.235 ;
        RECT 25.770 109.050 26.535 109.190 ;
        RECT 25.770 108.990 26.090 109.050 ;
        RECT 26.245 109.005 26.535 109.050 ;
        RECT 26.690 109.190 27.010 109.250 ;
        RECT 27.625 109.190 27.915 109.235 ;
        RECT 26.690 109.050 27.915 109.190 ;
        RECT 26.690 108.990 27.010 109.050 ;
        RECT 27.625 109.005 27.915 109.050 ;
        RECT 38.190 108.990 38.510 109.250 ;
        RECT 47.480 109.235 47.620 109.390 ;
        RECT 51.990 109.390 60.960 109.530 ;
        RECT 51.990 109.330 52.310 109.390 ;
        RECT 38.670 109.190 38.960 109.235 ;
        RECT 40.505 109.190 40.795 109.235 ;
        RECT 44.085 109.190 44.375 109.235 ;
        RECT 38.670 109.050 44.375 109.190 ;
        RECT 38.670 109.005 38.960 109.050 ;
        RECT 40.505 109.005 40.795 109.050 ;
        RECT 44.085 109.005 44.375 109.050 ;
        RECT 27.150 108.850 27.470 108.910 ;
        RECT 45.165 108.895 45.455 109.210 ;
        RECT 47.405 109.005 47.695 109.235 ;
        RECT 50.610 109.190 50.930 109.250 ;
        RECT 51.085 109.190 51.375 109.235 ;
        RECT 50.610 109.050 51.375 109.190 ;
        RECT 50.610 108.990 50.930 109.050 ;
        RECT 51.085 109.005 51.375 109.050 ;
        RECT 52.910 109.190 53.230 109.250 ;
        RECT 57.065 109.190 57.355 109.235 ;
        RECT 52.910 109.050 57.355 109.190 ;
        RECT 52.910 108.990 53.230 109.050 ;
        RECT 57.065 109.005 57.355 109.050 ;
        RECT 60.270 108.990 60.590 109.250 ;
        RECT 60.820 109.190 60.960 109.390 ;
        RECT 63.505 109.190 63.795 109.235 ;
        RECT 60.820 109.050 63.795 109.190 ;
        RECT 63.505 109.005 63.795 109.050 ;
        RECT 75.450 108.990 75.770 109.250 ;
        RECT 81.890 109.190 82.210 109.250 ;
        RECT 87.500 109.235 87.640 109.730 ;
        RECT 97.990 109.730 100.520 109.870 ;
        RECT 97.990 109.670 98.310 109.730 ;
        RECT 99.385 109.530 99.675 109.575 ;
        RECT 99.830 109.530 100.150 109.590 ;
        RECT 99.385 109.390 100.150 109.530 ;
        RECT 99.385 109.345 99.675 109.390 ;
        RECT 99.830 109.330 100.150 109.390 ;
        RECT 86.045 109.190 86.335 109.235 ;
        RECT 81.890 109.050 86.335 109.190 ;
        RECT 81.890 108.990 82.210 109.050 ;
        RECT 86.045 109.005 86.335 109.050 ;
        RECT 87.425 109.005 87.715 109.235 ;
        RECT 94.310 109.190 94.630 109.250 ;
        RECT 100.380 109.235 100.520 109.730 ;
        RECT 104.445 109.730 110.270 109.870 ;
        RECT 104.445 109.685 104.735 109.730 ;
        RECT 109.950 109.670 110.270 109.730 ;
        RECT 120.185 109.870 120.475 109.915 ;
        RECT 123.305 109.870 123.595 109.915 ;
        RECT 125.195 109.870 125.485 109.915 ;
        RECT 120.185 109.730 125.485 109.870 ;
        RECT 120.185 109.685 120.475 109.730 ;
        RECT 123.305 109.685 123.595 109.730 ;
        RECT 125.195 109.685 125.485 109.730 ;
        RECT 100.840 109.390 116.160 109.530 ;
        RECT 98.925 109.190 99.215 109.235 ;
        RECT 94.310 109.050 100.060 109.190 ;
        RECT 29.005 108.850 29.295 108.895 ;
        RECT 41.865 108.850 42.515 108.895 ;
        RECT 45.165 108.850 45.755 108.895 ;
        RECT 27.150 108.710 29.295 108.850 ;
        RECT 27.150 108.650 27.470 108.710 ;
        RECT 29.005 108.665 29.295 108.710 ;
        RECT 32.300 108.710 45.755 108.850 ;
        RECT 17.950 108.510 18.270 108.570 ;
        RECT 32.300 108.510 32.440 108.710 ;
        RECT 41.865 108.665 42.515 108.710 ;
        RECT 45.465 108.665 45.755 108.710 ;
        RECT 61.650 108.650 61.970 108.910 ;
        RECT 73.625 108.850 73.915 108.895 ;
        RECT 74.070 108.850 74.390 108.910 ;
        RECT 73.625 108.710 74.390 108.850 ;
        RECT 73.625 108.665 73.915 108.710 ;
        RECT 74.070 108.650 74.390 108.710 ;
        RECT 85.570 108.650 85.890 108.910 ;
        RECT 86.120 108.850 86.260 109.005 ;
        RECT 94.310 108.990 94.630 109.050 ;
        RECT 98.925 109.005 99.215 109.050 ;
        RECT 94.400 108.850 94.540 108.990 ;
        RECT 86.120 108.710 94.540 108.850 ;
        RECT 97.545 108.850 97.835 108.895 ;
        RECT 99.370 108.850 99.690 108.910 ;
        RECT 97.545 108.710 99.690 108.850 ;
        RECT 99.920 108.850 100.060 109.050 ;
        RECT 100.305 109.005 100.595 109.235 ;
        RECT 100.840 108.850 100.980 109.390 ;
        RECT 116.020 109.250 116.160 109.390 ;
        RECT 124.670 109.330 124.990 109.590 ;
        RECT 111.330 108.990 111.650 109.250 ;
        RECT 112.725 109.190 113.015 109.235 ;
        RECT 113.170 109.190 113.490 109.250 ;
        RECT 112.725 109.050 113.490 109.190 ;
        RECT 112.725 109.005 113.015 109.050 ;
        RECT 113.170 108.990 113.490 109.050 ;
        RECT 114.550 108.990 114.870 109.250 ;
        RECT 115.930 108.990 116.250 109.250 ;
        RECT 99.920 108.710 100.980 108.850 ;
        RECT 97.545 108.665 97.835 108.710 ;
        RECT 99.370 108.650 99.690 108.710 ;
        RECT 110.870 108.650 111.190 108.910 ;
        RECT 119.105 108.895 119.395 109.210 ;
        RECT 120.185 109.190 120.475 109.235 ;
        RECT 123.765 109.190 124.055 109.235 ;
        RECT 125.600 109.190 125.890 109.235 ;
        RECT 120.185 109.050 125.890 109.190 ;
        RECT 120.185 109.005 120.475 109.050 ;
        RECT 123.765 109.005 124.055 109.050 ;
        RECT 125.600 109.005 125.890 109.050 ;
        RECT 126.050 108.990 126.370 109.250 ;
        RECT 116.405 108.850 116.695 108.895 ;
        RECT 118.805 108.850 119.395 108.895 ;
        RECT 122.045 108.850 122.695 108.895 ;
        RECT 116.405 108.710 122.695 108.850 ;
        RECT 116.405 108.665 116.695 108.710 ;
        RECT 118.805 108.665 119.095 108.710 ;
        RECT 122.045 108.665 122.695 108.710 ;
        RECT 17.950 108.370 32.440 108.510 ;
        RECT 36.365 108.510 36.655 108.555 ;
        RECT 37.730 108.510 38.050 108.570 ;
        RECT 36.365 108.370 38.050 108.510 ;
        RECT 17.950 108.310 18.270 108.370 ;
        RECT 36.365 108.325 36.655 108.370 ;
        RECT 37.730 108.310 38.050 108.370 ;
        RECT 48.310 108.310 48.630 108.570 ;
        RECT 52.005 108.510 52.295 108.555 ;
        RECT 55.670 108.510 55.990 108.570 ;
        RECT 52.005 108.370 55.990 108.510 ;
        RECT 52.005 108.325 52.295 108.370 ;
        RECT 55.670 108.310 55.990 108.370 ;
        RECT 57.985 108.510 58.275 108.555 ;
        RECT 60.730 108.510 61.050 108.570 ;
        RECT 57.985 108.370 61.050 108.510 ;
        RECT 57.985 108.325 58.275 108.370 ;
        RECT 60.730 108.310 61.050 108.370 ;
        RECT 64.425 108.510 64.715 108.555 ;
        RECT 70.850 108.510 71.170 108.570 ;
        RECT 64.425 108.370 71.170 108.510 ;
        RECT 64.425 108.325 64.715 108.370 ;
        RECT 70.850 108.310 71.170 108.370 ;
        RECT 79.145 108.510 79.435 108.555 ;
        RECT 86.030 108.510 86.350 108.570 ;
        RECT 79.145 108.370 86.350 108.510 ;
        RECT 79.145 108.325 79.435 108.370 ;
        RECT 86.030 108.310 86.350 108.370 ;
        RECT 86.505 108.510 86.795 108.555 ;
        RECT 87.410 108.510 87.730 108.570 ;
        RECT 86.505 108.370 87.730 108.510 ;
        RECT 86.505 108.325 86.795 108.370 ;
        RECT 87.410 108.310 87.730 108.370 ;
        RECT 88.345 108.510 88.635 108.555 ;
        RECT 90.630 108.510 90.950 108.570 ;
        RECT 88.345 108.370 90.950 108.510 ;
        RECT 88.345 108.325 88.635 108.370 ;
        RECT 90.630 108.310 90.950 108.370 ;
        RECT 91.105 108.510 91.395 108.555 ;
        RECT 97.990 108.510 98.310 108.570 ;
        RECT 91.105 108.370 98.310 108.510 ;
        RECT 91.105 108.325 91.395 108.370 ;
        RECT 97.990 108.310 98.310 108.370 ;
        RECT 101.225 108.510 101.515 108.555 ;
        RECT 106.730 108.510 107.050 108.570 ;
        RECT 101.225 108.370 107.050 108.510 ;
        RECT 101.225 108.325 101.515 108.370 ;
        RECT 106.730 108.310 107.050 108.370 ;
        RECT 111.790 108.510 112.110 108.570 ;
        RECT 112.265 108.510 112.555 108.555 ;
        RECT 111.790 108.370 112.555 108.510 ;
        RECT 111.790 108.310 112.110 108.370 ;
        RECT 112.265 108.325 112.555 108.370 ;
        RECT 113.645 108.510 113.935 108.555 ;
        RECT 120.990 108.510 121.310 108.570 ;
        RECT 113.645 108.370 121.310 108.510 ;
        RECT 113.645 108.325 113.935 108.370 ;
        RECT 120.990 108.310 121.310 108.370 ;
        RECT 17.950 107.290 18.270 107.550 ;
        RECT 18.870 107.290 19.190 107.550 ;
        RECT 25.310 107.490 25.630 107.550 ;
        RECT 28.085 107.490 28.375 107.535 ;
        RECT 25.310 107.350 28.375 107.490 ;
        RECT 25.310 107.290 25.630 107.350 ;
        RECT 28.085 107.305 28.375 107.350 ;
        RECT 28.530 107.490 28.850 107.550 ;
        RECT 28.530 107.350 37.960 107.490 ;
        RECT 28.530 107.290 28.850 107.350 ;
        RECT 20.365 107.150 20.655 107.195 ;
        RECT 22.550 107.150 22.870 107.210 ;
        RECT 23.605 107.150 24.255 107.195 ;
        RECT 20.365 107.010 24.255 107.150 ;
        RECT 20.365 106.965 20.955 107.010 ;
        RECT 18.425 106.625 18.715 106.855 ;
        RECT 20.665 106.650 20.955 106.965 ;
        RECT 22.550 106.950 22.870 107.010 ;
        RECT 23.605 106.965 24.255 107.010 ;
        RECT 26.245 107.150 26.535 107.195 ;
        RECT 28.990 107.150 29.310 107.210 ;
        RECT 26.245 107.010 29.310 107.150 ;
        RECT 26.245 106.965 26.535 107.010 ;
        RECT 28.990 106.950 29.310 107.010 ;
        RECT 29.565 107.150 29.855 107.195 ;
        RECT 32.805 107.150 33.455 107.195 ;
        RECT 29.565 107.010 33.455 107.150 ;
        RECT 29.565 106.965 30.155 107.010 ;
        RECT 32.805 106.965 33.455 107.010 ;
        RECT 34.050 107.150 34.370 107.210 ;
        RECT 35.445 107.150 35.735 107.195 ;
        RECT 34.050 107.010 35.735 107.150 ;
        RECT 21.745 106.810 22.035 106.855 ;
        RECT 25.325 106.810 25.615 106.855 ;
        RECT 27.160 106.810 27.450 106.855 ;
        RECT 21.745 106.670 27.450 106.810 ;
        RECT 21.745 106.625 22.035 106.670 ;
        RECT 25.325 106.625 25.615 106.670 ;
        RECT 27.160 106.625 27.450 106.670 ;
        RECT 28.070 106.810 28.390 106.870 ;
        RECT 29.865 106.810 30.155 106.965 ;
        RECT 34.050 106.950 34.370 107.010 ;
        RECT 35.445 106.965 35.735 107.010 ;
        RECT 37.820 106.855 37.960 107.350 ;
        RECT 48.325 107.305 48.615 107.535 ;
        RECT 47.865 107.150 48.155 107.195 ;
        RECT 48.400 107.150 48.540 107.305 ;
        RECT 61.650 107.290 61.970 107.550 ;
        RECT 86.965 107.490 87.255 107.535 ;
        RECT 85.200 107.350 87.255 107.490 ;
        RECT 47.865 107.010 48.540 107.150 ;
        RECT 49.805 107.150 50.095 107.195 ;
        RECT 53.045 107.150 53.695 107.195 ;
        RECT 49.805 107.010 53.695 107.150 ;
        RECT 47.865 106.965 48.155 107.010 ;
        RECT 49.805 106.965 50.395 107.010 ;
        RECT 53.045 106.965 53.695 107.010 ;
        RECT 50.105 106.870 50.395 106.965 ;
        RECT 55.670 106.950 55.990 107.210 ;
        RECT 61.740 107.150 61.880 107.290 ;
        RECT 85.200 107.195 85.340 107.350 ;
        RECT 86.965 107.305 87.255 107.350 ;
        RECT 99.370 107.290 99.690 107.550 ;
        RECT 115.930 107.490 116.250 107.550 ;
        RECT 124.210 107.490 124.530 107.550 ;
        RECT 124.685 107.490 124.975 107.535 ;
        RECT 113.260 107.350 123.060 107.490 ;
        RECT 63.965 107.150 64.255 107.195 ;
        RECT 66.365 107.150 66.655 107.195 ;
        RECT 69.605 107.150 70.255 107.195 ;
        RECT 60.360 107.010 63.720 107.150 ;
        RECT 28.070 106.670 30.155 106.810 ;
        RECT 18.500 106.470 18.640 106.625 ;
        RECT 28.070 106.610 28.390 106.670 ;
        RECT 29.865 106.650 30.155 106.670 ;
        RECT 30.945 106.810 31.235 106.855 ;
        RECT 34.525 106.810 34.815 106.855 ;
        RECT 36.360 106.810 36.650 106.855 ;
        RECT 30.945 106.670 36.650 106.810 ;
        RECT 30.945 106.625 31.235 106.670 ;
        RECT 34.525 106.625 34.815 106.670 ;
        RECT 36.360 106.625 36.650 106.670 ;
        RECT 37.745 106.810 38.035 106.855 ;
        RECT 39.570 106.810 39.890 106.870 ;
        RECT 37.745 106.670 39.890 106.810 ;
        RECT 37.745 106.625 38.035 106.670 ;
        RECT 39.570 106.610 39.890 106.670 ;
        RECT 40.045 106.810 40.335 106.855 ;
        RECT 48.770 106.810 49.090 106.870 ;
        RECT 40.045 106.670 49.090 106.810 ;
        RECT 40.045 106.625 40.335 106.670 ;
        RECT 48.770 106.610 49.090 106.670 ;
        RECT 50.105 106.650 50.470 106.870 ;
        RECT 50.150 106.610 50.470 106.650 ;
        RECT 51.185 106.810 51.475 106.855 ;
        RECT 54.765 106.810 55.055 106.855 ;
        RECT 56.600 106.810 56.890 106.855 ;
        RECT 51.185 106.670 56.890 106.810 ;
        RECT 51.185 106.625 51.475 106.670 ;
        RECT 54.765 106.625 55.055 106.670 ;
        RECT 56.600 106.625 56.890 106.670 ;
        RECT 57.050 106.610 57.370 106.870 ;
        RECT 60.360 106.855 60.500 107.010 ;
        RECT 58.445 106.810 58.735 106.855 ;
        RECT 60.285 106.810 60.575 106.855 ;
        RECT 58.445 106.670 60.575 106.810 ;
        RECT 58.445 106.625 58.735 106.670 ;
        RECT 60.285 106.625 60.575 106.670 ;
        RECT 61.190 106.810 61.510 106.870 ;
        RECT 63.580 106.855 63.720 107.010 ;
        RECT 63.965 107.010 70.255 107.150 ;
        RECT 63.965 106.965 64.255 107.010 ;
        RECT 66.365 106.965 66.955 107.010 ;
        RECT 69.605 106.965 70.255 107.010 ;
        RECT 79.245 107.150 79.535 107.195 ;
        RECT 82.485 107.150 83.135 107.195 ;
        RECT 79.245 107.010 83.135 107.150 ;
        RECT 79.245 106.965 79.835 107.010 ;
        RECT 82.485 106.965 83.135 107.010 ;
        RECT 85.125 106.965 85.415 107.195 ;
        RECT 91.665 107.150 91.955 107.195 ;
        RECT 93.850 107.150 94.170 107.210 ;
        RECT 94.905 107.150 95.555 107.195 ;
        RECT 91.665 107.010 95.555 107.150 ;
        RECT 91.665 106.965 92.255 107.010 ;
        RECT 61.665 106.810 61.955 106.855 ;
        RECT 61.190 106.670 61.955 106.810 ;
        RECT 23.010 106.470 23.330 106.530 ;
        RECT 18.500 106.330 23.330 106.470 ;
        RECT 23.010 106.270 23.330 106.330 ;
        RECT 27.610 106.470 27.930 106.530 ;
        RECT 36.825 106.470 37.115 106.515 ;
        RECT 38.190 106.470 38.510 106.530 ;
        RECT 40.490 106.470 40.810 106.530 ;
        RECT 58.520 106.470 58.660 106.625 ;
        RECT 61.190 106.610 61.510 106.670 ;
        RECT 61.665 106.625 61.955 106.670 ;
        RECT 63.505 106.625 63.795 106.855 ;
        RECT 66.665 106.650 66.955 106.965 ;
        RECT 79.545 106.870 79.835 106.965 ;
        RECT 67.745 106.810 68.035 106.855 ;
        RECT 71.325 106.810 71.615 106.855 ;
        RECT 73.160 106.810 73.450 106.855 ;
        RECT 67.745 106.670 73.450 106.810 ;
        RECT 67.745 106.625 68.035 106.670 ;
        RECT 71.325 106.625 71.615 106.670 ;
        RECT 73.160 106.625 73.450 106.670 ;
        RECT 73.610 106.610 73.930 106.870 ;
        RECT 75.925 106.625 76.215 106.855 ;
        RECT 72.245 106.470 72.535 106.515 ;
        RECT 27.610 106.330 40.810 106.470 ;
        RECT 27.610 106.270 27.930 106.330 ;
        RECT 36.825 106.285 37.115 106.330 ;
        RECT 38.190 106.270 38.510 106.330 ;
        RECT 40.490 106.270 40.810 106.330 ;
        RECT 50.700 106.330 58.660 106.470 ;
        RECT 62.660 106.330 72.535 106.470 ;
        RECT 76.000 106.470 76.140 106.625 ;
        RECT 76.370 106.610 76.690 106.870 ;
        RECT 79.545 106.650 79.910 106.870 ;
        RECT 79.590 106.610 79.910 106.650 ;
        RECT 80.625 106.810 80.915 106.855 ;
        RECT 84.205 106.810 84.495 106.855 ;
        RECT 86.040 106.810 86.330 106.855 ;
        RECT 80.625 106.670 86.330 106.810 ;
        RECT 80.625 106.625 80.915 106.670 ;
        RECT 84.205 106.625 84.495 106.670 ;
        RECT 86.040 106.625 86.330 106.670 ;
        RECT 86.950 106.810 87.270 106.870 ;
        RECT 87.885 106.810 88.175 106.855 ;
        RECT 86.950 106.670 88.175 106.810 ;
        RECT 86.950 106.610 87.270 106.670 ;
        RECT 87.885 106.625 88.175 106.670 ;
        RECT 91.965 106.650 92.255 106.965 ;
        RECT 93.850 106.950 94.170 107.010 ;
        RECT 94.905 106.965 95.555 107.010 ;
        RECT 99.830 107.150 100.150 107.210 ;
        RECT 100.865 107.150 101.155 107.195 ;
        RECT 104.105 107.150 104.755 107.195 ;
        RECT 99.830 107.010 104.755 107.150 ;
        RECT 99.830 106.950 100.150 107.010 ;
        RECT 100.865 106.965 101.455 107.010 ;
        RECT 104.105 106.965 104.755 107.010 ;
        RECT 93.045 106.810 93.335 106.855 ;
        RECT 96.625 106.810 96.915 106.855 ;
        RECT 98.460 106.810 98.750 106.855 ;
        RECT 93.045 106.670 98.750 106.810 ;
        RECT 93.045 106.625 93.335 106.670 ;
        RECT 96.625 106.625 96.915 106.670 ;
        RECT 98.460 106.625 98.750 106.670 ;
        RECT 101.165 106.650 101.455 106.965 ;
        RECT 106.730 106.950 107.050 107.210 ;
        RECT 113.260 106.855 113.400 107.350 ;
        RECT 115.930 107.290 116.250 107.350 ;
        RECT 113.645 107.150 113.935 107.195 ;
        RECT 116.505 107.150 116.795 107.195 ;
        RECT 119.745 107.150 120.395 107.195 ;
        RECT 113.645 107.010 120.395 107.150 ;
        RECT 113.645 106.965 113.935 107.010 ;
        RECT 116.505 106.965 117.095 107.010 ;
        RECT 119.745 106.965 120.395 107.010 ;
        RECT 120.990 107.150 121.310 107.210 ;
        RECT 122.385 107.150 122.675 107.195 ;
        RECT 120.990 107.010 122.675 107.150 ;
        RECT 122.920 107.150 123.060 107.350 ;
        RECT 124.210 107.350 124.975 107.490 ;
        RECT 124.210 107.290 124.530 107.350 ;
        RECT 124.685 107.305 124.975 107.350 ;
        RECT 122.920 107.010 124.440 107.150 ;
        RECT 102.245 106.810 102.535 106.855 ;
        RECT 105.825 106.810 106.115 106.855 ;
        RECT 107.660 106.810 107.950 106.855 ;
        RECT 102.245 106.670 107.950 106.810 ;
        RECT 102.245 106.625 102.535 106.670 ;
        RECT 105.825 106.625 106.115 106.670 ;
        RECT 107.660 106.625 107.950 106.670 ;
        RECT 109.505 106.810 109.795 106.855 ;
        RECT 109.965 106.810 110.255 106.855 ;
        RECT 113.185 106.810 113.475 106.855 ;
        RECT 109.505 106.670 113.475 106.810 ;
        RECT 109.505 106.625 109.795 106.670 ;
        RECT 109.965 106.625 110.255 106.670 ;
        RECT 113.185 106.625 113.475 106.670 ;
        RECT 116.805 106.650 117.095 106.965 ;
        RECT 120.990 106.950 121.310 107.010 ;
        RECT 122.385 106.965 122.675 107.010 ;
        RECT 124.300 106.855 124.440 107.010 ;
        RECT 117.885 106.810 118.175 106.855 ;
        RECT 121.465 106.810 121.755 106.855 ;
        RECT 123.300 106.810 123.590 106.855 ;
        RECT 117.885 106.670 123.590 106.810 ;
        RECT 117.885 106.625 118.175 106.670 ;
        RECT 121.465 106.625 121.755 106.670 ;
        RECT 123.300 106.625 123.590 106.670 ;
        RECT 124.225 106.625 124.515 106.855 ;
        RECT 81.890 106.470 82.210 106.530 ;
        RECT 76.000 106.330 82.210 106.470 ;
        RECT 50.700 106.190 50.840 106.330 ;
        RECT 21.745 106.130 22.035 106.175 ;
        RECT 24.865 106.130 25.155 106.175 ;
        RECT 26.755 106.130 27.045 106.175 ;
        RECT 21.745 105.990 27.045 106.130 ;
        RECT 21.745 105.945 22.035 105.990 ;
        RECT 24.865 105.945 25.155 105.990 ;
        RECT 26.755 105.945 27.045 105.990 ;
        RECT 30.945 106.130 31.235 106.175 ;
        RECT 34.065 106.130 34.355 106.175 ;
        RECT 35.955 106.130 36.245 106.175 ;
        RECT 30.945 105.990 36.245 106.130 ;
        RECT 30.945 105.945 31.235 105.990 ;
        RECT 34.065 105.945 34.355 105.990 ;
        RECT 35.955 105.945 36.245 105.990 ;
        RECT 39.570 106.130 39.890 106.190 ;
        RECT 50.610 106.130 50.930 106.190 ;
        RECT 62.660 106.175 62.800 106.330 ;
        RECT 72.245 106.285 72.535 106.330 ;
        RECT 81.890 106.270 82.210 106.330 ;
        RECT 85.110 106.470 85.430 106.530 ;
        RECT 86.505 106.470 86.795 106.515 ;
        RECT 85.110 106.330 86.795 106.470 ;
        RECT 85.110 106.270 85.430 106.330 ;
        RECT 86.505 106.285 86.795 106.330 ;
        RECT 97.530 106.270 97.850 106.530 ;
        RECT 98.910 106.270 99.230 106.530 ;
        RECT 106.730 106.470 107.050 106.530 ;
        RECT 108.125 106.470 108.415 106.515 ;
        RECT 112.250 106.470 112.570 106.530 ;
        RECT 120.070 106.470 120.390 106.530 ;
        RECT 123.765 106.470 124.055 106.515 ;
        RECT 126.050 106.470 126.370 106.530 ;
        RECT 106.730 106.330 126.370 106.470 ;
        RECT 106.730 106.270 107.050 106.330 ;
        RECT 108.125 106.285 108.415 106.330 ;
        RECT 112.250 106.270 112.570 106.330 ;
        RECT 120.070 106.270 120.390 106.330 ;
        RECT 123.765 106.285 124.055 106.330 ;
        RECT 126.050 106.270 126.370 106.330 ;
        RECT 39.570 105.990 50.930 106.130 ;
        RECT 39.570 105.930 39.890 105.990 ;
        RECT 50.610 105.930 50.930 105.990 ;
        RECT 51.185 106.130 51.475 106.175 ;
        RECT 54.305 106.130 54.595 106.175 ;
        RECT 56.195 106.130 56.485 106.175 ;
        RECT 51.185 105.990 56.485 106.130 ;
        RECT 51.185 105.945 51.475 105.990 ;
        RECT 54.305 105.945 54.595 105.990 ;
        RECT 56.195 105.945 56.485 105.990 ;
        RECT 62.585 105.945 62.875 106.175 ;
        RECT 64.410 106.130 64.730 106.190 ;
        RECT 63.120 105.990 64.730 106.130 ;
        RECT 38.205 105.790 38.495 105.835 ;
        RECT 41.410 105.790 41.730 105.850 ;
        RECT 38.205 105.650 41.730 105.790 ;
        RECT 38.205 105.605 38.495 105.650 ;
        RECT 41.410 105.590 41.730 105.650 ;
        RECT 56.590 105.790 56.910 105.850 ;
        RECT 57.985 105.790 58.275 105.835 ;
        RECT 56.590 105.650 58.275 105.790 ;
        RECT 56.590 105.590 56.910 105.650 ;
        RECT 57.985 105.605 58.275 105.650 ;
        RECT 60.745 105.790 61.035 105.835 ;
        RECT 63.120 105.790 63.260 105.990 ;
        RECT 64.410 105.930 64.730 105.990 ;
        RECT 67.745 106.130 68.035 106.175 ;
        RECT 70.865 106.130 71.155 106.175 ;
        RECT 72.755 106.130 73.045 106.175 ;
        RECT 67.745 105.990 73.045 106.130 ;
        RECT 67.745 105.945 68.035 105.990 ;
        RECT 70.865 105.945 71.155 105.990 ;
        RECT 72.755 105.945 73.045 105.990 ;
        RECT 75.465 106.130 75.755 106.175 ;
        RECT 78.210 106.130 78.530 106.190 ;
        RECT 75.465 105.990 78.530 106.130 ;
        RECT 75.465 105.945 75.755 105.990 ;
        RECT 78.210 105.930 78.530 105.990 ;
        RECT 80.625 106.130 80.915 106.175 ;
        RECT 83.745 106.130 84.035 106.175 ;
        RECT 85.635 106.130 85.925 106.175 ;
        RECT 80.625 105.990 85.925 106.130 ;
        RECT 80.625 105.945 80.915 105.990 ;
        RECT 83.745 105.945 84.035 105.990 ;
        RECT 85.635 105.945 85.925 105.990 ;
        RECT 93.045 106.130 93.335 106.175 ;
        RECT 96.165 106.130 96.455 106.175 ;
        RECT 98.055 106.130 98.345 106.175 ;
        RECT 93.045 105.990 98.345 106.130 ;
        RECT 93.045 105.945 93.335 105.990 ;
        RECT 96.165 105.945 96.455 105.990 ;
        RECT 98.055 105.945 98.345 105.990 ;
        RECT 102.245 106.130 102.535 106.175 ;
        RECT 105.365 106.130 105.655 106.175 ;
        RECT 107.255 106.130 107.545 106.175 ;
        RECT 102.245 105.990 107.545 106.130 ;
        RECT 102.245 105.945 102.535 105.990 ;
        RECT 105.365 105.945 105.655 105.990 ;
        RECT 107.255 105.945 107.545 105.990 ;
        RECT 117.885 106.130 118.175 106.175 ;
        RECT 121.005 106.130 121.295 106.175 ;
        RECT 122.895 106.130 123.185 106.175 ;
        RECT 117.885 105.990 123.185 106.130 ;
        RECT 117.885 105.945 118.175 105.990 ;
        RECT 121.005 105.945 121.295 105.990 ;
        RECT 122.895 105.945 123.185 105.990 ;
        RECT 60.745 105.650 63.260 105.790 ;
        RECT 63.950 105.790 64.270 105.850 ;
        RECT 64.885 105.790 65.175 105.835 ;
        RECT 63.950 105.650 65.175 105.790 ;
        RECT 60.745 105.605 61.035 105.650 ;
        RECT 63.950 105.590 64.270 105.650 ;
        RECT 64.885 105.605 65.175 105.650 ;
        RECT 77.290 105.590 77.610 105.850 ;
        RECT 77.750 105.590 78.070 105.850 ;
        RECT 90.170 105.590 90.490 105.850 ;
        RECT 109.030 105.590 109.350 105.850 ;
        RECT 110.410 105.590 110.730 105.850 ;
        RECT 115.010 105.590 115.330 105.850 ;
        RECT 22.550 104.770 22.870 104.830 ;
        RECT 26.705 104.770 26.995 104.815 ;
        RECT 22.550 104.630 26.995 104.770 ;
        RECT 22.550 104.570 22.870 104.630 ;
        RECT 26.705 104.585 26.995 104.630 ;
        RECT 28.070 104.570 28.390 104.830 ;
        RECT 28.990 104.570 29.310 104.830 ;
        RECT 50.150 104.770 50.470 104.830 ;
        RECT 52.005 104.770 52.295 104.815 ;
        RECT 50.150 104.630 52.295 104.770 ;
        RECT 50.150 104.570 50.470 104.630 ;
        RECT 52.005 104.585 52.295 104.630 ;
        RECT 74.070 104.770 74.390 104.830 ;
        RECT 76.385 104.770 76.675 104.815 ;
        RECT 74.070 104.630 76.675 104.770 ;
        RECT 74.070 104.570 74.390 104.630 ;
        RECT 76.385 104.585 76.675 104.630 ;
        RECT 85.570 104.570 85.890 104.830 ;
        RECT 95.705 104.770 95.995 104.815 ;
        RECT 97.530 104.770 97.850 104.830 ;
        RECT 106.730 104.770 107.050 104.830 ;
        RECT 87.960 104.630 94.540 104.770 ;
        RECT 27.150 104.230 27.470 104.490 ;
        RECT 31.305 104.430 31.595 104.475 ;
        RECT 34.050 104.430 34.370 104.490 ;
        RECT 31.305 104.290 34.370 104.430 ;
        RECT 31.305 104.245 31.595 104.290 ;
        RECT 34.050 104.230 34.370 104.290 ;
        RECT 34.625 104.430 34.915 104.475 ;
        RECT 37.745 104.430 38.035 104.475 ;
        RECT 39.635 104.430 39.925 104.475 ;
        RECT 34.625 104.290 39.925 104.430 ;
        RECT 34.625 104.245 34.915 104.290 ;
        RECT 37.745 104.245 38.035 104.290 ;
        RECT 39.635 104.245 39.925 104.290 ;
        RECT 43.825 104.430 44.115 104.475 ;
        RECT 46.945 104.430 47.235 104.475 ;
        RECT 48.835 104.430 49.125 104.475 ;
        RECT 43.825 104.290 49.125 104.430 ;
        RECT 43.825 104.245 44.115 104.290 ;
        RECT 46.945 104.245 47.235 104.290 ;
        RECT 48.835 104.245 49.125 104.290 ;
        RECT 57.165 104.430 57.455 104.475 ;
        RECT 60.285 104.430 60.575 104.475 ;
        RECT 62.175 104.430 62.465 104.475 ;
        RECT 57.165 104.290 62.465 104.430 ;
        RECT 57.165 104.245 57.455 104.290 ;
        RECT 60.285 104.245 60.575 104.290 ;
        RECT 62.175 104.245 62.465 104.290 ;
        RECT 66.365 104.430 66.655 104.475 ;
        RECT 69.485 104.430 69.775 104.475 ;
        RECT 71.375 104.430 71.665 104.475 ;
        RECT 66.365 104.290 71.665 104.430 ;
        RECT 66.365 104.245 66.655 104.290 ;
        RECT 69.485 104.245 69.775 104.290 ;
        RECT 71.375 104.245 71.665 104.290 ;
        RECT 79.245 104.430 79.535 104.475 ;
        RECT 82.365 104.430 82.655 104.475 ;
        RECT 84.255 104.430 84.545 104.475 ;
        RECT 87.960 104.430 88.100 104.630 ;
        RECT 79.245 104.290 84.545 104.430 ;
        RECT 79.245 104.245 79.535 104.290 ;
        RECT 82.365 104.245 82.655 104.290 ;
        RECT 84.255 104.245 84.545 104.290 ;
        RECT 85.200 104.290 88.100 104.430 ;
        RECT 88.445 104.430 88.735 104.475 ;
        RECT 91.565 104.430 91.855 104.475 ;
        RECT 93.455 104.430 93.745 104.475 ;
        RECT 88.445 104.290 93.745 104.430 ;
        RECT 27.240 104.090 27.380 104.230 ;
        RECT 85.200 104.150 85.340 104.290 ;
        RECT 88.445 104.245 88.735 104.290 ;
        RECT 91.565 104.245 91.855 104.290 ;
        RECT 93.455 104.245 93.745 104.290 ;
        RECT 94.400 104.430 94.540 104.630 ;
        RECT 95.705 104.630 97.850 104.770 ;
        RECT 95.705 104.585 95.995 104.630 ;
        RECT 97.530 104.570 97.850 104.630 ;
        RECT 102.220 104.630 107.050 104.770 ;
        RECT 98.910 104.430 99.230 104.490 ;
        RECT 94.400 104.290 99.230 104.430 ;
        RECT 31.765 104.090 32.055 104.135 ;
        RECT 27.240 103.950 32.055 104.090 ;
        RECT 31.765 103.905 32.055 103.950 ;
        RECT 40.950 103.890 41.270 104.150 ;
        RECT 48.310 103.890 48.630 104.150 ;
        RECT 61.190 104.090 61.510 104.150 ;
        RECT 61.665 104.090 61.955 104.135 ;
        RECT 61.190 103.950 61.955 104.090 ;
        RECT 61.190 103.890 61.510 103.950 ;
        RECT 61.665 103.905 61.955 103.950 ;
        RECT 63.045 104.090 63.335 104.135 ;
        RECT 72.245 104.090 72.535 104.135 ;
        RECT 73.610 104.090 73.930 104.150 ;
        RECT 63.045 103.950 73.930 104.090 ;
        RECT 63.045 103.905 63.335 103.950 ;
        RECT 72.245 103.905 72.535 103.950 ;
        RECT 73.610 103.890 73.930 103.950 ;
        RECT 77.290 104.090 77.610 104.150 ;
        RECT 83.745 104.090 84.035 104.135 ;
        RECT 77.290 103.950 84.035 104.090 ;
        RECT 77.290 103.890 77.610 103.950 ;
        RECT 83.745 103.905 84.035 103.950 ;
        RECT 85.110 103.890 85.430 104.150 ;
        RECT 90.630 104.090 90.950 104.150 ;
        RECT 94.400 104.135 94.540 104.290 ;
        RECT 98.910 104.230 99.230 104.290 ;
        RECT 102.220 104.135 102.360 104.630 ;
        RECT 106.730 104.570 107.050 104.630 ;
        RECT 110.870 104.770 111.190 104.830 ;
        RECT 111.345 104.770 111.635 104.815 ;
        RECT 110.870 104.630 111.635 104.770 ;
        RECT 110.870 104.570 111.190 104.630 ;
        RECT 111.345 104.585 111.635 104.630 ;
        RECT 103.015 104.430 103.305 104.475 ;
        RECT 104.905 104.430 105.195 104.475 ;
        RECT 108.025 104.430 108.315 104.475 ;
        RECT 103.015 104.290 108.315 104.430 ;
        RECT 103.015 104.245 103.305 104.290 ;
        RECT 104.905 104.245 105.195 104.290 ;
        RECT 108.025 104.245 108.315 104.290 ;
        RECT 114.205 104.430 114.495 104.475 ;
        RECT 117.325 104.430 117.615 104.475 ;
        RECT 119.215 104.430 119.505 104.475 ;
        RECT 114.205 104.290 119.505 104.430 ;
        RECT 114.205 104.245 114.495 104.290 ;
        RECT 117.325 104.245 117.615 104.290 ;
        RECT 119.215 104.245 119.505 104.290 ;
        RECT 92.945 104.090 93.235 104.135 ;
        RECT 90.630 103.950 93.235 104.090 ;
        RECT 90.630 103.890 90.950 103.950 ;
        RECT 92.945 103.905 93.235 103.950 ;
        RECT 94.325 103.905 94.615 104.135 ;
        RECT 102.145 103.905 102.435 104.135 ;
        RECT 103.525 104.090 103.815 104.135 ;
        RECT 106.270 104.090 106.590 104.150 ;
        RECT 103.525 103.950 106.590 104.090 ;
        RECT 103.525 103.905 103.815 103.950 ;
        RECT 106.270 103.890 106.590 103.950 ;
        RECT 111.790 104.090 112.110 104.150 ;
        RECT 118.705 104.090 118.995 104.135 ;
        RECT 111.790 103.950 118.995 104.090 ;
        RECT 111.790 103.890 112.110 103.950 ;
        RECT 118.705 103.905 118.995 103.950 ;
        RECT 120.070 103.890 120.390 104.150 ;
        RECT 23.010 103.750 23.330 103.810 ;
        RECT 27.165 103.750 27.455 103.795 ;
        RECT 27.625 103.750 27.915 103.795 ;
        RECT 28.530 103.750 28.850 103.810 ;
        RECT 23.010 103.610 28.850 103.750 ;
        RECT 23.010 103.550 23.330 103.610 ;
        RECT 27.165 103.565 27.455 103.610 ;
        RECT 27.625 103.565 27.915 103.610 ;
        RECT 28.530 103.550 28.850 103.610 ;
        RECT 29.925 103.565 30.215 103.795 ;
        RECT 30.385 103.750 30.675 103.795 ;
        RECT 30.830 103.750 31.150 103.810 ;
        RECT 30.385 103.610 31.150 103.750 ;
        RECT 30.385 103.565 30.675 103.610 ;
        RECT 30.000 103.070 30.140 103.565 ;
        RECT 30.830 103.550 31.150 103.610 ;
        RECT 33.545 103.455 33.835 103.770 ;
        RECT 34.625 103.750 34.915 103.795 ;
        RECT 38.205 103.750 38.495 103.795 ;
        RECT 40.040 103.750 40.330 103.795 ;
        RECT 34.625 103.610 40.330 103.750 ;
        RECT 34.625 103.565 34.915 103.610 ;
        RECT 38.205 103.565 38.495 103.610 ;
        RECT 40.040 103.565 40.330 103.610 ;
        RECT 40.490 103.550 40.810 103.810 ;
        RECT 33.245 103.410 33.835 103.455 ;
        RECT 36.485 103.410 37.135 103.455 ;
        RECT 38.650 103.410 38.970 103.470 ;
        RECT 33.245 103.270 38.970 103.410 ;
        RECT 33.245 103.225 33.535 103.270 ;
        RECT 36.485 103.225 37.135 103.270 ;
        RECT 38.650 103.210 38.970 103.270 ;
        RECT 39.110 103.210 39.430 103.470 ;
        RECT 35.430 103.070 35.750 103.130 ;
        RECT 30.000 102.930 35.750 103.070 ;
        RECT 40.580 103.070 40.720 103.550 ;
        RECT 41.410 103.410 41.730 103.470 ;
        RECT 42.745 103.455 43.035 103.770 ;
        RECT 43.825 103.750 44.115 103.795 ;
        RECT 47.405 103.750 47.695 103.795 ;
        RECT 49.240 103.750 49.530 103.795 ;
        RECT 43.825 103.610 49.530 103.750 ;
        RECT 43.825 103.565 44.115 103.610 ;
        RECT 47.405 103.565 47.695 103.610 ;
        RECT 49.240 103.565 49.530 103.610 ;
        RECT 49.705 103.565 49.995 103.795 ;
        RECT 50.610 103.750 50.930 103.810 ;
        RECT 52.465 103.750 52.755 103.795 ;
        RECT 50.610 103.610 52.755 103.750 ;
        RECT 42.445 103.410 43.035 103.455 ;
        RECT 45.685 103.410 46.335 103.455 ;
        RECT 41.410 103.270 46.335 103.410 ;
        RECT 41.410 103.210 41.730 103.270 ;
        RECT 42.445 103.225 42.735 103.270 ;
        RECT 45.685 103.225 46.335 103.270 ;
        RECT 49.780 103.070 49.920 103.565 ;
        RECT 50.610 103.550 50.930 103.610 ;
        RECT 52.465 103.565 52.755 103.610 ;
        RECT 56.085 103.455 56.375 103.770 ;
        RECT 57.165 103.750 57.455 103.795 ;
        RECT 60.745 103.750 61.035 103.795 ;
        RECT 62.580 103.750 62.870 103.795 ;
        RECT 57.165 103.610 62.870 103.750 ;
        RECT 57.165 103.565 57.455 103.610 ;
        RECT 60.745 103.565 61.035 103.610 ;
        RECT 62.580 103.565 62.870 103.610 ;
        RECT 55.785 103.410 56.375 103.455 ;
        RECT 56.590 103.410 56.910 103.470 ;
        RECT 59.025 103.410 59.675 103.455 ;
        RECT 55.785 103.270 59.675 103.410 ;
        RECT 55.785 103.225 56.075 103.270 ;
        RECT 56.590 103.210 56.910 103.270 ;
        RECT 59.025 103.225 59.675 103.270 ;
        RECT 64.410 103.410 64.730 103.470 ;
        RECT 65.285 103.455 65.575 103.770 ;
        RECT 66.365 103.750 66.655 103.795 ;
        RECT 69.945 103.750 70.235 103.795 ;
        RECT 71.780 103.750 72.070 103.795 ;
        RECT 78.210 103.770 78.530 103.810 ;
        RECT 66.365 103.610 72.070 103.750 ;
        RECT 66.365 103.565 66.655 103.610 ;
        RECT 69.945 103.565 70.235 103.610 ;
        RECT 71.780 103.565 72.070 103.610 ;
        RECT 78.165 103.550 78.530 103.770 ;
        RECT 79.245 103.750 79.535 103.795 ;
        RECT 82.825 103.750 83.115 103.795 ;
        RECT 84.660 103.750 84.950 103.795 ;
        RECT 87.410 103.770 87.730 103.810 ;
        RECT 79.245 103.610 84.950 103.750 ;
        RECT 79.245 103.565 79.535 103.610 ;
        RECT 82.825 103.565 83.115 103.610 ;
        RECT 84.660 103.565 84.950 103.610 ;
        RECT 87.365 103.550 87.730 103.770 ;
        RECT 88.445 103.750 88.735 103.795 ;
        RECT 92.025 103.750 92.315 103.795 ;
        RECT 93.860 103.750 94.150 103.795 ;
        RECT 88.445 103.610 94.150 103.750 ;
        RECT 88.445 103.565 88.735 103.610 ;
        RECT 92.025 103.565 92.315 103.610 ;
        RECT 93.860 103.565 94.150 103.610 ;
        RECT 94.785 103.565 95.075 103.795 ;
        RECT 102.610 103.750 102.900 103.795 ;
        RECT 104.445 103.750 104.735 103.795 ;
        RECT 108.025 103.750 108.315 103.795 ;
        RECT 102.610 103.610 108.315 103.750 ;
        RECT 102.610 103.565 102.900 103.610 ;
        RECT 104.445 103.565 104.735 103.610 ;
        RECT 108.025 103.565 108.315 103.610 ;
        RECT 109.030 103.770 109.350 103.810 ;
        RECT 64.985 103.410 65.575 103.455 ;
        RECT 68.225 103.410 68.875 103.455 ;
        RECT 64.410 103.270 68.875 103.410 ;
        RECT 64.410 103.210 64.730 103.270 ;
        RECT 64.985 103.225 65.275 103.270 ;
        RECT 68.225 103.225 68.875 103.270 ;
        RECT 70.850 103.210 71.170 103.470 ;
        RECT 78.165 103.455 78.455 103.550 ;
        RECT 87.365 103.455 87.655 103.550 ;
        RECT 77.865 103.410 78.455 103.455 ;
        RECT 81.105 103.410 81.755 103.455 ;
        RECT 77.865 103.270 81.755 103.410 ;
        RECT 77.865 103.225 78.155 103.270 ;
        RECT 81.105 103.225 81.755 103.270 ;
        RECT 87.065 103.410 87.655 103.455 ;
        RECT 90.305 103.410 90.955 103.455 ;
        RECT 87.065 103.270 90.955 103.410 ;
        RECT 87.065 103.225 87.355 103.270 ;
        RECT 90.305 103.225 90.955 103.270 ;
        RECT 40.580 102.930 49.920 103.070 ;
        RECT 35.430 102.870 35.750 102.930 ;
        RECT 54.290 102.870 54.610 103.130 ;
        RECT 61.650 103.070 61.970 103.130 ;
        RECT 63.505 103.070 63.795 103.115 ;
        RECT 61.650 102.930 63.795 103.070 ;
        RECT 61.650 102.870 61.970 102.930 ;
        RECT 63.505 102.885 63.795 102.930 ;
        RECT 81.890 103.070 82.210 103.130 ;
        RECT 94.860 103.070 95.000 103.565 ;
        RECT 109.030 103.550 109.395 103.770 ;
        RECT 109.105 103.455 109.395 103.550 ;
        RECT 105.805 103.410 106.455 103.455 ;
        RECT 109.105 103.410 109.695 103.455 ;
        RECT 105.805 103.270 109.695 103.410 ;
        RECT 105.805 103.225 106.455 103.270 ;
        RECT 109.405 103.225 109.695 103.270 ;
        RECT 110.410 103.410 110.730 103.470 ;
        RECT 113.125 103.455 113.415 103.770 ;
        RECT 114.205 103.750 114.495 103.795 ;
        RECT 117.785 103.750 118.075 103.795 ;
        RECT 119.620 103.750 119.910 103.795 ;
        RECT 114.205 103.610 119.910 103.750 ;
        RECT 114.205 103.565 114.495 103.610 ;
        RECT 117.785 103.565 118.075 103.610 ;
        RECT 119.620 103.565 119.910 103.610 ;
        RECT 112.825 103.410 113.415 103.455 ;
        RECT 116.065 103.410 116.715 103.455 ;
        RECT 110.410 103.270 116.715 103.410 ;
        RECT 110.410 103.210 110.730 103.270 ;
        RECT 112.825 103.225 113.115 103.270 ;
        RECT 116.065 103.225 116.715 103.270 ;
        RECT 81.890 102.930 95.000 103.070 ;
        RECT 81.890 102.870 82.210 102.930 ;
        RECT 110.870 102.870 111.190 103.130 ;
        RECT 125.130 102.870 125.450 103.130 ;
        RECT 38.650 101.850 38.970 102.110 ;
        RECT 39.110 102.050 39.430 102.110 ;
        RECT 39.585 102.050 39.875 102.095 ;
        RECT 39.110 101.910 39.875 102.050 ;
        RECT 39.110 101.850 39.430 101.910 ;
        RECT 39.585 101.865 39.875 101.910 ;
        RECT 36.825 101.710 37.115 101.755 ;
        RECT 40.950 101.710 41.270 101.770 ;
        RECT 36.825 101.570 41.270 101.710 ;
        RECT 36.825 101.525 37.115 101.570 ;
        RECT 40.950 101.510 41.270 101.570 ;
        RECT 49.705 101.710 49.995 101.755 ;
        RECT 54.290 101.710 54.610 101.770 ;
        RECT 49.705 101.570 54.610 101.710 ;
        RECT 49.705 101.525 49.995 101.570 ;
        RECT 54.290 101.510 54.610 101.570 ;
        RECT 61.650 101.510 61.970 101.770 ;
        RECT 63.505 101.710 63.795 101.755 ;
        RECT 63.950 101.710 64.270 101.770 ;
        RECT 63.505 101.570 64.270 101.710 ;
        RECT 63.505 101.525 63.795 101.570 ;
        RECT 63.950 101.510 64.270 101.570 ;
        RECT 76.385 101.710 76.675 101.755 ;
        RECT 77.750 101.710 78.070 101.770 ;
        RECT 76.385 101.570 78.070 101.710 ;
        RECT 76.385 101.525 76.675 101.570 ;
        RECT 77.750 101.510 78.070 101.570 ;
        RECT 89.265 101.710 89.555 101.755 ;
        RECT 90.170 101.710 90.490 101.770 ;
        RECT 89.265 101.570 90.490 101.710 ;
        RECT 89.265 101.525 89.555 101.570 ;
        RECT 90.170 101.510 90.490 101.570 ;
        RECT 110.870 101.510 111.190 101.770 ;
        RECT 115.010 101.510 115.330 101.770 ;
        RECT 39.125 101.370 39.415 101.415 ;
        RECT 39.570 101.370 39.890 101.430 ;
        RECT 39.125 101.230 39.890 101.370 ;
        RECT 39.125 101.185 39.415 101.230 ;
        RECT 39.570 101.170 39.890 101.230 ;
        RECT 40.505 101.370 40.795 101.415 ;
        RECT 42.330 101.370 42.650 101.430 ;
        RECT 40.505 101.230 42.650 101.370 ;
        RECT 40.505 101.185 40.795 101.230 ;
        RECT 42.330 101.170 42.650 101.230 ;
        RECT 75.450 101.370 75.770 101.430 ;
        RECT 125.130 101.370 125.450 101.430 ;
        RECT 75.450 101.230 125.450 101.370 ;
        RECT 75.450 101.170 75.770 101.230 ;
        RECT 125.130 101.170 125.450 101.230 ;
        RECT 30.385 100.690 30.675 100.735 ;
        RECT 44.170 100.690 44.490 100.750 ;
        RECT 30.385 100.550 44.490 100.690 ;
        RECT 30.385 100.505 30.675 100.550 ;
        RECT 44.170 100.490 44.490 100.550 ;
        RECT 43.265 100.350 43.555 100.395 ;
        RECT 54.750 100.350 55.070 100.410 ;
        RECT 43.265 100.210 55.070 100.350 ;
        RECT 43.265 100.165 43.555 100.210 ;
        RECT 54.750 100.150 55.070 100.210 ;
        RECT 55.225 100.350 55.515 100.395 ;
        RECT 60.730 100.350 61.050 100.410 ;
        RECT 55.225 100.210 61.050 100.350 ;
        RECT 55.225 100.165 55.515 100.210 ;
        RECT 60.730 100.150 61.050 100.210 ;
        RECT 68.090 100.350 68.410 100.410 ;
        RECT 69.945 100.350 70.235 100.395 ;
        RECT 68.090 100.210 70.235 100.350 ;
        RECT 68.090 100.150 68.410 100.210 ;
        RECT 69.945 100.165 70.235 100.210 ;
        RECT 80.050 100.350 80.370 100.410 ;
        RECT 82.825 100.350 83.115 100.395 ;
        RECT 80.050 100.210 83.115 100.350 ;
        RECT 80.050 100.150 80.370 100.210 ;
        RECT 82.825 100.165 83.115 100.210 ;
        RECT 93.850 100.350 94.170 100.410 ;
        RECT 95.705 100.350 95.995 100.395 ;
        RECT 93.850 100.210 95.995 100.350 ;
        RECT 93.850 100.150 94.170 100.210 ;
        RECT 95.705 100.165 95.995 100.210 ;
        RECT 103.970 100.350 104.290 100.410 ;
        RECT 104.445 100.350 104.735 100.395 ;
        RECT 103.970 100.210 104.735 100.350 ;
        RECT 103.970 100.150 104.290 100.210 ;
        RECT 104.445 100.165 104.735 100.210 ;
        RECT 115.930 100.350 116.250 100.410 ;
        RECT 121.465 100.350 121.755 100.395 ;
        RECT 115.930 100.210 121.755 100.350 ;
        RECT 115.930 100.150 116.250 100.210 ;
        RECT 121.465 100.165 121.755 100.210 ;
        RECT 21.115 74.380 23.065 74.390 ;
        RECT 19.415 73.240 23.065 74.380 ;
        RECT 19.415 73.230 21.125 73.240 ;
        RECT 28.135 73.230 30.305 74.410 ;
        RECT 32.315 74.390 34.265 74.400 ;
        RECT 30.615 73.250 34.265 74.390 ;
        RECT 30.615 73.240 32.325 73.250 ;
        RECT 39.425 73.200 41.595 74.380 ;
        RECT 43.535 74.360 45.485 74.370 ;
        RECT 41.835 73.220 45.485 74.360 ;
        RECT 54.785 74.340 56.735 74.350 ;
        RECT 41.835 73.210 43.545 73.220 ;
        RECT 50.005 73.140 52.175 74.320 ;
        RECT 53.085 73.200 56.735 74.340 ;
        RECT 53.085 73.190 54.795 73.200 ;
        RECT 61.425 73.170 63.595 74.350 ;
        RECT 66.005 74.330 67.955 74.340 ;
        RECT 64.305 73.190 67.955 74.330 ;
        RECT 64.305 73.180 66.015 73.190 ;
        RECT 72.535 73.180 74.705 74.360 ;
        RECT 77.245 74.320 79.195 74.330 ;
        RECT 75.545 73.180 79.195 74.320 ;
        RECT 75.545 73.170 77.255 73.180 ;
        RECT 83.805 73.170 85.975 74.350 ;
        RECT 88.495 74.330 90.445 74.340 ;
        RECT 86.795 73.190 90.445 74.330 ;
        RECT 99.775 74.320 101.725 74.330 ;
        RECT 86.795 73.180 88.505 73.190 ;
        RECT 94.995 73.110 97.165 74.290 ;
        RECT 98.075 73.180 101.725 74.320 ;
        RECT 98.075 73.170 99.785 73.180 ;
        RECT 106.405 73.160 108.575 74.340 ;
        RECT 111.045 74.320 112.995 74.330 ;
        RECT 109.345 73.180 112.995 74.320 ;
        RECT 109.345 73.170 111.055 73.180 ;
        RECT 117.605 73.160 119.775 74.340 ;
        RECT 122.295 74.320 124.245 74.330 ;
        RECT 120.595 73.180 124.245 74.320 ;
        RECT 129.455 73.240 131.625 74.420 ;
        RECT 120.595 73.170 122.305 73.180 ;
        RECT 26.495 65.190 26.725 65.320 ;
        RECT 26.435 55.240 26.805 65.190 ;
        RECT 27.635 65.150 27.865 65.320 ;
        RECT 27.565 55.200 27.935 65.150 ;
        RECT 28.925 65.140 29.155 65.320 ;
        RECT 37.695 65.200 37.925 65.330 ;
        RECT 28.835 55.250 29.255 65.140 ;
        RECT 37.635 55.250 38.005 65.200 ;
        RECT 38.835 65.160 39.065 65.330 ;
        RECT 38.765 55.210 39.135 65.160 ;
        RECT 40.125 65.150 40.355 65.330 ;
        RECT 48.915 65.170 49.145 65.300 ;
        RECT 40.035 55.260 40.455 65.150 ;
        RECT 48.855 55.220 49.225 65.170 ;
        RECT 50.055 65.130 50.285 65.300 ;
        RECT 49.985 55.180 50.355 65.130 ;
        RECT 51.345 65.120 51.575 65.300 ;
        RECT 60.165 65.150 60.395 65.280 ;
        RECT 51.255 55.230 51.675 65.120 ;
        RECT 60.105 55.200 60.475 65.150 ;
        RECT 61.305 65.110 61.535 65.280 ;
        RECT 61.235 55.160 61.605 65.110 ;
        RECT 62.595 65.100 62.825 65.280 ;
        RECT 71.385 65.140 71.615 65.270 ;
        RECT 62.505 55.210 62.925 65.100 ;
        RECT 71.325 55.190 71.695 65.140 ;
        RECT 72.525 65.100 72.755 65.270 ;
        RECT 72.455 55.150 72.825 65.100 ;
        RECT 73.815 65.090 74.045 65.270 ;
        RECT 82.625 65.130 82.855 65.260 ;
        RECT 73.725 55.200 74.145 65.090 ;
        RECT 82.565 55.180 82.935 65.130 ;
        RECT 83.765 65.090 83.995 65.260 ;
        RECT 83.695 55.140 84.065 65.090 ;
        RECT 85.055 65.080 85.285 65.260 ;
        RECT 93.875 65.140 94.105 65.270 ;
        RECT 84.965 55.190 85.385 65.080 ;
        RECT 93.815 55.190 94.185 65.140 ;
        RECT 95.015 65.100 95.245 65.270 ;
        RECT 94.945 55.150 95.315 65.100 ;
        RECT 96.305 65.090 96.535 65.270 ;
        RECT 105.155 65.130 105.385 65.260 ;
        RECT 96.215 55.200 96.635 65.090 ;
        RECT 105.095 55.180 105.465 65.130 ;
        RECT 106.295 65.090 106.525 65.260 ;
        RECT 106.225 55.140 106.595 65.090 ;
        RECT 107.585 65.080 107.815 65.260 ;
        RECT 116.425 65.130 116.655 65.260 ;
        RECT 107.495 55.190 107.915 65.080 ;
        RECT 116.365 55.180 116.735 65.130 ;
        RECT 117.565 65.090 117.795 65.260 ;
        RECT 117.495 55.140 117.865 65.090 ;
        RECT 118.855 65.080 119.085 65.260 ;
        RECT 127.675 65.130 127.905 65.260 ;
        RECT 118.765 55.190 119.185 65.080 ;
        RECT 127.615 55.180 127.985 65.130 ;
        RECT 128.815 65.090 129.045 65.260 ;
        RECT 128.745 55.140 129.115 65.090 ;
        RECT 130.105 65.080 130.335 65.260 ;
        RECT 130.015 55.190 130.435 65.080 ;
        RECT 21.655 52.320 22.115 52.550 ;
        RECT 25.625 52.280 26.255 52.560 ;
        RECT 25.735 52.240 26.195 52.280 ;
        RECT 27.665 52.240 28.125 52.470 ;
        RECT 32.855 52.330 33.315 52.560 ;
        RECT 36.825 52.290 37.455 52.570 ;
        RECT 36.935 52.250 37.395 52.290 ;
        RECT 38.865 52.250 39.325 52.480 ;
        RECT 44.075 52.300 44.535 52.530 ;
        RECT 48.045 52.260 48.675 52.540 ;
        RECT 48.155 52.220 48.615 52.260 ;
        RECT 50.085 52.220 50.545 52.450 ;
        RECT 55.325 52.280 55.785 52.510 ;
        RECT 59.295 52.240 59.925 52.520 ;
        RECT 59.405 52.200 59.865 52.240 ;
        RECT 61.335 52.200 61.795 52.430 ;
        RECT 66.545 52.270 67.005 52.500 ;
        RECT 70.515 52.230 71.145 52.510 ;
        RECT 70.625 52.190 71.085 52.230 ;
        RECT 72.555 52.190 73.015 52.420 ;
        RECT 77.785 52.260 78.245 52.490 ;
        RECT 81.755 52.220 82.385 52.500 ;
        RECT 81.865 52.180 82.325 52.220 ;
        RECT 83.795 52.180 84.255 52.410 ;
        RECT 89.035 52.270 89.495 52.500 ;
        RECT 93.005 52.230 93.635 52.510 ;
        RECT 93.115 52.190 93.575 52.230 ;
        RECT 95.045 52.190 95.505 52.420 ;
        RECT 100.315 52.260 100.775 52.490 ;
        RECT 104.285 52.220 104.915 52.500 ;
        RECT 104.395 52.180 104.855 52.220 ;
        RECT 106.325 52.180 106.785 52.410 ;
        RECT 111.585 52.260 112.045 52.490 ;
        RECT 115.555 52.220 116.185 52.500 ;
        RECT 115.665 52.180 116.125 52.220 ;
        RECT 117.595 52.180 118.055 52.410 ;
        RECT 122.835 52.260 123.295 52.490 ;
        RECT 126.805 52.220 127.435 52.500 ;
        RECT 126.915 52.180 127.375 52.220 ;
        RECT 128.845 52.180 129.305 52.410 ;
        RECT 22.165 51.890 22.395 52.115 ;
        RECT 26.245 51.970 26.475 52.035 ;
        RECT 27.385 51.970 27.615 52.035 ;
        RECT 22.155 50.210 22.525 51.890 ;
        RECT 22.165 50.115 22.395 50.210 ;
        RECT 21.525 49.670 22.245 49.930 ;
        RECT 21.385 47.490 22.105 47.750 ;
        RECT 22.015 47.190 22.245 47.340 ;
        RECT 22.005 46.450 22.375 47.190 ;
        RECT 26.185 46.970 26.585 51.970 ;
        RECT 27.265 46.970 27.665 51.970 ;
        RECT 33.365 51.900 33.595 52.125 ;
        RECT 37.445 51.980 37.675 52.045 ;
        RECT 38.585 51.980 38.815 52.045 ;
        RECT 33.355 50.220 33.725 51.900 ;
        RECT 33.365 50.125 33.595 50.220 ;
        RECT 32.725 49.680 33.445 49.940 ;
        RECT 32.585 47.500 33.305 47.760 ;
        RECT 33.215 47.200 33.445 47.350 ;
        RECT 25.735 46.600 26.195 46.830 ;
        RECT 27.665 46.710 28.125 46.830 ;
        RECT 27.515 46.600 28.125 46.710 ;
        RECT 22.015 46.340 22.245 46.450 ;
        RECT 27.515 46.430 28.095 46.600 ;
        RECT 33.205 46.460 33.575 47.200 ;
        RECT 37.385 46.980 37.785 51.980 ;
        RECT 38.465 46.980 38.865 51.980 ;
        RECT 44.585 51.870 44.815 52.095 ;
        RECT 48.665 51.950 48.895 52.015 ;
        RECT 49.805 51.950 50.035 52.015 ;
        RECT 44.575 50.190 44.945 51.870 ;
        RECT 44.585 50.095 44.815 50.190 ;
        RECT 43.945 49.650 44.665 49.910 ;
        RECT 43.805 47.470 44.525 47.730 ;
        RECT 44.435 47.170 44.665 47.320 ;
        RECT 36.935 46.610 37.395 46.840 ;
        RECT 38.865 46.720 39.325 46.840 ;
        RECT 38.715 46.610 39.325 46.720 ;
        RECT 33.215 46.350 33.445 46.460 ;
        RECT 38.715 46.440 39.295 46.610 ;
        RECT 44.425 46.430 44.795 47.170 ;
        RECT 48.605 46.950 49.005 51.950 ;
        RECT 49.685 46.950 50.085 51.950 ;
        RECT 55.835 51.850 56.065 52.075 ;
        RECT 59.915 51.930 60.145 51.995 ;
        RECT 61.055 51.930 61.285 51.995 ;
        RECT 55.825 50.170 56.195 51.850 ;
        RECT 55.835 50.075 56.065 50.170 ;
        RECT 55.195 49.630 55.915 49.890 ;
        RECT 55.055 47.450 55.775 47.710 ;
        RECT 55.685 47.150 55.915 47.300 ;
        RECT 48.155 46.580 48.615 46.810 ;
        RECT 50.085 46.690 50.545 46.810 ;
        RECT 49.935 46.580 50.545 46.690 ;
        RECT 44.435 46.320 44.665 46.430 ;
        RECT 49.935 46.410 50.515 46.580 ;
        RECT 55.675 46.410 56.045 47.150 ;
        RECT 59.855 46.930 60.255 51.930 ;
        RECT 60.935 46.930 61.335 51.930 ;
        RECT 67.055 51.840 67.285 52.065 ;
        RECT 71.135 51.920 71.365 51.985 ;
        RECT 72.275 51.920 72.505 51.985 ;
        RECT 67.045 50.160 67.415 51.840 ;
        RECT 67.055 50.065 67.285 50.160 ;
        RECT 66.415 49.620 67.135 49.880 ;
        RECT 66.275 47.440 66.995 47.700 ;
        RECT 66.905 47.140 67.135 47.290 ;
        RECT 59.405 46.560 59.865 46.790 ;
        RECT 61.335 46.670 61.795 46.790 ;
        RECT 61.185 46.560 61.795 46.670 ;
        RECT 55.685 46.300 55.915 46.410 ;
        RECT 61.185 46.390 61.765 46.560 ;
        RECT 66.895 46.400 67.265 47.140 ;
        RECT 71.075 46.920 71.475 51.920 ;
        RECT 72.155 46.920 72.555 51.920 ;
        RECT 78.295 51.830 78.525 52.055 ;
        RECT 82.375 51.910 82.605 51.975 ;
        RECT 83.515 51.910 83.745 51.975 ;
        RECT 78.285 50.150 78.655 51.830 ;
        RECT 78.295 50.055 78.525 50.150 ;
        RECT 77.655 49.610 78.375 49.870 ;
        RECT 77.515 47.430 78.235 47.690 ;
        RECT 78.145 47.130 78.375 47.280 ;
        RECT 70.625 46.550 71.085 46.780 ;
        RECT 72.555 46.660 73.015 46.780 ;
        RECT 72.405 46.550 73.015 46.660 ;
        RECT 66.905 46.290 67.135 46.400 ;
        RECT 72.405 46.380 72.985 46.550 ;
        RECT 78.135 46.390 78.505 47.130 ;
        RECT 82.315 46.910 82.715 51.910 ;
        RECT 83.395 46.910 83.795 51.910 ;
        RECT 89.545 51.840 89.775 52.065 ;
        RECT 93.625 51.920 93.855 51.985 ;
        RECT 94.765 51.920 94.995 51.985 ;
        RECT 89.535 50.160 89.905 51.840 ;
        RECT 89.545 50.065 89.775 50.160 ;
        RECT 88.905 49.620 89.625 49.880 ;
        RECT 88.765 47.440 89.485 47.700 ;
        RECT 89.395 47.140 89.625 47.290 ;
        RECT 81.865 46.540 82.325 46.770 ;
        RECT 83.795 46.650 84.255 46.770 ;
        RECT 83.645 46.540 84.255 46.650 ;
        RECT 78.145 46.280 78.375 46.390 ;
        RECT 83.645 46.370 84.225 46.540 ;
        RECT 89.385 46.400 89.755 47.140 ;
        RECT 93.565 46.920 93.965 51.920 ;
        RECT 94.645 46.920 95.045 51.920 ;
        RECT 100.825 51.830 101.055 52.055 ;
        RECT 104.905 51.910 105.135 51.975 ;
        RECT 106.045 51.910 106.275 51.975 ;
        RECT 100.815 50.150 101.185 51.830 ;
        RECT 100.825 50.055 101.055 50.150 ;
        RECT 100.185 49.610 100.905 49.870 ;
        RECT 100.045 47.430 100.765 47.690 ;
        RECT 100.675 47.130 100.905 47.280 ;
        RECT 93.115 46.550 93.575 46.780 ;
        RECT 95.045 46.660 95.505 46.780 ;
        RECT 94.895 46.550 95.505 46.660 ;
        RECT 89.395 46.290 89.625 46.400 ;
        RECT 94.895 46.380 95.475 46.550 ;
        RECT 100.665 46.390 101.035 47.130 ;
        RECT 104.845 46.910 105.245 51.910 ;
        RECT 105.925 46.910 106.325 51.910 ;
        RECT 112.095 51.830 112.325 52.055 ;
        RECT 116.175 51.910 116.405 51.975 ;
        RECT 117.315 51.910 117.545 51.975 ;
        RECT 112.085 50.150 112.455 51.830 ;
        RECT 112.095 50.055 112.325 50.150 ;
        RECT 111.455 49.610 112.175 49.870 ;
        RECT 111.315 47.430 112.035 47.690 ;
        RECT 111.945 47.130 112.175 47.280 ;
        RECT 104.395 46.540 104.855 46.770 ;
        RECT 106.325 46.650 106.785 46.770 ;
        RECT 106.175 46.540 106.785 46.650 ;
        RECT 100.675 46.280 100.905 46.390 ;
        RECT 106.175 46.370 106.755 46.540 ;
        RECT 111.935 46.390 112.305 47.130 ;
        RECT 116.115 46.910 116.515 51.910 ;
        RECT 117.195 46.910 117.595 51.910 ;
        RECT 123.345 51.830 123.575 52.055 ;
        RECT 127.425 51.910 127.655 51.975 ;
        RECT 128.565 51.910 128.795 51.975 ;
        RECT 123.335 50.150 123.705 51.830 ;
        RECT 123.345 50.055 123.575 50.150 ;
        RECT 122.705 49.610 123.425 49.870 ;
        RECT 122.565 47.430 123.285 47.690 ;
        RECT 123.195 47.130 123.425 47.280 ;
        RECT 115.665 46.540 116.125 46.770 ;
        RECT 117.595 46.650 118.055 46.770 ;
        RECT 117.445 46.540 118.055 46.650 ;
        RECT 111.945 46.280 112.175 46.390 ;
        RECT 117.445 46.370 118.025 46.540 ;
        RECT 123.185 46.390 123.555 47.130 ;
        RECT 127.365 46.910 127.765 51.910 ;
        RECT 128.445 46.910 128.845 51.910 ;
        RECT 126.915 46.540 127.375 46.770 ;
        RECT 128.845 46.650 129.305 46.770 ;
        RECT 128.695 46.540 129.305 46.650 ;
        RECT 123.195 46.280 123.425 46.390 ;
        RECT 128.695 46.370 129.275 46.540 ;
        RECT 21.505 45.950 21.965 46.180 ;
        RECT 32.705 45.960 33.165 46.190 ;
        RECT 43.925 45.930 44.385 46.160 ;
        RECT 55.175 45.910 55.635 46.140 ;
        RECT 66.395 45.900 66.855 46.130 ;
        RECT 77.635 45.890 78.095 46.120 ;
        RECT 88.885 45.900 89.345 46.130 ;
        RECT 100.165 45.890 100.625 46.120 ;
        RECT 111.435 45.890 111.895 46.120 ;
        RECT 122.685 45.890 123.145 46.120 ;
        RECT 26.775 39.230 27.235 39.460 ;
        RECT 38.055 39.230 38.515 39.460 ;
        RECT 49.345 39.210 49.805 39.440 ;
        RECT 60.565 39.210 61.025 39.440 ;
        RECT 71.765 39.210 72.225 39.440 ;
        RECT 83.055 39.200 83.515 39.430 ;
        RECT 94.295 39.220 94.755 39.450 ;
        RECT 105.505 39.240 105.965 39.470 ;
        RECT 116.705 39.280 117.165 39.510 ;
        RECT 127.915 39.300 128.375 39.530 ;
        RECT 20.645 38.810 21.225 38.980 ;
        RECT 26.495 38.960 26.725 39.070 ;
        RECT 20.615 38.700 21.225 38.810 ;
        RECT 20.615 38.580 21.075 38.700 ;
        RECT 22.545 38.580 23.005 38.810 ;
        RECT 21.075 33.440 21.475 38.440 ;
        RECT 22.155 33.440 22.555 38.440 ;
        RECT 26.365 38.220 26.735 38.960 ;
        RECT 31.925 38.810 32.505 38.980 ;
        RECT 37.775 38.960 38.005 39.070 ;
        RECT 31.895 38.700 32.505 38.810 ;
        RECT 31.895 38.580 32.355 38.700 ;
        RECT 33.825 38.580 34.285 38.810 ;
        RECT 26.495 38.070 26.725 38.220 ;
        RECT 26.635 37.660 27.355 37.920 ;
        RECT 26.495 35.480 27.215 35.740 ;
        RECT 26.345 35.200 26.575 35.295 ;
        RECT 26.215 33.520 26.585 35.200 ;
        RECT 21.125 33.375 21.355 33.440 ;
        RECT 22.265 33.375 22.495 33.440 ;
        RECT 26.345 33.295 26.575 33.520 ;
        RECT 32.355 33.440 32.755 38.440 ;
        RECT 33.435 33.440 33.835 38.440 ;
        RECT 37.645 38.220 38.015 38.960 ;
        RECT 43.215 38.790 43.795 38.960 ;
        RECT 49.065 38.940 49.295 39.050 ;
        RECT 43.185 38.680 43.795 38.790 ;
        RECT 43.185 38.560 43.645 38.680 ;
        RECT 45.115 38.560 45.575 38.790 ;
        RECT 37.775 38.070 38.005 38.220 ;
        RECT 37.915 37.660 38.635 37.920 ;
        RECT 37.775 35.480 38.495 35.740 ;
        RECT 37.625 35.200 37.855 35.295 ;
        RECT 37.495 33.520 37.865 35.200 ;
        RECT 32.405 33.375 32.635 33.440 ;
        RECT 33.545 33.375 33.775 33.440 ;
        RECT 37.625 33.295 37.855 33.520 ;
        RECT 43.645 33.420 44.045 38.420 ;
        RECT 44.725 33.420 45.125 38.420 ;
        RECT 48.935 38.200 49.305 38.940 ;
        RECT 54.435 38.790 55.015 38.960 ;
        RECT 60.285 38.940 60.515 39.050 ;
        RECT 54.405 38.680 55.015 38.790 ;
        RECT 54.405 38.560 54.865 38.680 ;
        RECT 56.335 38.560 56.795 38.790 ;
        RECT 49.065 38.050 49.295 38.200 ;
        RECT 49.205 37.640 49.925 37.900 ;
        RECT 49.065 35.460 49.785 35.720 ;
        RECT 48.915 35.180 49.145 35.275 ;
        RECT 48.785 33.500 49.155 35.180 ;
        RECT 43.695 33.355 43.925 33.420 ;
        RECT 44.835 33.355 45.065 33.420 ;
        RECT 48.915 33.275 49.145 33.500 ;
        RECT 54.865 33.420 55.265 38.420 ;
        RECT 55.945 33.420 56.345 38.420 ;
        RECT 60.155 38.200 60.525 38.940 ;
        RECT 65.635 38.790 66.215 38.960 ;
        RECT 71.485 38.940 71.715 39.050 ;
        RECT 65.605 38.680 66.215 38.790 ;
        RECT 65.605 38.560 66.065 38.680 ;
        RECT 67.535 38.560 67.995 38.790 ;
        RECT 60.285 38.050 60.515 38.200 ;
        RECT 60.425 37.640 61.145 37.900 ;
        RECT 60.285 35.460 61.005 35.720 ;
        RECT 60.135 35.180 60.365 35.275 ;
        RECT 60.005 33.500 60.375 35.180 ;
        RECT 54.915 33.355 55.145 33.420 ;
        RECT 56.055 33.355 56.285 33.420 ;
        RECT 60.135 33.275 60.365 33.500 ;
        RECT 66.065 33.420 66.465 38.420 ;
        RECT 67.145 33.420 67.545 38.420 ;
        RECT 71.355 38.200 71.725 38.940 ;
        RECT 76.925 38.780 77.505 38.950 ;
        RECT 82.775 38.930 83.005 39.040 ;
        RECT 76.895 38.670 77.505 38.780 ;
        RECT 76.895 38.550 77.355 38.670 ;
        RECT 78.825 38.550 79.285 38.780 ;
        RECT 71.485 38.050 71.715 38.200 ;
        RECT 71.625 37.640 72.345 37.900 ;
        RECT 71.485 35.460 72.205 35.720 ;
        RECT 71.335 35.180 71.565 35.275 ;
        RECT 71.205 33.500 71.575 35.180 ;
        RECT 66.115 33.355 66.345 33.420 ;
        RECT 67.255 33.355 67.485 33.420 ;
        RECT 71.335 33.275 71.565 33.500 ;
        RECT 77.355 33.410 77.755 38.410 ;
        RECT 78.435 33.410 78.835 38.410 ;
        RECT 82.645 38.190 83.015 38.930 ;
        RECT 88.165 38.800 88.745 38.970 ;
        RECT 94.015 38.950 94.245 39.060 ;
        RECT 88.135 38.690 88.745 38.800 ;
        RECT 88.135 38.570 88.595 38.690 ;
        RECT 90.065 38.570 90.525 38.800 ;
        RECT 82.775 38.040 83.005 38.190 ;
        RECT 82.915 37.630 83.635 37.890 ;
        RECT 82.775 35.450 83.495 35.710 ;
        RECT 82.625 35.170 82.855 35.265 ;
        RECT 82.495 33.490 82.865 35.170 ;
        RECT 77.405 33.345 77.635 33.410 ;
        RECT 78.545 33.345 78.775 33.410 ;
        RECT 82.625 33.265 82.855 33.490 ;
        RECT 88.595 33.430 88.995 38.430 ;
        RECT 89.675 33.430 90.075 38.430 ;
        RECT 93.885 38.210 94.255 38.950 ;
        RECT 99.375 38.820 99.955 38.990 ;
        RECT 105.225 38.970 105.455 39.080 ;
        RECT 99.345 38.710 99.955 38.820 ;
        RECT 99.345 38.590 99.805 38.710 ;
        RECT 101.275 38.590 101.735 38.820 ;
        RECT 94.015 38.060 94.245 38.210 ;
        RECT 94.155 37.650 94.875 37.910 ;
        RECT 94.015 35.470 94.735 35.730 ;
        RECT 93.865 35.190 94.095 35.285 ;
        RECT 93.735 33.510 94.105 35.190 ;
        RECT 88.645 33.365 88.875 33.430 ;
        RECT 89.785 33.365 90.015 33.430 ;
        RECT 93.865 33.285 94.095 33.510 ;
        RECT 99.805 33.450 100.205 38.450 ;
        RECT 100.885 33.450 101.285 38.450 ;
        RECT 105.095 38.230 105.465 38.970 ;
        RECT 110.575 38.860 111.155 39.030 ;
        RECT 116.425 39.010 116.655 39.120 ;
        RECT 110.545 38.750 111.155 38.860 ;
        RECT 110.545 38.630 111.005 38.750 ;
        RECT 112.475 38.630 112.935 38.860 ;
        RECT 105.225 38.080 105.455 38.230 ;
        RECT 105.365 37.670 106.085 37.930 ;
        RECT 105.225 35.490 105.945 35.750 ;
        RECT 105.075 35.210 105.305 35.305 ;
        RECT 104.945 33.530 105.315 35.210 ;
        RECT 99.855 33.385 100.085 33.450 ;
        RECT 100.995 33.385 101.225 33.450 ;
        RECT 105.075 33.305 105.305 33.530 ;
        RECT 111.005 33.490 111.405 38.490 ;
        RECT 112.085 33.490 112.485 38.490 ;
        RECT 116.295 38.270 116.665 39.010 ;
        RECT 121.785 38.880 122.365 39.050 ;
        RECT 127.635 39.030 127.865 39.140 ;
        RECT 121.755 38.770 122.365 38.880 ;
        RECT 121.755 38.650 122.215 38.770 ;
        RECT 123.685 38.650 124.145 38.880 ;
        RECT 116.425 38.120 116.655 38.270 ;
        RECT 116.565 37.710 117.285 37.970 ;
        RECT 116.425 35.530 117.145 35.790 ;
        RECT 116.275 35.250 116.505 35.345 ;
        RECT 116.145 33.570 116.515 35.250 ;
        RECT 111.055 33.425 111.285 33.490 ;
        RECT 112.195 33.425 112.425 33.490 ;
        RECT 116.275 33.345 116.505 33.570 ;
        RECT 122.215 33.510 122.615 38.510 ;
        RECT 123.295 33.510 123.695 38.510 ;
        RECT 127.505 38.290 127.875 39.030 ;
        RECT 127.635 38.140 127.865 38.290 ;
        RECT 127.775 37.730 128.495 37.990 ;
        RECT 127.635 35.550 128.355 35.810 ;
        RECT 127.485 35.270 127.715 35.365 ;
        RECT 127.355 33.590 127.725 35.270 ;
        RECT 122.265 33.445 122.495 33.510 ;
        RECT 123.405 33.445 123.635 33.510 ;
        RECT 127.485 33.365 127.715 33.590 ;
        RECT 20.615 32.940 21.075 33.170 ;
        RECT 22.545 33.130 23.005 33.170 ;
        RECT 22.485 32.850 23.115 33.130 ;
        RECT 26.625 32.860 27.085 33.090 ;
        RECT 31.895 32.940 32.355 33.170 ;
        RECT 33.825 33.130 34.285 33.170 ;
        RECT 33.765 32.850 34.395 33.130 ;
        RECT 37.905 32.860 38.365 33.090 ;
        RECT 43.185 32.920 43.645 33.150 ;
        RECT 45.115 33.110 45.575 33.150 ;
        RECT 45.055 32.830 45.685 33.110 ;
        RECT 49.195 32.840 49.655 33.070 ;
        RECT 54.405 32.920 54.865 33.150 ;
        RECT 56.335 33.110 56.795 33.150 ;
        RECT 56.275 32.830 56.905 33.110 ;
        RECT 60.415 32.840 60.875 33.070 ;
        RECT 65.605 32.920 66.065 33.150 ;
        RECT 67.535 33.110 67.995 33.150 ;
        RECT 67.475 32.830 68.105 33.110 ;
        RECT 71.615 32.840 72.075 33.070 ;
        RECT 76.895 32.910 77.355 33.140 ;
        RECT 78.825 33.100 79.285 33.140 ;
        RECT 78.765 32.820 79.395 33.100 ;
        RECT 82.905 32.830 83.365 33.060 ;
        RECT 88.135 32.930 88.595 33.160 ;
        RECT 90.065 33.120 90.525 33.160 ;
        RECT 90.005 32.840 90.635 33.120 ;
        RECT 94.145 32.850 94.605 33.080 ;
        RECT 99.345 32.950 99.805 33.180 ;
        RECT 101.275 33.140 101.735 33.180 ;
        RECT 101.215 32.860 101.845 33.140 ;
        RECT 105.355 32.870 105.815 33.100 ;
        RECT 110.545 32.990 111.005 33.220 ;
        RECT 112.475 33.180 112.935 33.220 ;
        RECT 112.415 32.900 113.045 33.180 ;
        RECT 116.555 32.910 117.015 33.140 ;
        RECT 121.755 33.010 122.215 33.240 ;
        RECT 123.685 33.200 124.145 33.240 ;
        RECT 123.625 32.920 124.255 33.200 ;
        RECT 127.765 32.930 128.225 33.160 ;
        RECT 19.485 20.270 19.905 30.160 ;
        RECT 19.585 20.090 19.815 20.270 ;
        RECT 20.805 20.260 21.175 30.210 ;
        RECT 20.875 20.090 21.105 20.260 ;
        RECT 21.935 20.220 22.305 30.170 ;
        RECT 30.765 20.270 31.185 30.160 ;
        RECT 22.015 20.090 22.245 20.220 ;
        RECT 30.865 20.090 31.095 20.270 ;
        RECT 32.085 20.260 32.455 30.210 ;
        RECT 32.155 20.090 32.385 20.260 ;
        RECT 33.215 20.220 33.585 30.170 ;
        RECT 42.055 20.250 42.475 30.140 ;
        RECT 33.295 20.090 33.525 20.220 ;
        RECT 42.155 20.070 42.385 20.250 ;
        RECT 43.375 20.240 43.745 30.190 ;
        RECT 43.445 20.070 43.675 20.240 ;
        RECT 44.505 20.200 44.875 30.150 ;
        RECT 53.275 20.250 53.695 30.140 ;
        RECT 44.585 20.070 44.815 20.200 ;
        RECT 53.375 20.070 53.605 20.250 ;
        RECT 54.595 20.240 54.965 30.190 ;
        RECT 54.665 20.070 54.895 20.240 ;
        RECT 55.725 20.200 56.095 30.150 ;
        RECT 64.475 20.250 64.895 30.140 ;
        RECT 55.805 20.070 56.035 20.200 ;
        RECT 64.575 20.070 64.805 20.250 ;
        RECT 65.795 20.240 66.165 30.190 ;
        RECT 65.865 20.070 66.095 20.240 ;
        RECT 66.925 20.200 67.295 30.150 ;
        RECT 75.765 20.240 76.185 30.130 ;
        RECT 67.005 20.070 67.235 20.200 ;
        RECT 75.865 20.060 76.095 20.240 ;
        RECT 77.085 20.230 77.455 30.180 ;
        RECT 77.155 20.060 77.385 20.230 ;
        RECT 78.215 20.190 78.585 30.140 ;
        RECT 87.005 20.260 87.425 30.150 ;
        RECT 78.295 20.060 78.525 20.190 ;
        RECT 87.105 20.080 87.335 20.260 ;
        RECT 88.325 20.250 88.695 30.200 ;
        RECT 88.395 20.080 88.625 20.250 ;
        RECT 89.455 20.210 89.825 30.160 ;
        RECT 98.215 20.280 98.635 30.170 ;
        RECT 89.535 20.080 89.765 20.210 ;
        RECT 98.315 20.100 98.545 20.280 ;
        RECT 99.535 20.270 99.905 30.220 ;
        RECT 99.605 20.100 99.835 20.270 ;
        RECT 100.665 20.230 101.035 30.180 ;
        RECT 109.415 20.320 109.835 30.210 ;
        RECT 100.745 20.100 100.975 20.230 ;
        RECT 109.515 20.140 109.745 20.320 ;
        RECT 110.735 20.310 111.105 30.260 ;
        RECT 110.805 20.140 111.035 20.310 ;
        RECT 111.865 20.270 112.235 30.220 ;
        RECT 120.625 20.340 121.045 30.230 ;
        RECT 111.945 20.140 112.175 20.270 ;
        RECT 120.725 20.160 120.955 20.340 ;
        RECT 121.945 20.330 122.315 30.280 ;
        RECT 122.015 20.160 122.245 20.330 ;
        RECT 123.075 20.290 123.445 30.240 ;
        RECT 123.155 20.160 123.385 20.290 ;
        RECT 128.755 12.240 130.465 12.250 ;
        RECT 117.545 12.220 119.255 12.230 ;
        RECT 106.345 12.180 108.055 12.190 ;
        RECT 27.615 12.170 29.325 12.180 ;
        RECT 38.895 12.170 40.605 12.180 ;
        RECT 25.675 11.030 29.325 12.170 ;
        RECT 36.955 11.030 40.605 12.170 ;
        RECT 95.135 12.160 96.845 12.170 ;
        RECT 50.185 12.150 51.895 12.160 ;
        RECT 61.405 12.150 63.115 12.160 ;
        RECT 72.605 12.150 74.315 12.160 ;
        RECT 25.675 11.020 27.625 11.030 ;
        RECT 36.955 11.020 38.905 11.030 ;
        RECT 48.245 11.010 51.895 12.150 ;
        RECT 59.465 11.010 63.115 12.150 ;
        RECT 70.665 11.010 74.315 12.150 ;
        RECT 83.895 12.140 85.605 12.150 ;
        RECT 48.245 11.000 50.195 11.010 ;
        RECT 59.465 11.000 61.415 11.010 ;
        RECT 70.665 11.000 72.615 11.010 ;
        RECT 81.955 11.000 85.605 12.140 ;
        RECT 93.195 11.020 96.845 12.160 ;
        RECT 104.405 11.040 108.055 12.180 ;
        RECT 115.605 11.080 119.255 12.220 ;
        RECT 126.815 11.100 130.465 12.240 ;
        RECT 126.815 11.090 128.765 11.100 ;
        RECT 115.605 11.070 117.555 11.080 ;
        RECT 104.405 11.030 106.355 11.040 ;
        RECT 93.195 11.010 95.145 11.020 ;
        RECT 81.955 10.990 83.905 11.000 ;
      LAYER met2 ;
        RECT 81.000 207.220 81.260 207.540 ;
        RECT 71.340 206.880 71.600 207.200 ;
        RECT 75.480 206.880 75.740 207.200 ;
        RECT 71.400 205.500 71.540 206.880 ;
        RECT 75.020 206.200 75.280 206.520 ;
        RECT 75.080 205.500 75.220 206.200 ;
        RECT 71.340 205.180 71.600 205.500 ;
        RECT 75.020 205.180 75.280 205.500 ;
        RECT 65.360 203.480 65.620 203.800 ;
        RECT 69.040 203.480 69.300 203.800 ;
        RECT 61.680 201.780 61.940 202.100 ;
        RECT 60.300 201.440 60.560 201.760 ;
        RECT 55.240 196.000 55.500 196.320 ;
        RECT 52.020 195.320 52.280 195.640 ;
        RECT 52.080 194.280 52.220 195.320 ;
        RECT 52.020 193.960 52.280 194.280 ;
        RECT 37.760 193.280 38.020 193.600 ;
        RECT 45.120 193.280 45.380 193.600 ;
        RECT 37.820 188.500 37.960 193.280 ;
        RECT 45.180 191.900 45.320 193.280 ;
        RECT 50.640 192.600 50.900 192.920 ;
        RECT 52.940 192.600 53.200 192.920 ;
        RECT 45.120 191.580 45.380 191.900 ;
        RECT 42.820 190.900 43.080 191.220 ;
        RECT 47.880 190.900 48.140 191.220 ;
        RECT 38.220 190.220 38.480 190.540 ;
        RECT 34.540 188.180 34.800 188.500 ;
        RECT 35.920 188.180 36.180 188.500 ;
        RECT 37.760 188.180 38.020 188.500 ;
        RECT 30.400 187.840 30.660 188.160 ;
        RECT 25.800 185.120 26.060 185.440 ;
        RECT 25.860 179.320 26.000 185.120 ;
        RECT 30.460 185.100 30.600 187.840 ;
        RECT 34.600 185.440 34.740 188.180 ;
        RECT 35.980 186.120 36.120 188.180 ;
        RECT 35.920 185.800 36.180 186.120 ;
        RECT 35.460 185.460 35.720 185.780 ;
        RECT 34.540 185.120 34.800 185.440 ;
        RECT 27.180 184.780 27.440 185.100 ;
        RECT 30.400 184.780 30.660 185.100 ;
        RECT 27.240 183.740 27.380 184.780 ;
        RECT 31.320 184.440 31.580 184.760 ;
        RECT 27.180 183.420 27.440 183.740 ;
        RECT 26.260 179.340 26.520 179.660 ;
        RECT 27.640 179.340 27.900 179.660 ;
        RECT 25.800 179.000 26.060 179.320 ;
        RECT 26.320 178.300 26.460 179.340 ;
        RECT 27.700 178.300 27.840 179.340 ;
        RECT 26.260 177.980 26.520 178.300 ;
        RECT 27.640 177.980 27.900 178.300 ;
        RECT 26.260 177.300 26.520 177.620 ;
        RECT 28.100 177.300 28.360 177.620 ;
        RECT 29.940 177.300 30.200 177.620 ;
        RECT 26.320 174.560 26.460 177.300 ;
        RECT 27.640 176.280 27.900 176.600 ;
        RECT 27.700 174.560 27.840 176.280 ;
        RECT 28.160 175.240 28.300 177.300 ;
        RECT 30.000 175.580 30.140 177.300 ;
        RECT 29.940 175.260 30.200 175.580 ;
        RECT 28.100 174.920 28.360 175.240 ;
        RECT 26.260 174.240 26.520 174.560 ;
        RECT 27.640 174.240 27.900 174.560 ;
        RECT 31.380 173.880 31.520 184.440 ;
        RECT 34.080 183.080 34.340 183.400 ;
        RECT 34.140 174.900 34.280 183.080 ;
        RECT 34.540 182.740 34.800 183.060 ;
        RECT 34.600 180.340 34.740 182.740 ;
        RECT 35.520 182.720 35.660 185.460 ;
        RECT 36.380 184.440 36.640 184.760 ;
        RECT 35.460 182.400 35.720 182.720 ;
        RECT 34.540 180.020 34.800 180.340 ;
        RECT 34.080 174.580 34.340 174.900 ;
        RECT 31.320 173.560 31.580 173.880 ;
        RECT 31.380 169.120 31.520 173.560 ;
        RECT 34.600 172.180 34.740 180.020 ;
        RECT 35.000 176.960 35.260 177.280 ;
        RECT 35.060 174.560 35.200 176.960 ;
        RECT 35.520 176.600 35.660 182.400 ;
        RECT 36.440 182.380 36.580 184.440 ;
        RECT 36.380 182.060 36.640 182.380 ;
        RECT 36.440 180.000 36.580 182.060 ;
        RECT 36.380 179.680 36.640 180.000 ;
        RECT 35.460 176.280 35.720 176.600 ;
        RECT 35.520 175.240 35.660 176.280 ;
        RECT 35.460 174.920 35.720 175.240 ;
        RECT 35.000 174.240 35.260 174.560 ;
        RECT 35.920 174.240 36.180 174.560 ;
        RECT 35.980 172.520 36.120 174.240 ;
        RECT 35.920 172.200 36.180 172.520 ;
        RECT 34.540 171.860 34.800 172.180 ;
        RECT 35.460 171.180 35.720 171.500 ;
        RECT 22.580 168.800 22.840 169.120 ;
        RECT 31.320 168.800 31.580 169.120 ;
        RECT 34.080 168.800 34.340 169.120 ;
        RECT 22.640 167.080 22.780 168.800 ;
        RECT 27.640 168.120 27.900 168.440 ;
        RECT 22.580 166.760 22.840 167.080 ;
        RECT 25.800 166.080 26.060 166.400 ;
        RECT 27.180 166.080 27.440 166.400 ;
        RECT 25.860 164.700 26.000 166.080 ;
        RECT 25.800 164.380 26.060 164.700 ;
        RECT 26.720 163.360 26.980 163.680 ;
        RECT 26.260 162.680 26.520 163.000 ;
        RECT 18.900 161.320 19.160 161.640 ;
        RECT 18.960 159.260 19.100 161.320 ;
        RECT 25.800 160.640 26.060 160.960 ;
        RECT 21.660 159.960 21.920 160.280 ;
        RECT 18.900 158.940 19.160 159.260 ;
        RECT 21.720 158.580 21.860 159.960 ;
        RECT 25.860 159.260 26.000 160.640 ;
        RECT 26.320 160.140 26.460 162.680 ;
        RECT 26.780 161.980 26.920 163.360 ;
        RECT 26.720 161.660 26.980 161.980 ;
        RECT 27.240 161.300 27.380 166.080 ;
        RECT 27.700 163.340 27.840 168.120 ;
        RECT 31.380 167.420 31.520 168.800 ;
        RECT 31.320 167.100 31.580 167.420 ;
        RECT 34.140 165.720 34.280 168.800 ;
        RECT 35.000 168.120 35.260 168.440 ;
        RECT 35.060 166.400 35.200 168.120 ;
        RECT 35.000 166.080 35.260 166.400 ;
        RECT 34.080 165.400 34.340 165.720 ;
        RECT 27.640 163.020 27.900 163.340 ;
        RECT 27.180 160.980 27.440 161.300 ;
        RECT 26.320 160.000 26.920 160.140 ;
        RECT 25.800 158.940 26.060 159.260 ;
        RECT 21.200 158.260 21.460 158.580 ;
        RECT 21.660 158.260 21.920 158.580 ;
        RECT 18.900 157.920 19.160 158.240 ;
        RECT 18.960 144.980 19.100 157.920 ;
        RECT 19.360 157.240 19.620 157.560 ;
        RECT 19.420 156.200 19.560 157.240 ;
        RECT 19.360 155.880 19.620 156.200 ;
        RECT 21.260 153.140 21.400 158.260 ;
        RECT 21.660 157.240 21.920 157.560 ;
        RECT 21.720 156.540 21.860 157.240 ;
        RECT 26.780 156.540 26.920 160.000 ;
        RECT 21.660 156.220 21.920 156.540 ;
        RECT 26.720 156.220 26.980 156.540 ;
        RECT 21.720 153.140 21.860 156.220 ;
        RECT 27.240 155.940 27.380 160.980 ;
        RECT 31.320 160.300 31.580 160.620 ;
        RECT 30.400 159.960 30.660 160.280 ;
        RECT 25.860 155.800 27.380 155.940 ;
        RECT 25.860 155.520 26.000 155.800 ;
        RECT 25.800 155.200 26.060 155.520 ;
        RECT 26.720 155.200 26.980 155.520 ;
        RECT 21.200 152.820 21.460 153.140 ;
        RECT 21.660 152.820 21.920 153.140 ;
        RECT 20.740 150.440 21.000 150.760 ;
        RECT 20.800 145.660 20.940 150.440 ;
        RECT 21.260 147.700 21.400 152.820 ;
        RECT 25.340 152.480 25.600 152.800 ;
        RECT 22.580 151.800 22.840 152.120 ;
        RECT 22.640 149.400 22.780 151.800 ;
        RECT 23.500 149.760 23.760 150.080 ;
        RECT 22.580 149.080 22.840 149.400 ;
        RECT 22.120 147.720 22.380 148.040 ;
        RECT 21.200 147.380 21.460 147.700 ;
        RECT 22.180 146.680 22.320 147.720 ;
        RECT 22.640 147.360 22.780 149.080 ;
        RECT 23.560 148.380 23.700 149.760 ;
        RECT 23.500 148.060 23.760 148.380 ;
        RECT 23.960 147.380 24.220 147.700 ;
        RECT 22.580 147.040 22.840 147.360 ;
        RECT 24.020 146.680 24.160 147.380 ;
        RECT 25.400 147.360 25.540 152.480 ;
        RECT 25.860 150.080 26.000 155.200 ;
        RECT 26.780 153.820 26.920 155.200 ;
        RECT 26.720 153.500 26.980 153.820 ;
        RECT 30.460 153.140 30.600 159.960 ;
        RECT 31.380 158.920 31.520 160.300 ;
        RECT 31.320 158.600 31.580 158.920 ;
        RECT 31.380 153.480 31.520 158.600 ;
        RECT 34.140 155.520 34.280 165.400 ;
        RECT 35.060 161.980 35.200 166.080 ;
        RECT 35.000 161.660 35.260 161.980 ;
        RECT 35.000 160.980 35.260 161.300 ;
        RECT 34.540 160.640 34.800 160.960 ;
        RECT 34.600 156.540 34.740 160.640 ;
        RECT 35.060 159.260 35.200 160.980 ;
        RECT 35.000 158.940 35.260 159.260 ;
        RECT 34.540 156.220 34.800 156.540 ;
        RECT 34.080 155.200 34.340 155.520 ;
        RECT 31.320 153.160 31.580 153.480 ;
        RECT 30.400 152.820 30.660 153.140 ;
        RECT 31.380 152.540 31.520 153.160 ;
        RECT 34.600 152.800 34.740 156.220 ;
        RECT 30.920 152.400 31.520 152.540 ;
        RECT 34.540 152.480 34.800 152.800 ;
        RECT 25.800 149.760 26.060 150.080 ;
        RECT 30.920 147.360 31.060 152.400 ;
        RECT 31.320 151.800 31.580 152.120 ;
        RECT 33.160 151.800 33.420 152.120 ;
        RECT 35.000 151.800 35.260 152.120 ;
        RECT 31.380 150.760 31.520 151.800 ;
        RECT 33.220 151.180 33.360 151.800 ;
        RECT 33.220 151.040 34.740 151.180 ;
        RECT 31.320 150.440 31.580 150.760 ;
        RECT 34.600 150.420 34.740 151.040 ;
        RECT 34.540 150.100 34.800 150.420 ;
        RECT 25.340 147.040 25.600 147.360 ;
        RECT 29.480 147.040 29.740 147.360 ;
        RECT 30.860 147.040 31.120 147.360 ;
        RECT 22.120 146.360 22.380 146.680 ;
        RECT 23.960 146.360 24.220 146.680 ;
        RECT 22.180 145.660 22.320 146.360 ;
        RECT 25.400 145.660 25.540 147.040 ;
        RECT 29.540 146.680 29.680 147.040 ;
        RECT 25.800 146.360 26.060 146.680 ;
        RECT 27.180 146.360 27.440 146.680 ;
        RECT 29.480 146.360 29.740 146.680 ;
        RECT 20.740 145.340 21.000 145.660 ;
        RECT 22.120 145.340 22.380 145.660 ;
        RECT 25.340 145.340 25.600 145.660 ;
        RECT 25.400 144.980 25.540 145.340 ;
        RECT 25.860 145.320 26.000 146.360 ;
        RECT 25.800 145.000 26.060 145.320 ;
        RECT 18.900 144.660 19.160 144.980 ;
        RECT 25.340 144.660 25.600 144.980 ;
        RECT 27.240 144.640 27.380 146.360 ;
        RECT 27.180 144.320 27.440 144.640 ;
        RECT 35.060 141.920 35.200 151.800 ;
        RECT 35.520 142.600 35.660 171.180 ;
        RECT 35.920 170.840 36.180 171.160 ;
        RECT 35.980 166.140 36.120 170.840 ;
        RECT 36.440 169.460 36.580 179.680 ;
        RECT 37.300 179.340 37.560 179.660 ;
        RECT 37.360 174.560 37.500 179.340 ;
        RECT 37.820 179.320 37.960 188.180 ;
        RECT 38.280 186.460 38.420 190.220 ;
        RECT 40.060 189.880 40.320 190.200 ;
        RECT 38.220 186.140 38.480 186.460 ;
        RECT 39.600 184.780 39.860 185.100 ;
        RECT 39.660 182.040 39.800 184.780 ;
        RECT 40.120 182.720 40.260 189.880 ;
        RECT 41.440 187.160 41.700 187.480 ;
        RECT 41.500 184.760 41.640 187.160 ;
        RECT 40.980 184.440 41.240 184.760 ;
        RECT 41.440 184.440 41.700 184.760 ;
        RECT 41.900 184.440 42.160 184.760 ;
        RECT 40.060 182.400 40.320 182.720 ;
        RECT 39.600 181.720 39.860 182.040 ;
        RECT 39.140 179.680 39.400 180.000 ;
        RECT 37.760 179.000 38.020 179.320 ;
        RECT 38.680 179.000 38.940 179.320 ;
        RECT 37.820 177.620 37.960 179.000 ;
        RECT 38.740 177.960 38.880 179.000 ;
        RECT 39.200 178.300 39.340 179.680 ;
        RECT 39.660 178.300 39.800 181.720 ;
        RECT 39.140 177.980 39.400 178.300 ;
        RECT 39.600 177.980 39.860 178.300 ;
        RECT 40.120 177.960 40.260 182.400 ;
        RECT 41.040 181.020 41.180 184.440 ;
        RECT 40.980 180.700 41.240 181.020 ;
        RECT 38.680 177.640 38.940 177.960 ;
        RECT 40.060 177.640 40.320 177.960 ;
        RECT 37.760 177.300 38.020 177.620 ;
        RECT 37.300 174.240 37.560 174.560 ;
        RECT 37.360 172.180 37.500 174.240 ;
        RECT 37.300 171.860 37.560 172.180 ;
        RECT 36.380 169.140 36.640 169.460 ;
        RECT 37.820 169.120 37.960 177.300 ;
        RECT 40.060 176.280 40.320 176.600 ;
        RECT 40.120 174.900 40.260 176.280 ;
        RECT 40.520 174.920 40.780 175.240 ;
        RECT 40.060 174.580 40.320 174.900 ;
        RECT 38.220 173.900 38.480 174.220 ;
        RECT 37.760 168.800 38.020 169.120 ;
        RECT 36.370 166.565 36.650 166.935 ;
        RECT 37.300 166.760 37.560 167.080 ;
        RECT 36.380 166.420 36.640 166.565 ;
        RECT 35.980 166.000 36.580 166.140 ;
        RECT 35.920 162.680 36.180 163.000 ;
        RECT 35.980 158.580 36.120 162.680 ;
        RECT 35.920 158.260 36.180 158.580 ;
        RECT 35.920 148.060 36.180 148.380 ;
        RECT 35.980 147.360 36.120 148.060 ;
        RECT 35.920 147.040 36.180 147.360 ;
        RECT 35.920 142.620 36.180 142.940 ;
        RECT 35.460 142.280 35.720 142.600 ;
        RECT 35.000 141.600 35.260 141.920 ;
        RECT 24.880 140.920 25.140 141.240 ;
        RECT 18.440 139.560 18.700 139.880 ;
        RECT 17.060 135.820 17.320 136.140 ;
        RECT 17.120 134.100 17.260 135.820 ;
        RECT 18.500 134.780 18.640 139.560 ;
        RECT 23.500 138.880 23.760 139.200 ;
        RECT 19.360 138.200 19.620 138.520 ;
        RECT 19.420 134.780 19.560 138.200 ;
        RECT 23.560 137.500 23.700 138.880 ;
        RECT 23.500 137.180 23.760 137.500 ;
        RECT 21.200 136.160 21.460 136.480 ;
        RECT 23.500 136.160 23.760 136.480 ;
        RECT 21.260 134.780 21.400 136.160 ;
        RECT 18.440 134.460 18.700 134.780 ;
        RECT 19.360 134.460 19.620 134.780 ;
        RECT 21.200 134.460 21.460 134.780 ;
        RECT 17.060 133.780 17.320 134.100 ;
        RECT 19.420 131.040 19.560 134.460 ;
        RECT 20.740 133.440 21.000 133.760 ;
        RECT 20.800 131.380 20.940 133.440 ;
        RECT 20.740 131.060 21.000 131.380 ;
        RECT 19.360 130.720 19.620 131.040 ;
        RECT 20.800 129.420 20.940 131.060 ;
        RECT 23.040 130.040 23.300 130.360 ;
        RECT 20.800 129.280 21.400 129.420 ;
        RECT 20.740 128.680 21.000 129.000 ;
        RECT 20.800 125.600 20.940 128.680 ;
        RECT 21.260 126.280 21.400 129.280 ;
        RECT 21.200 125.960 21.460 126.280 ;
        RECT 20.740 125.280 21.000 125.600 ;
        RECT 18.900 122.900 19.160 123.220 ;
        RECT 14.300 114.740 14.560 115.060 ;
        RECT 14.360 91.170 14.500 114.740 ;
        RECT 17.980 108.280 18.240 108.600 ;
        RECT 18.040 107.580 18.180 108.280 ;
        RECT 18.960 107.580 19.100 122.900 ;
        RECT 21.260 120.500 21.400 125.960 ;
        RECT 23.100 125.600 23.240 130.040 ;
        RECT 21.660 125.280 21.920 125.600 ;
        RECT 23.040 125.280 23.300 125.600 ;
        RECT 21.720 120.840 21.860 125.280 ;
        RECT 23.560 120.840 23.700 136.160 ;
        RECT 23.960 135.480 24.220 135.800 ;
        RECT 24.020 134.440 24.160 135.480 ;
        RECT 23.960 134.120 24.220 134.440 ;
        RECT 24.420 130.380 24.680 130.700 ;
        RECT 24.480 129.340 24.620 130.380 ;
        RECT 24.420 129.020 24.680 129.340 ;
        RECT 24.420 128.000 24.680 128.320 ;
        RECT 24.480 126.620 24.620 128.000 ;
        RECT 24.420 126.300 24.680 126.620 ;
        RECT 24.940 126.020 25.080 140.920 ;
        RECT 35.980 140.220 36.120 142.620 ;
        RECT 35.920 139.900 36.180 140.220 ;
        RECT 25.800 139.560 26.060 139.880 ;
        RECT 24.480 125.880 25.080 126.020 ;
        RECT 23.960 121.880 24.220 122.200 ;
        RECT 21.660 120.520 21.920 120.840 ;
        RECT 22.580 120.520 22.840 120.840 ;
        RECT 23.500 120.520 23.760 120.840 ;
        RECT 21.200 120.180 21.460 120.500 ;
        RECT 21.200 119.160 21.460 119.480 ;
        RECT 22.120 119.160 22.380 119.480 ;
        RECT 21.260 118.460 21.400 119.160 ;
        RECT 21.200 118.140 21.460 118.460 ;
        RECT 21.660 117.800 21.920 118.120 ;
        RECT 21.720 115.740 21.860 117.800 ;
        RECT 21.660 115.420 21.920 115.740 ;
        RECT 20.740 113.720 21.000 114.040 ;
        RECT 20.800 112.680 20.940 113.720 ;
        RECT 22.180 113.020 22.320 119.160 ;
        RECT 22.640 114.720 22.780 120.520 ;
        RECT 23.040 119.160 23.300 119.480 ;
        RECT 23.100 114.720 23.240 119.160 ;
        RECT 24.020 117.860 24.160 121.880 ;
        RECT 24.480 121.260 24.620 125.880 ;
        RECT 25.860 122.620 26.000 139.560 ;
        RECT 26.260 138.880 26.520 139.200 ;
        RECT 26.320 133.760 26.460 138.880 ;
        RECT 30.860 138.540 31.120 138.860 ;
        RECT 30.920 135.800 31.060 138.540 ;
        RECT 36.440 136.820 36.580 166.000 ;
        RECT 37.360 164.360 37.500 166.760 ;
        RECT 37.820 166.060 37.960 168.800 ;
        RECT 37.760 165.740 38.020 166.060 ;
        RECT 37.820 164.700 37.960 165.740 ;
        RECT 37.760 164.380 38.020 164.700 ;
        RECT 37.300 164.040 37.560 164.360 ;
        RECT 37.820 164.020 37.960 164.380 ;
        RECT 37.760 163.700 38.020 164.020 ;
        RECT 37.300 152.480 37.560 152.800 ;
        RECT 37.360 150.760 37.500 152.480 ;
        RECT 37.300 150.440 37.560 150.760 ;
        RECT 37.360 146.680 37.500 150.440 ;
        RECT 37.300 146.360 37.560 146.680 ;
        RECT 36.840 144.320 37.100 144.640 ;
        RECT 34.080 136.500 34.340 136.820 ;
        RECT 36.380 136.500 36.640 136.820 ;
        RECT 30.400 135.480 30.660 135.800 ;
        RECT 30.860 135.480 31.120 135.800 ;
        RECT 32.700 135.480 32.960 135.800 ;
        RECT 30.460 134.180 30.600 135.480 ;
        RECT 30.920 134.780 31.060 135.480 ;
        RECT 30.860 134.460 31.120 134.780 ;
        RECT 31.780 134.180 32.040 134.440 ;
        RECT 30.460 134.120 32.040 134.180 ;
        RECT 30.460 134.040 31.980 134.120 ;
        RECT 32.760 134.100 32.900 135.480 ;
        RECT 26.260 133.440 26.520 133.760 ;
        RECT 26.320 128.660 26.460 133.440 ;
        RECT 30.460 132.060 30.600 134.040 ;
        RECT 32.700 133.780 32.960 134.100 ;
        RECT 34.140 133.760 34.280 136.500 ;
        RECT 35.460 135.480 35.720 135.800 ;
        RECT 34.080 133.670 34.340 133.760 ;
        RECT 34.080 133.530 34.740 133.670 ;
        RECT 34.080 133.440 34.340 133.530 ;
        RECT 30.860 132.760 31.120 133.080 ;
        RECT 30.400 131.740 30.660 132.060 ;
        RECT 27.640 130.040 27.900 130.360 ;
        RECT 26.260 128.340 26.520 128.660 ;
        RECT 26.320 123.560 26.460 128.340 ;
        RECT 27.180 125.280 27.440 125.600 ;
        RECT 26.720 124.600 26.980 124.920 ;
        RECT 26.260 123.240 26.520 123.560 ;
        RECT 25.860 122.480 26.460 122.620 ;
        RECT 24.480 121.120 26.000 121.260 ;
        RECT 25.340 119.160 25.600 119.480 ;
        RECT 24.020 117.720 25.080 117.860 ;
        RECT 25.400 117.780 25.540 119.160 ;
        RECT 22.580 114.400 22.840 114.720 ;
        RECT 23.040 114.400 23.300 114.720 ;
        RECT 23.960 113.720 24.220 114.040 ;
        RECT 22.120 112.700 22.380 113.020 ;
        RECT 20.740 112.360 21.000 112.680 ;
        RECT 24.020 112.340 24.160 113.720 ;
        RECT 23.960 112.020 24.220 112.340 ;
        RECT 20.280 111.000 20.540 111.320 ;
        RECT 17.980 107.260 18.240 107.580 ;
        RECT 18.900 107.260 19.160 107.580 ;
        RECT 20.340 91.170 20.480 111.000 ;
        RECT 23.040 108.960 23.300 109.280 ;
        RECT 22.580 106.920 22.840 107.240 ;
        RECT 22.640 104.860 22.780 106.920 ;
        RECT 23.100 106.560 23.240 108.960 ;
        RECT 23.040 106.240 23.300 106.560 ;
        RECT 22.580 104.540 22.840 104.860 ;
        RECT 23.100 103.840 23.240 106.240 ;
        RECT 23.040 103.520 23.300 103.840 ;
        RECT 24.940 101.540 25.080 117.720 ;
        RECT 25.340 117.460 25.600 117.780 ;
        RECT 25.340 114.060 25.600 114.380 ;
        RECT 25.400 107.580 25.540 114.060 ;
        RECT 25.860 109.280 26.000 121.120 ;
        RECT 26.320 111.840 26.460 122.480 ;
        RECT 26.780 120.160 26.920 124.600 ;
        RECT 27.240 120.500 27.380 125.280 ;
        RECT 27.700 125.260 27.840 130.040 ;
        RECT 28.100 127.660 28.360 127.980 ;
        RECT 28.160 125.600 28.300 127.660 ;
        RECT 28.100 125.280 28.360 125.600 ;
        RECT 27.640 124.940 27.900 125.260 ;
        RECT 27.180 120.180 27.440 120.500 ;
        RECT 26.720 119.840 26.980 120.160 ;
        RECT 30.400 119.160 30.660 119.480 ;
        RECT 30.460 118.120 30.600 119.160 ;
        RECT 30.400 117.800 30.660 118.120 ;
        RECT 26.720 117.460 26.980 117.780 ;
        RECT 26.780 112.420 26.920 117.460 ;
        RECT 26.780 112.340 27.840 112.420 ;
        RECT 28.100 112.360 28.360 112.680 ;
        RECT 26.720 112.280 27.840 112.340 ;
        RECT 26.720 112.020 26.980 112.280 ;
        RECT 26.320 111.700 26.920 111.840 ;
        RECT 26.780 109.280 26.920 111.700 ;
        RECT 25.800 108.960 26.060 109.280 ;
        RECT 26.720 108.960 26.980 109.280 ;
        RECT 27.180 108.620 27.440 108.940 ;
        RECT 25.340 107.260 25.600 107.580 ;
        RECT 27.240 104.520 27.380 108.620 ;
        RECT 27.700 106.560 27.840 112.280 ;
        RECT 28.160 110.300 28.300 112.360 ;
        RECT 28.560 111.680 28.820 112.000 ;
        RECT 28.620 110.300 28.760 111.680 ;
        RECT 28.100 109.980 28.360 110.300 ;
        RECT 28.560 109.980 28.820 110.300 ;
        RECT 28.560 107.260 28.820 107.580 ;
        RECT 28.100 106.580 28.360 106.900 ;
        RECT 27.640 106.240 27.900 106.560 ;
        RECT 28.160 104.860 28.300 106.580 ;
        RECT 28.100 104.540 28.360 104.860 ;
        RECT 27.180 104.200 27.440 104.520 ;
        RECT 28.620 103.840 28.760 107.260 ;
        RECT 29.020 106.920 29.280 107.240 ;
        RECT 29.080 104.860 29.220 106.920 ;
        RECT 29.020 104.540 29.280 104.860 ;
        RECT 30.920 103.840 31.060 132.760 ;
        RECT 34.080 130.380 34.340 130.700 ;
        RECT 34.140 129.340 34.280 130.380 ;
        RECT 34.080 129.020 34.340 129.340 ;
        RECT 31.320 128.340 31.580 128.660 ;
        RECT 31.380 122.540 31.520 128.340 ;
        RECT 34.600 125.940 34.740 133.530 ;
        RECT 35.000 133.440 35.260 133.760 ;
        RECT 35.060 128.320 35.200 133.440 ;
        RECT 35.000 128.000 35.260 128.320 ;
        RECT 34.540 125.620 34.800 125.940 ;
        RECT 35.060 124.920 35.200 128.000 ;
        RECT 34.540 124.600 34.800 124.920 ;
        RECT 35.000 124.600 35.260 124.920 ;
        RECT 34.600 123.220 34.740 124.600 ;
        RECT 34.540 122.900 34.800 123.220 ;
        RECT 31.320 122.220 31.580 122.540 ;
        RECT 31.380 120.750 31.520 122.220 ;
        RECT 34.600 121.180 34.740 122.900 ;
        RECT 34.540 120.860 34.800 121.180 ;
        RECT 31.780 120.750 32.040 120.840 ;
        RECT 31.380 120.610 32.040 120.750 ;
        RECT 31.780 120.520 32.040 120.610 ;
        RECT 31.840 120.160 31.980 120.520 ;
        RECT 31.780 119.840 32.040 120.160 ;
        RECT 35.060 118.460 35.200 124.600 ;
        RECT 35.000 118.140 35.260 118.460 ;
        RECT 31.320 113.720 31.580 114.040 ;
        RECT 28.560 103.520 28.820 103.840 ;
        RECT 30.860 103.520 31.120 103.840 ;
        RECT 24.940 101.400 26.460 101.540 ;
        RECT 26.320 91.170 26.460 101.400 ;
        RECT 14.290 89.420 14.570 91.170 ;
        RECT 20.270 89.850 20.550 91.170 ;
        RECT 13.920 85.550 15.140 89.420 ;
        RECT 19.910 85.980 21.130 89.850 ;
        RECT 26.250 88.990 26.530 91.170 ;
        RECT 31.380 90.660 31.520 113.720 ;
        RECT 34.080 106.920 34.340 107.240 ;
        RECT 34.140 104.520 34.280 106.920 ;
        RECT 34.080 104.200 34.340 104.520 ;
        RECT 35.520 103.160 35.660 135.480 ;
        RECT 36.380 134.010 36.640 134.100 ;
        RECT 36.900 134.010 37.040 144.320 ;
        RECT 37.300 137.180 37.560 137.500 ;
        RECT 36.380 133.870 37.040 134.010 ;
        RECT 36.380 133.780 36.640 133.870 ;
        RECT 36.900 131.380 37.040 133.870 ;
        RECT 36.840 131.060 37.100 131.380 ;
        RECT 37.360 129.340 37.500 137.180 ;
        RECT 38.280 134.440 38.420 173.900 ;
        RECT 40.120 172.180 40.260 174.580 ;
        RECT 40.060 171.860 40.320 172.180 ;
        RECT 38.680 166.420 38.940 166.740 ;
        RECT 38.740 161.980 38.880 166.420 ;
        RECT 40.060 165.400 40.320 165.720 ;
        RECT 40.120 163.340 40.260 165.400 ;
        RECT 40.060 163.020 40.320 163.340 ;
        RECT 38.680 161.660 38.940 161.980 ;
        RECT 40.060 154.520 40.320 154.840 ;
        RECT 39.600 153.160 39.860 153.480 ;
        RECT 39.660 152.800 39.800 153.160 ;
        RECT 39.600 152.480 39.860 152.800 ;
        RECT 38.680 146.360 38.940 146.680 ;
        RECT 39.600 146.590 39.860 146.680 ;
        RECT 39.200 146.450 39.860 146.590 ;
        RECT 38.220 134.120 38.480 134.440 ;
        RECT 38.740 134.100 38.880 146.360 ;
        RECT 39.200 137.160 39.340 146.450 ;
        RECT 39.600 146.360 39.860 146.450 ;
        RECT 40.120 139.200 40.260 154.520 ;
        RECT 40.060 138.880 40.320 139.200 ;
        RECT 39.600 138.200 39.860 138.520 ;
        RECT 39.660 137.500 39.800 138.200 ;
        RECT 39.600 137.180 39.860 137.500 ;
        RECT 39.140 136.840 39.400 137.160 ;
        RECT 40.060 135.820 40.320 136.140 ;
        RECT 40.120 134.440 40.260 135.820 ;
        RECT 40.060 134.120 40.320 134.440 ;
        RECT 38.680 133.780 38.940 134.100 ;
        RECT 40.580 133.760 40.720 174.920 ;
        RECT 41.500 173.940 41.640 184.440 ;
        RECT 41.960 183.060 42.100 184.440 ;
        RECT 42.880 183.740 43.020 190.900 ;
        RECT 47.940 188.160 48.080 190.900 ;
        RECT 50.700 188.160 50.840 192.600 ;
        RECT 52.480 190.560 52.740 190.880 ;
        RECT 52.540 189.180 52.680 190.560 ;
        RECT 52.480 188.860 52.740 189.180 ;
        RECT 47.880 187.840 48.140 188.160 ;
        RECT 50.640 187.840 50.900 188.160 ;
        RECT 43.280 185.800 43.540 186.120 ;
        RECT 42.820 183.420 43.080 183.740 ;
        RECT 41.900 182.740 42.160 183.060 ;
        RECT 43.340 182.720 43.480 185.800 ;
        RECT 47.940 185.780 48.080 187.840 ;
        RECT 47.880 185.460 48.140 185.780 ;
        RECT 46.040 184.440 46.300 184.760 ;
        RECT 46.100 183.740 46.240 184.440 ;
        RECT 46.040 183.420 46.300 183.740 ;
        RECT 43.280 182.400 43.540 182.720 ;
        RECT 41.900 182.060 42.160 182.380 ;
        RECT 41.960 174.560 42.100 182.060 ;
        RECT 47.940 182.040 48.080 185.460 ;
        RECT 49.720 182.740 49.980 183.060 ;
        RECT 47.880 181.720 48.140 182.040 ;
        RECT 49.780 181.020 49.920 182.740 ;
        RECT 49.720 180.700 49.980 181.020 ;
        RECT 49.260 180.360 49.520 180.680 ;
        RECT 43.740 179.680 44.000 180.000 ;
        RECT 43.280 177.300 43.540 177.620 ;
        RECT 43.340 174.900 43.480 177.300 ;
        RECT 43.280 174.580 43.540 174.900 ;
        RECT 43.800 174.560 43.940 179.680 ;
        RECT 45.580 179.340 45.840 179.660 ;
        RECT 45.640 177.620 45.780 179.340 ;
        RECT 49.320 178.300 49.460 180.360 ;
        RECT 49.260 177.980 49.520 178.300 ;
        RECT 48.340 177.640 48.600 177.960 ;
        RECT 45.580 177.300 45.840 177.620 ;
        RECT 47.420 176.280 47.680 176.600 ;
        RECT 47.880 176.280 48.140 176.600 ;
        RECT 44.660 174.920 44.920 175.240 ;
        RECT 44.720 174.560 44.860 174.920 ;
        RECT 41.900 174.240 42.160 174.560 ;
        RECT 43.740 174.240 44.000 174.560 ;
        RECT 44.660 174.240 44.920 174.560 ;
        RECT 41.040 173.800 41.640 173.940 ;
        RECT 41.040 172.180 41.180 173.800 ;
        RECT 40.980 171.860 41.240 172.180 ;
        RECT 41.440 171.860 41.700 172.180 ;
        RECT 41.500 169.800 41.640 171.860 ;
        RECT 41.440 169.480 41.700 169.800 ;
        RECT 43.280 169.480 43.540 169.800 ;
        RECT 41.440 168.120 41.700 168.440 ;
        RECT 40.980 166.420 41.240 166.740 ;
        RECT 41.040 161.980 41.180 166.420 ;
        RECT 40.980 161.660 41.240 161.980 ;
        RECT 40.980 158.260 41.240 158.580 ;
        RECT 41.040 150.420 41.180 158.260 ;
        RECT 40.980 150.100 41.240 150.420 ;
        RECT 40.980 149.420 41.240 149.740 ;
        RECT 41.040 147.360 41.180 149.420 ;
        RECT 40.980 147.040 41.240 147.360 ;
        RECT 40.980 144.660 41.240 144.980 ;
        RECT 41.040 142.600 41.180 144.660 ;
        RECT 40.980 142.280 41.240 142.600 ;
        RECT 41.500 139.880 41.640 168.120 ;
        RECT 41.900 165.400 42.160 165.720 ;
        RECT 41.960 164.020 42.100 165.400 ;
        RECT 41.900 163.700 42.160 164.020 ;
        RECT 42.360 157.920 42.620 158.240 ;
        RECT 41.900 157.580 42.160 157.900 ;
        RECT 41.960 155.860 42.100 157.580 ;
        RECT 42.420 155.860 42.560 157.920 ;
        RECT 42.820 157.240 43.080 157.560 ;
        RECT 42.880 156.200 43.020 157.240 ;
        RECT 42.820 155.880 43.080 156.200 ;
        RECT 43.340 155.860 43.480 169.480 ;
        RECT 44.720 169.120 44.860 174.240 ;
        RECT 46.040 173.900 46.300 174.220 ;
        RECT 46.500 173.900 46.760 174.220 ;
        RECT 44.660 168.800 44.920 169.120 ;
        RECT 45.580 165.740 45.840 166.060 ;
        RECT 45.640 164.020 45.780 165.740 ;
        RECT 45.580 163.700 45.840 164.020 ;
        RECT 43.740 163.020 44.000 163.340 ;
        RECT 43.800 158.240 43.940 163.020 ;
        RECT 45.580 162.680 45.840 163.000 ;
        RECT 45.640 161.300 45.780 162.680 ;
        RECT 45.580 160.980 45.840 161.300 ;
        RECT 43.740 157.920 44.000 158.240 ;
        RECT 45.120 157.240 45.380 157.560 ;
        RECT 45.580 157.240 45.840 157.560 ;
        RECT 45.180 155.860 45.320 157.240 ;
        RECT 41.900 155.540 42.160 155.860 ;
        RECT 42.360 155.540 42.620 155.860 ;
        RECT 43.280 155.540 43.540 155.860 ;
        RECT 45.120 155.540 45.380 155.860 ;
        RECT 43.740 154.520 44.000 154.840 ;
        RECT 42.820 153.500 43.080 153.820 ;
        RECT 42.360 153.160 42.620 153.480 ;
        RECT 41.900 152.480 42.160 152.800 ;
        RECT 41.960 148.380 42.100 152.480 ;
        RECT 42.420 150.420 42.560 153.160 ;
        RECT 42.880 153.140 43.020 153.500 ;
        RECT 42.820 152.820 43.080 153.140 ;
        RECT 42.880 150.420 43.020 152.820 ;
        RECT 42.360 150.100 42.620 150.420 ;
        RECT 42.820 150.100 43.080 150.420 ;
        RECT 41.900 148.060 42.160 148.380 ;
        RECT 42.420 148.040 42.560 150.100 ;
        RECT 42.360 147.720 42.620 148.040 ;
        RECT 41.440 139.560 41.700 139.880 ;
        RECT 41.440 138.540 41.700 138.860 ;
        RECT 41.500 136.480 41.640 138.540 ;
        RECT 41.440 136.160 41.700 136.480 ;
        RECT 40.520 133.440 40.780 133.760 ;
        RECT 40.980 133.100 41.240 133.420 ;
        RECT 39.140 132.760 39.400 133.080 ;
        RECT 37.300 129.020 37.560 129.340 ;
        RECT 38.220 128.340 38.480 128.660 ;
        RECT 37.760 125.620 38.020 125.940 ;
        RECT 36.830 124.405 37.110 124.775 ;
        RECT 37.300 124.600 37.560 124.920 ;
        RECT 36.900 123.560 37.040 124.405 ;
        RECT 36.840 123.240 37.100 123.560 ;
        RECT 35.920 117.120 36.180 117.440 ;
        RECT 35.980 113.020 36.120 117.120 ;
        RECT 35.920 112.700 36.180 113.020 ;
        RECT 37.360 112.340 37.500 124.600 ;
        RECT 37.820 122.880 37.960 125.620 ;
        RECT 38.280 125.600 38.420 128.340 ;
        RECT 39.200 125.600 39.340 132.760 ;
        RECT 41.040 131.040 41.180 133.100 ;
        RECT 41.500 132.060 41.640 136.160 ;
        RECT 42.360 135.480 42.620 135.800 ;
        RECT 41.440 131.740 41.700 132.060 ;
        RECT 40.520 130.720 40.780 131.040 ;
        RECT 40.980 130.720 41.240 131.040 ;
        RECT 38.220 125.280 38.480 125.600 ;
        RECT 39.140 125.280 39.400 125.600 ;
        RECT 39.600 125.280 39.860 125.600 ;
        RECT 39.660 124.830 39.800 125.280 ;
        RECT 39.200 124.690 39.800 124.830 ;
        RECT 39.200 122.880 39.340 124.690 ;
        RECT 37.760 122.560 38.020 122.880 ;
        RECT 39.140 122.560 39.400 122.880 ;
        RECT 37.820 121.180 37.960 122.560 ;
        RECT 37.760 120.860 38.020 121.180 ;
        RECT 39.200 119.480 39.340 122.560 ;
        RECT 40.580 120.500 40.720 130.720 ;
        RECT 41.500 128.660 41.640 131.740 ;
        RECT 41.440 128.340 41.700 128.660 ;
        RECT 41.440 121.880 41.700 122.200 ;
        RECT 40.520 120.180 40.780 120.500 ;
        RECT 39.600 119.840 39.860 120.160 ;
        RECT 39.140 119.160 39.400 119.480 ;
        RECT 39.200 118.460 39.340 119.160 ;
        RECT 39.140 118.140 39.400 118.460 ;
        RECT 38.220 117.460 38.480 117.780 ;
        RECT 37.300 112.020 37.560 112.340 ;
        RECT 38.280 109.280 38.420 117.460 ;
        RECT 39.660 115.740 39.800 119.840 ;
        RECT 40.580 117.780 40.720 120.180 ;
        RECT 40.520 117.460 40.780 117.780 ;
        RECT 39.600 115.420 39.860 115.740 ;
        RECT 41.500 114.720 41.640 121.880 ;
        RECT 41.440 114.400 41.700 114.720 ;
        RECT 38.220 108.960 38.480 109.280 ;
        RECT 37.760 108.280 38.020 108.600 ;
        RECT 35.460 102.840 35.720 103.160 ;
        RECT 37.820 100.180 37.960 108.280 ;
        RECT 38.280 106.560 38.420 108.960 ;
        RECT 39.600 106.580 39.860 106.900 ;
        RECT 38.220 106.240 38.480 106.560 ;
        RECT 39.660 106.220 39.800 106.580 ;
        RECT 40.520 106.240 40.780 106.560 ;
        RECT 39.600 105.900 39.860 106.220 ;
        RECT 38.680 103.180 38.940 103.500 ;
        RECT 39.140 103.180 39.400 103.500 ;
        RECT 38.740 102.140 38.880 103.180 ;
        RECT 39.200 102.140 39.340 103.180 ;
        RECT 38.680 101.820 38.940 102.140 ;
        RECT 39.140 101.820 39.400 102.140 ;
        RECT 39.660 101.460 39.800 105.900 ;
        RECT 40.580 103.840 40.720 106.240 ;
        RECT 41.440 105.560 41.700 105.880 ;
        RECT 40.980 103.860 41.240 104.180 ;
        RECT 40.520 103.520 40.780 103.840 ;
        RECT 41.040 101.800 41.180 103.860 ;
        RECT 41.500 103.500 41.640 105.560 ;
        RECT 41.440 103.180 41.700 103.500 ;
        RECT 40.980 101.480 41.240 101.800 ;
        RECT 42.420 101.460 42.560 135.480 ;
        RECT 43.800 134.100 43.940 154.520 ;
        RECT 44.660 149.080 44.920 149.400 ;
        RECT 44.200 137.180 44.460 137.500 ;
        RECT 43.740 133.780 44.000 134.100 ;
        RECT 43.280 132.760 43.540 133.080 ;
        RECT 42.820 125.620 43.080 125.940 ;
        RECT 42.880 120.160 43.020 125.620 ;
        RECT 43.340 125.260 43.480 132.760 ;
        RECT 43.280 124.940 43.540 125.260 ;
        RECT 44.260 124.920 44.400 137.180 ;
        RECT 44.720 136.480 44.860 149.080 ;
        RECT 45.640 139.540 45.780 157.240 ;
        RECT 45.580 139.220 45.840 139.540 ;
        RECT 46.100 139.200 46.240 173.900 ;
        RECT 46.560 150.420 46.700 173.900 ;
        RECT 46.960 165.400 47.220 165.720 ;
        RECT 47.020 163.680 47.160 165.400 ;
        RECT 46.960 163.360 47.220 163.680 ;
        RECT 47.480 160.140 47.620 176.280 ;
        RECT 47.020 160.000 47.620 160.140 ;
        RECT 46.500 150.100 46.760 150.420 ;
        RECT 47.020 148.460 47.160 160.000 ;
        RECT 47.420 157.240 47.680 157.560 ;
        RECT 47.480 150.420 47.620 157.240 ;
        RECT 47.420 150.100 47.680 150.420 ;
        RECT 47.420 149.080 47.680 149.400 ;
        RECT 46.560 148.320 47.160 148.460 ;
        RECT 46.040 138.880 46.300 139.200 ;
        RECT 45.580 138.200 45.840 138.520 ;
        RECT 44.660 136.160 44.920 136.480 ;
        RECT 44.660 132.760 44.920 133.080 ;
        RECT 44.200 124.600 44.460 124.920 ;
        RECT 42.820 119.840 43.080 120.160 ;
        RECT 43.280 117.800 43.540 118.120 ;
        RECT 43.340 115.060 43.480 117.800 ;
        RECT 43.280 114.740 43.540 115.060 ;
        RECT 42.820 114.060 43.080 114.380 ;
        RECT 42.880 110.300 43.020 114.060 ;
        RECT 42.820 109.980 43.080 110.300 ;
        RECT 44.720 109.620 44.860 132.760 ;
        RECT 45.640 125.600 45.780 138.200 ;
        RECT 46.560 136.820 46.700 148.320 ;
        RECT 46.960 142.620 47.220 142.940 ;
        RECT 46.500 136.500 46.760 136.820 ;
        RECT 46.040 135.820 46.300 136.140 ;
        RECT 46.100 134.780 46.240 135.820 ;
        RECT 46.040 134.460 46.300 134.780 ;
        RECT 47.020 132.060 47.160 142.620 ;
        RECT 46.960 131.740 47.220 132.060 ;
        RECT 46.960 130.720 47.220 131.040 ;
        RECT 47.020 128.660 47.160 130.720 ;
        RECT 47.480 129.340 47.620 149.080 ;
        RECT 47.940 142.260 48.080 176.280 ;
        RECT 48.400 174.560 48.540 177.640 ;
        RECT 49.320 177.620 49.460 177.980 ;
        RECT 50.700 177.620 50.840 187.840 ;
        RECT 53.000 180.340 53.140 192.600 ;
        RECT 54.320 189.880 54.580 190.200 ;
        RECT 54.780 189.880 55.040 190.200 ;
        RECT 54.380 181.950 54.520 189.880 ;
        RECT 54.840 188.840 54.980 189.880 ;
        RECT 54.780 188.520 55.040 188.840 ;
        RECT 55.300 185.780 55.440 196.000 ;
        RECT 56.620 195.320 56.880 195.640 ;
        RECT 56.680 194.280 56.820 195.320 ;
        RECT 56.620 193.960 56.880 194.280 ;
        RECT 58.920 193.960 59.180 194.280 ;
        RECT 58.980 191.900 59.120 193.960 ;
        RECT 60.360 193.600 60.500 201.440 ;
        RECT 61.740 200.060 61.880 201.780 ;
        RECT 65.420 201.420 65.560 203.480 ;
        RECT 65.360 201.100 65.620 201.420 ;
        RECT 69.100 201.080 69.240 203.480 ;
        RECT 70.420 201.100 70.680 201.420 ;
        RECT 69.040 200.760 69.300 201.080 ;
        RECT 69.100 200.060 69.240 200.760 ;
        RECT 61.680 199.740 61.940 200.060 ;
        RECT 69.040 199.740 69.300 200.060 ;
        RECT 70.480 199.380 70.620 201.100 ;
        RECT 66.740 199.060 67.000 199.380 ;
        RECT 70.420 199.060 70.680 199.380 ;
        RECT 66.800 197.340 66.940 199.060 ;
        RECT 70.480 198.700 70.620 199.060 ;
        RECT 70.420 198.380 70.680 198.700 ;
        RECT 67.660 198.040 67.920 198.360 ;
        RECT 70.880 198.040 71.140 198.360 ;
        RECT 66.740 197.020 67.000 197.340 ;
        RECT 66.740 193.620 67.000 193.940 ;
        RECT 60.300 193.280 60.560 193.600 ;
        RECT 63.980 193.280 64.240 193.600 ;
        RECT 58.920 191.580 59.180 191.900 ;
        RECT 64.040 190.540 64.180 193.280 ;
        RECT 66.280 192.600 66.540 192.920 ;
        RECT 66.340 190.540 66.480 192.600 ;
        RECT 63.980 190.220 64.240 190.540 ;
        RECT 66.280 190.220 66.540 190.540 ;
        RECT 55.240 185.460 55.500 185.780 ;
        RECT 55.300 183.060 55.440 185.460 ;
        RECT 64.040 185.440 64.180 190.220 ;
        RECT 63.980 185.120 64.240 185.440 ;
        RECT 61.680 184.780 61.940 185.100 ;
        RECT 61.740 183.740 61.880 184.780 ;
        RECT 61.680 183.420 61.940 183.740 ;
        RECT 55.240 182.740 55.500 183.060 ;
        RECT 56.620 182.740 56.880 183.060 ;
        RECT 56.160 182.060 56.420 182.380 ;
        RECT 54.380 181.810 54.980 181.950 ;
        RECT 54.320 180.700 54.580 181.020 ;
        RECT 52.940 180.250 53.200 180.340 ;
        RECT 52.940 180.110 54.060 180.250 ;
        RECT 52.940 180.020 53.200 180.110 ;
        RECT 52.940 177.980 53.200 178.300 ;
        RECT 53.000 177.620 53.140 177.980 ;
        RECT 53.920 177.620 54.060 180.110 ;
        RECT 54.380 180.000 54.520 180.700 ;
        RECT 54.320 179.680 54.580 180.000 ;
        RECT 54.380 178.300 54.520 179.680 ;
        RECT 54.840 179.320 54.980 181.810 ;
        RECT 55.700 181.720 55.960 182.040 ;
        RECT 55.760 179.660 55.900 181.720 ;
        RECT 55.700 179.340 55.960 179.660 ;
        RECT 54.780 179.000 55.040 179.320 ;
        RECT 54.320 177.980 54.580 178.300 ;
        RECT 49.260 177.300 49.520 177.620 ;
        RECT 50.640 177.300 50.900 177.620 ;
        RECT 52.940 177.300 53.200 177.620 ;
        RECT 53.860 177.300 54.120 177.620 ;
        RECT 49.320 175.240 49.460 177.300 ;
        RECT 49.720 176.280 49.980 176.600 ;
        RECT 49.260 174.920 49.520 175.240 ;
        RECT 48.340 174.240 48.600 174.560 ;
        RECT 48.400 173.880 48.540 174.240 ;
        RECT 48.340 173.560 48.600 173.880 ;
        RECT 48.400 168.780 48.540 173.560 ;
        RECT 48.340 168.460 48.600 168.780 ;
        RECT 48.800 165.400 49.060 165.720 ;
        RECT 48.860 160.620 49.000 165.400 ;
        RECT 48.800 160.300 49.060 160.620 ;
        RECT 48.860 158.240 49.000 160.300 ;
        RECT 49.260 158.600 49.520 158.920 ;
        RECT 49.320 158.240 49.460 158.600 ;
        RECT 48.340 157.920 48.600 158.240 ;
        RECT 48.800 157.920 49.060 158.240 ;
        RECT 49.260 157.920 49.520 158.240 ;
        RECT 48.400 155.770 48.540 157.920 ;
        RECT 48.800 155.770 49.060 155.860 ;
        RECT 48.400 155.630 49.060 155.770 ;
        RECT 48.800 155.540 49.060 155.630 ;
        RECT 49.320 155.180 49.460 157.920 ;
        RECT 49.260 154.860 49.520 155.180 ;
        RECT 49.780 150.420 49.920 176.280 ;
        RECT 52.480 174.240 52.740 174.560 ;
        RECT 52.540 172.860 52.680 174.240 ;
        RECT 54.840 174.220 54.980 179.000 ;
        RECT 55.240 177.300 55.500 177.620 ;
        RECT 55.300 175.580 55.440 177.300 ;
        RECT 56.220 177.280 56.360 182.060 ;
        RECT 56.160 176.960 56.420 177.280 ;
        RECT 55.240 175.260 55.500 175.580 ;
        RECT 56.220 174.900 56.360 176.960 ;
        RECT 56.160 174.580 56.420 174.900 ;
        RECT 54.780 173.900 55.040 174.220 ;
        RECT 52.480 172.540 52.740 172.860 ;
        RECT 53.400 171.860 53.660 172.180 ;
        RECT 53.460 171.695 53.600 171.860 ;
        RECT 53.390 171.325 53.670 171.695 ;
        RECT 56.680 170.140 56.820 182.740 ;
        RECT 57.080 182.400 57.340 182.720 ;
        RECT 57.140 176.940 57.280 182.400 ;
        RECT 61.220 181.720 61.480 182.040 ;
        RECT 61.280 179.660 61.420 181.720 ;
        RECT 64.040 180.000 64.180 185.120 ;
        RECT 65.820 182.400 66.080 182.720 ;
        RECT 65.880 180.000 66.020 182.400 ;
        RECT 63.980 179.680 64.240 180.000 ;
        RECT 65.820 179.680 66.080 180.000 ;
        RECT 61.220 179.340 61.480 179.660 ;
        RECT 58.000 177.300 58.260 177.620 ;
        RECT 57.080 176.620 57.340 176.940 ;
        RECT 57.530 176.765 57.810 177.135 ;
        RECT 57.600 176.600 57.740 176.765 ;
        RECT 57.540 176.280 57.800 176.600 ;
        RECT 58.060 174.560 58.200 177.300 ;
        RECT 59.840 176.280 60.100 176.600 ;
        RECT 59.900 174.900 60.040 176.280 ;
        RECT 59.840 174.580 60.100 174.900 ;
        RECT 58.000 174.240 58.260 174.560 ;
        RECT 61.220 173.560 61.480 173.880 ;
        RECT 61.280 172.520 61.420 173.560 ;
        RECT 61.220 172.200 61.480 172.520 ;
        RECT 64.040 171.840 64.180 179.680 ;
        RECT 66.270 179.485 66.550 179.855 ;
        RECT 66.280 179.340 66.540 179.485 ;
        RECT 65.360 179.000 65.620 179.320 ;
        RECT 65.420 177.815 65.560 179.000 ;
        RECT 65.350 177.445 65.630 177.815 ;
        RECT 66.340 176.940 66.480 179.340 ;
        RECT 66.280 176.620 66.540 176.940 ;
        RECT 64.440 176.280 64.700 176.600 ;
        RECT 64.500 175.240 64.640 176.280 ;
        RECT 64.440 174.920 64.700 175.240 ;
        RECT 66.800 174.900 66.940 193.620 ;
        RECT 66.740 174.580 67.000 174.900 ;
        RECT 64.440 171.860 64.700 172.180 ;
        RECT 63.980 171.520 64.240 171.840 ;
        RECT 57.540 170.840 57.800 171.160 ;
        RECT 56.620 169.820 56.880 170.140 ;
        RECT 57.600 169.120 57.740 170.840 ;
        RECT 57.540 168.800 57.800 169.120 ;
        RECT 54.320 166.760 54.580 167.080 ;
        RECT 54.380 166.400 54.520 166.760 ;
        RECT 57.600 166.400 57.740 168.800 ;
        RECT 64.040 166.400 64.180 171.520 ;
        RECT 64.500 170.140 64.640 171.860 ;
        RECT 64.440 169.820 64.700 170.140 ;
        RECT 64.500 167.420 64.640 169.820 ;
        RECT 64.900 168.120 65.160 168.440 ;
        RECT 64.440 167.100 64.700 167.420 ;
        RECT 64.440 166.420 64.700 166.740 ;
        RECT 54.320 166.080 54.580 166.400 ;
        RECT 54.780 166.080 55.040 166.400 ;
        RECT 57.540 166.080 57.800 166.400 ;
        RECT 63.980 166.080 64.240 166.400 ;
        RECT 51.100 163.700 51.360 164.020 ;
        RECT 53.860 163.700 54.120 164.020 ;
        RECT 51.160 160.960 51.300 163.700 ;
        RECT 51.560 162.680 51.820 163.000 ;
        RECT 51.620 161.640 51.760 162.680 ;
        RECT 51.560 161.320 51.820 161.640 ;
        RECT 53.920 161.300 54.060 163.700 ;
        RECT 54.320 162.680 54.580 163.000 ;
        RECT 54.380 161.300 54.520 162.680 ;
        RECT 52.940 160.980 53.200 161.300 ;
        RECT 53.860 160.980 54.120 161.300 ;
        RECT 54.320 160.980 54.580 161.300 ;
        RECT 51.100 160.640 51.360 160.960 ;
        RECT 52.020 158.600 52.280 158.920 ;
        RECT 52.080 158.240 52.220 158.600 ;
        RECT 53.000 158.240 53.140 160.980 ;
        RECT 54.840 159.260 54.980 166.080 ;
        RECT 58.460 165.400 58.720 165.720 ;
        RECT 58.520 163.340 58.660 165.400 ;
        RECT 64.040 163.680 64.180 166.080 ;
        RECT 63.980 163.360 64.240 163.680 ;
        RECT 58.460 163.020 58.720 163.340 ;
        RECT 62.140 163.020 62.400 163.340 ;
        RECT 62.200 161.980 62.340 163.020 ;
        RECT 62.140 161.660 62.400 161.980 ;
        RECT 55.700 159.960 55.960 160.280 ;
        RECT 54.780 158.940 55.040 159.260 ;
        RECT 55.760 158.240 55.900 159.960 ;
        RECT 52.020 157.920 52.280 158.240 ;
        RECT 52.940 157.920 53.200 158.240 ;
        RECT 55.700 157.920 55.960 158.240 ;
        RECT 57.080 157.920 57.340 158.240 ;
        RECT 63.520 157.920 63.780 158.240 ;
        RECT 52.080 157.560 52.220 157.920 ;
        RECT 50.180 157.240 50.440 157.560 ;
        RECT 52.020 157.240 52.280 157.560 ;
        RECT 50.240 150.420 50.380 157.240 ;
        RECT 52.080 155.860 52.220 157.240 ;
        RECT 52.020 155.540 52.280 155.860 ;
        RECT 50.640 154.520 50.900 154.840 ;
        RECT 53.860 154.520 54.120 154.840 ;
        RECT 48.800 150.100 49.060 150.420 ;
        RECT 49.720 150.100 49.980 150.420 ;
        RECT 50.180 150.100 50.440 150.420 ;
        RECT 48.340 149.080 48.600 149.400 ;
        RECT 47.880 141.940 48.140 142.260 ;
        RECT 47.880 136.160 48.140 136.480 ;
        RECT 47.940 134.780 48.080 136.160 ;
        RECT 47.880 134.460 48.140 134.780 ;
        RECT 48.400 130.700 48.540 149.080 ;
        RECT 48.860 148.380 49.000 150.100 ;
        RECT 48.800 148.060 49.060 148.380 ;
        RECT 50.180 141.940 50.440 142.260 ;
        RECT 48.800 139.900 49.060 140.220 ;
        RECT 48.860 139.540 49.000 139.900 ;
        RECT 48.800 139.220 49.060 139.540 ;
        RECT 49.720 139.110 49.980 139.200 ;
        RECT 50.240 139.110 50.380 141.940 ;
        RECT 50.700 141.920 50.840 154.520 ;
        RECT 51.560 152.480 51.820 152.800 ;
        RECT 51.100 150.100 51.360 150.420 ;
        RECT 51.160 142.260 51.300 150.100 ;
        RECT 51.620 145.320 51.760 152.480 ;
        RECT 53.400 150.780 53.660 151.100 ;
        RECT 52.020 149.080 52.280 149.400 ;
        RECT 51.560 145.000 51.820 145.320 ;
        RECT 51.620 142.940 51.760 145.000 ;
        RECT 51.560 142.620 51.820 142.940 ;
        RECT 51.100 141.940 51.360 142.260 ;
        RECT 50.640 141.600 50.900 141.920 ;
        RECT 51.100 140.920 51.360 141.240 ;
        RECT 51.560 140.920 51.820 141.240 ;
        RECT 51.160 140.220 51.300 140.920 ;
        RECT 50.640 139.900 50.900 140.220 ;
        RECT 51.100 139.900 51.360 140.220 ;
        RECT 49.720 138.970 50.380 139.110 ;
        RECT 49.720 138.880 49.980 138.970 ;
        RECT 48.800 138.540 49.060 138.860 ;
        RECT 48.860 134.100 49.000 138.540 ;
        RECT 49.780 134.100 49.920 138.880 ;
        RECT 48.800 133.780 49.060 134.100 ;
        RECT 49.720 133.780 49.980 134.100 ;
        RECT 49.780 133.080 49.920 133.780 ;
        RECT 49.720 132.760 49.980 133.080 ;
        RECT 48.340 130.380 48.600 130.700 ;
        RECT 47.420 129.020 47.680 129.340 ;
        RECT 46.960 128.340 47.220 128.660 ;
        RECT 45.580 125.280 45.840 125.600 ;
        RECT 46.500 125.510 46.760 125.600 ;
        RECT 47.020 125.510 47.160 128.340 ;
        RECT 46.500 125.370 47.160 125.510 ;
        RECT 46.500 125.280 46.760 125.370 ;
        RECT 47.880 125.280 48.140 125.600 ;
        RECT 46.500 124.600 46.760 124.920 ;
        RECT 45.580 122.220 45.840 122.540 ;
        RECT 45.120 117.460 45.380 117.780 ;
        RECT 45.180 115.740 45.320 117.460 ;
        RECT 45.120 115.420 45.380 115.740 ;
        RECT 45.640 114.720 45.780 122.220 ;
        RECT 46.560 120.500 46.700 124.600 ;
        RECT 46.500 120.180 46.760 120.500 ;
        RECT 47.940 119.820 48.080 125.280 ;
        RECT 50.180 122.220 50.440 122.540 ;
        RECT 50.240 120.160 50.380 122.220 ;
        RECT 50.180 119.840 50.440 120.160 ;
        RECT 47.880 119.500 48.140 119.820 ;
        RECT 47.940 118.460 48.080 119.500 ;
        RECT 48.800 119.160 49.060 119.480 ;
        RECT 49.720 119.160 49.980 119.480 ;
        RECT 47.880 118.140 48.140 118.460 ;
        RECT 48.860 114.720 49.000 119.160 ;
        RECT 49.780 114.720 49.920 119.160 ;
        RECT 45.580 114.400 45.840 114.720 ;
        RECT 48.800 114.400 49.060 114.720 ;
        RECT 49.720 114.400 49.980 114.720 ;
        RECT 44.660 109.300 44.920 109.620 ;
        RECT 50.700 109.280 50.840 139.900 ;
        RECT 51.620 139.540 51.760 140.920 ;
        RECT 51.560 139.220 51.820 139.540 ;
        RECT 51.620 133.500 51.760 139.220 ;
        RECT 51.160 133.420 51.760 133.500 ;
        RECT 51.100 133.360 51.760 133.420 ;
        RECT 51.100 133.100 51.360 133.360 ;
        RECT 51.100 124.940 51.360 125.260 ;
        RECT 51.160 124.775 51.300 124.940 ;
        RECT 51.090 124.405 51.370 124.775 ;
        RECT 51.100 119.160 51.360 119.480 ;
        RECT 51.160 118.120 51.300 119.160 ;
        RECT 51.100 117.800 51.360 118.120 ;
        RECT 52.080 109.620 52.220 149.080 ;
        RECT 52.480 146.700 52.740 147.020 ;
        RECT 52.540 143.960 52.680 146.700 ;
        RECT 52.940 146.360 53.200 146.680 ;
        RECT 53.000 144.980 53.140 146.360 ;
        RECT 52.940 144.660 53.200 144.980 ;
        RECT 53.460 144.380 53.600 150.780 ;
        RECT 53.920 150.420 54.060 154.520 ;
        RECT 57.140 152.800 57.280 157.920 ;
        RECT 63.580 155.860 63.720 157.920 ;
        RECT 60.300 155.540 60.560 155.860 ;
        RECT 63.520 155.540 63.780 155.860 ;
        RECT 60.360 153.480 60.500 155.540 ;
        RECT 64.040 155.520 64.180 163.360 ;
        RECT 64.500 158.240 64.640 166.420 ;
        RECT 64.440 157.920 64.700 158.240 ;
        RECT 64.500 156.540 64.640 157.920 ;
        RECT 64.440 156.220 64.700 156.540 ;
        RECT 60.760 155.200 61.020 155.520 ;
        RECT 63.980 155.200 64.240 155.520 ;
        RECT 60.300 153.160 60.560 153.480 ;
        RECT 57.080 152.480 57.340 152.800 ;
        RECT 59.840 152.030 60.100 152.120 ;
        RECT 59.840 151.890 60.500 152.030 ;
        RECT 59.840 151.800 60.100 151.890 ;
        RECT 60.360 150.500 60.500 151.890 ;
        RECT 60.820 151.100 60.960 155.200 ;
        RECT 64.040 153.140 64.180 155.200 ;
        RECT 63.980 152.820 64.240 153.140 ;
        RECT 60.760 150.780 61.020 151.100 ;
        RECT 59.440 150.420 60.500 150.500 ;
        RECT 53.860 150.100 54.120 150.420 ;
        RECT 54.780 150.100 55.040 150.420 ;
        RECT 59.380 150.360 60.500 150.420 ;
        RECT 59.380 150.100 59.640 150.360 ;
        RECT 63.980 150.100 64.240 150.420 ;
        RECT 53.920 147.700 54.060 150.100 ;
        RECT 53.860 147.380 54.120 147.700 ;
        RECT 54.320 147.380 54.580 147.700 ;
        RECT 53.000 144.240 53.600 144.380 ;
        RECT 52.480 143.640 52.740 143.960 ;
        RECT 52.540 139.540 52.680 143.640 ;
        RECT 52.480 139.220 52.740 139.540 ;
        RECT 52.540 136.480 52.680 139.220 ;
        RECT 52.480 136.160 52.740 136.480 ;
        RECT 52.020 109.300 52.280 109.620 ;
        RECT 53.000 109.280 53.140 144.240 ;
        RECT 54.380 136.820 54.520 147.380 ;
        RECT 54.840 147.215 54.980 150.100 ;
        RECT 57.080 149.760 57.340 150.080 ;
        RECT 56.620 149.420 56.880 149.740 ;
        RECT 56.680 147.360 56.820 149.420 ;
        RECT 57.140 148.040 57.280 149.760 ;
        RECT 57.080 147.720 57.340 148.040 ;
        RECT 54.770 146.845 55.050 147.215 ;
        RECT 56.620 147.040 56.880 147.360 ;
        RECT 57.140 147.270 57.280 147.720 ;
        RECT 57.540 147.270 57.800 147.360 ;
        RECT 57.140 147.130 57.800 147.270 ;
        RECT 58.920 147.215 59.180 147.360 ;
        RECT 54.840 141.830 54.980 146.845 ;
        RECT 56.680 145.660 56.820 147.040 ;
        RECT 56.620 145.340 56.880 145.660 ;
        RECT 56.160 145.000 56.420 145.320 ;
        RECT 55.240 141.830 55.500 141.920 ;
        RECT 54.840 141.690 55.500 141.830 ;
        RECT 55.240 141.600 55.500 141.690 ;
        RECT 55.300 138.860 55.440 141.600 ;
        RECT 55.700 139.220 55.960 139.540 ;
        RECT 55.240 138.540 55.500 138.860 ;
        RECT 54.320 136.500 54.580 136.820 ;
        RECT 54.380 136.220 54.520 136.500 ;
        RECT 54.380 136.080 54.980 136.220 ;
        RECT 54.320 135.480 54.580 135.800 ;
        RECT 53.400 134.120 53.660 134.440 ;
        RECT 53.460 129.340 53.600 134.120 ;
        RECT 54.380 133.080 54.520 135.480 ;
        RECT 54.320 132.760 54.580 133.080 ;
        RECT 53.400 129.020 53.660 129.340 ;
        RECT 54.840 128.320 54.980 136.080 ;
        RECT 55.300 134.100 55.440 138.540 ;
        RECT 55.760 134.440 55.900 139.220 ;
        RECT 56.220 139.200 56.360 145.000 ;
        RECT 57.140 141.580 57.280 147.130 ;
        RECT 57.540 147.040 57.800 147.130 ;
        RECT 58.910 146.845 59.190 147.215 ;
        RECT 59.440 147.020 59.580 150.100 ;
        RECT 59.380 146.700 59.640 147.020 ;
        RECT 61.680 146.700 61.940 147.020 ;
        RECT 61.740 145.320 61.880 146.700 ;
        RECT 64.040 146.680 64.180 150.100 ;
        RECT 63.980 146.360 64.240 146.680 ;
        RECT 59.380 145.000 59.640 145.320 ;
        RECT 61.680 145.000 61.940 145.320 ;
        RECT 58.920 143.640 59.180 143.960 ;
        RECT 58.980 141.580 59.120 143.640 ;
        RECT 59.440 142.940 59.580 145.000 ;
        RECT 64.440 144.660 64.700 144.980 ;
        RECT 59.380 142.620 59.640 142.940 ;
        RECT 61.220 141.940 61.480 142.260 ;
        RECT 57.080 141.260 57.340 141.580 ;
        RECT 58.920 141.260 59.180 141.580 ;
        RECT 56.160 138.880 56.420 139.200 ;
        RECT 60.300 135.480 60.560 135.800 ;
        RECT 55.700 134.120 55.960 134.440 ;
        RECT 55.240 133.780 55.500 134.100 ;
        RECT 60.360 133.760 60.500 135.480 ;
        RECT 60.300 133.440 60.560 133.760 ;
        RECT 56.620 132.760 56.880 133.080 ;
        RECT 56.680 129.340 56.820 132.760 ;
        RECT 56.160 129.020 56.420 129.340 ;
        RECT 56.620 129.020 56.880 129.340 ;
        RECT 54.780 128.000 55.040 128.320 ;
        RECT 54.840 126.280 54.980 128.000 ;
        RECT 54.780 125.960 55.040 126.280 ;
        RECT 56.220 125.940 56.360 129.020 ;
        RECT 60.300 127.320 60.560 127.640 ;
        RECT 56.160 125.620 56.420 125.940 ;
        RECT 56.220 123.900 56.360 125.620 ;
        RECT 57.540 124.600 57.800 124.920 ;
        RECT 56.160 123.580 56.420 123.900 ;
        RECT 56.620 123.240 56.880 123.560 ;
        RECT 56.680 118.460 56.820 123.240 ;
        RECT 57.600 122.880 57.740 124.600 ;
        RECT 60.360 123.220 60.500 127.320 ;
        RECT 60.300 122.900 60.560 123.220 ;
        RECT 57.540 122.560 57.800 122.880 ;
        RECT 57.600 119.820 57.740 122.560 ;
        RECT 60.300 119.840 60.560 120.160 ;
        RECT 57.540 119.500 57.800 119.820 ;
        RECT 57.600 118.540 57.740 119.500 ;
        RECT 56.620 118.140 56.880 118.460 ;
        RECT 57.140 118.400 57.740 118.540 ;
        RECT 57.140 117.440 57.280 118.400 ;
        RECT 60.360 117.780 60.500 119.840 ;
        RECT 60.300 117.460 60.560 117.780 ;
        RECT 54.780 117.120 55.040 117.440 ;
        RECT 57.080 117.120 57.340 117.440 ;
        RECT 54.840 115.740 54.980 117.120 ;
        RECT 54.780 115.420 55.040 115.740 ;
        RECT 50.640 108.960 50.900 109.280 ;
        RECT 52.940 108.960 53.200 109.280 ;
        RECT 48.340 108.280 48.600 108.600 ;
        RECT 55.700 108.280 55.960 108.600 ;
        RECT 48.400 104.180 48.540 108.280 ;
        RECT 55.760 107.240 55.900 108.280 ;
        RECT 55.700 106.920 55.960 107.240 ;
        RECT 57.140 106.900 57.280 117.120 ;
        RECT 60.300 114.740 60.560 115.060 ;
        RECT 60.360 109.280 60.500 114.740 ;
        RECT 60.300 108.960 60.560 109.280 ;
        RECT 60.760 108.280 61.020 108.600 ;
        RECT 48.800 106.580 49.060 106.900 ;
        RECT 50.180 106.580 50.440 106.900 ;
        RECT 57.080 106.580 57.340 106.900 ;
        RECT 48.340 103.860 48.600 104.180 ;
        RECT 39.600 101.140 39.860 101.460 ;
        RECT 42.360 101.140 42.620 101.460 ;
        RECT 44.200 100.460 44.460 100.780 ;
        RECT 37.820 100.040 38.420 100.180 ;
        RECT 38.280 91.170 38.420 100.040 ;
        RECT 44.260 91.170 44.400 100.460 ;
        RECT 32.230 90.660 32.510 91.170 ;
        RECT 31.380 90.520 32.510 90.660 ;
        RECT 32.230 89.380 32.510 90.520 ;
        RECT 25.730 85.120 26.950 88.990 ;
        RECT 31.780 85.510 33.000 89.380 ;
        RECT 38.210 89.290 38.490 91.170 ;
        RECT 44.190 89.530 44.470 91.170 ;
        RECT 48.860 90.660 49.000 106.580 ;
        RECT 50.240 104.860 50.380 106.580 ;
        RECT 60.820 106.300 60.960 108.280 ;
        RECT 61.280 106.900 61.420 141.940 ;
        RECT 63.980 139.900 64.240 140.220 ;
        RECT 64.040 137.160 64.180 139.900 ;
        RECT 64.500 139.880 64.640 144.660 ;
        RECT 64.960 140.300 65.100 168.120 ;
        RECT 67.720 166.400 67.860 198.040 ;
        RECT 70.420 197.020 70.680 197.340 ;
        RECT 69.040 192.600 69.300 192.920 ;
        RECT 69.100 191.560 69.240 192.600 ;
        RECT 69.040 191.240 69.300 191.560 ;
        RECT 69.100 188.160 69.240 191.240 ;
        RECT 70.480 190.880 70.620 197.020 ;
        RECT 70.420 190.560 70.680 190.880 ;
        RECT 69.040 187.840 69.300 188.160 ;
        RECT 69.100 182.720 69.240 187.840 ;
        RECT 69.040 182.400 69.300 182.720 ;
        RECT 69.500 182.060 69.760 182.380 ;
        RECT 68.580 180.420 68.840 180.680 ;
        RECT 68.580 180.360 69.240 180.420 ;
        RECT 68.640 180.280 69.240 180.360 ;
        RECT 69.560 180.340 69.700 182.060 ;
        RECT 68.580 179.680 68.840 180.000 ;
        RECT 69.100 179.740 69.240 180.280 ;
        RECT 69.500 180.020 69.760 180.340 ;
        RECT 70.940 180.250 71.080 198.040 ;
        RECT 71.400 194.280 71.540 205.180 ;
        RECT 75.540 202.780 75.680 206.880 ;
        RECT 75.940 206.200 76.200 206.520 ;
        RECT 76.000 205.160 76.140 206.200 ;
        RECT 75.940 204.840 76.200 205.160 ;
        RECT 77.780 203.480 78.040 203.800 ;
        RECT 79.160 203.480 79.420 203.800 ;
        RECT 75.480 202.460 75.740 202.780 ;
        RECT 72.260 201.780 72.520 202.100 ;
        RECT 72.320 200.060 72.460 201.780 ;
        RECT 73.640 201.100 73.900 201.420 ;
        RECT 72.260 199.740 72.520 200.060 ;
        RECT 72.320 199.040 72.460 199.740 ;
        RECT 72.260 198.720 72.520 199.040 ;
        RECT 73.700 196.660 73.840 201.100 ;
        RECT 74.100 199.400 74.360 199.720 ;
        RECT 74.160 198.700 74.300 199.400 ;
        RECT 75.540 198.700 75.680 202.460 ;
        RECT 77.840 202.100 77.980 203.480 ;
        RECT 79.220 202.780 79.360 203.480 ;
        RECT 79.160 202.460 79.420 202.780 ;
        RECT 77.780 201.780 78.040 202.100 ;
        RECT 78.240 201.440 78.500 201.760 ;
        RECT 76.860 201.100 77.120 201.420 ;
        RECT 76.920 200.060 77.060 201.100 ;
        RECT 77.320 200.760 77.580 201.080 ;
        RECT 76.860 199.740 77.120 200.060 ;
        RECT 75.940 199.400 76.200 199.720 ;
        RECT 74.100 198.380 74.360 198.700 ;
        RECT 75.480 198.380 75.740 198.700 ;
        RECT 74.160 196.660 74.300 198.380 ;
        RECT 73.180 196.340 73.440 196.660 ;
        RECT 73.640 196.340 73.900 196.660 ;
        RECT 74.100 196.340 74.360 196.660 ;
        RECT 73.240 195.640 73.380 196.340 ;
        RECT 73.180 195.320 73.440 195.640 ;
        RECT 71.340 193.960 71.600 194.280 ;
        RECT 73.700 193.940 73.840 196.340 ;
        RECT 74.160 193.940 74.300 196.340 ;
        RECT 75.540 196.320 75.680 198.380 ;
        RECT 75.480 196.000 75.740 196.320 ;
        RECT 74.560 195.320 74.820 195.640 ;
        RECT 73.640 193.620 73.900 193.940 ;
        RECT 74.100 193.620 74.360 193.940 ;
        RECT 73.180 190.560 73.440 190.880 ;
        RECT 73.240 189.180 73.380 190.560 ;
        RECT 73.180 188.860 73.440 189.180 ;
        RECT 74.160 188.070 74.300 193.620 ;
        RECT 74.620 193.600 74.760 195.320 ;
        RECT 74.560 193.280 74.820 193.600 ;
        RECT 75.540 192.920 75.680 196.000 ;
        RECT 76.000 195.980 76.140 199.400 ;
        RECT 77.380 198.700 77.520 200.760 ;
        RECT 78.300 200.060 78.440 201.440 ;
        RECT 78.700 200.760 78.960 201.080 ;
        RECT 78.240 199.740 78.500 200.060 ;
        RECT 78.760 199.380 78.900 200.760 ;
        RECT 81.060 199.720 81.200 207.220 ;
        RECT 88.360 204.160 88.620 204.480 ;
        RECT 88.420 202.100 88.560 204.160 ;
        RECT 84.680 201.780 84.940 202.100 ;
        RECT 88.360 201.780 88.620 202.100 ;
        RECT 83.300 201.100 83.560 201.420 ;
        RECT 83.360 200.060 83.500 201.100 ;
        RECT 84.740 200.060 84.880 201.780 ;
        RECT 88.420 201.330 88.560 201.780 ;
        RECT 87.500 201.190 88.560 201.330 ;
        RECT 83.300 199.740 83.560 200.060 ;
        RECT 84.680 199.740 84.940 200.060 ;
        RECT 81.000 199.400 81.260 199.720 ;
        RECT 78.700 199.060 78.960 199.380 ;
        RECT 83.760 199.060 84.020 199.380 ;
        RECT 77.780 198.720 78.040 199.040 ;
        RECT 77.320 198.380 77.580 198.700 ;
        RECT 76.400 196.680 76.660 197.000 ;
        RECT 75.940 195.660 76.200 195.980 ;
        RECT 76.000 194.620 76.140 195.660 ;
        RECT 75.940 194.300 76.200 194.620 ;
        RECT 75.940 193.280 76.200 193.600 ;
        RECT 75.480 192.600 75.740 192.920 ;
        RECT 75.540 190.880 75.680 192.600 ;
        RECT 75.480 190.790 75.740 190.880 ;
        RECT 73.700 187.930 74.300 188.070 ;
        RECT 75.080 190.650 75.740 190.790 ;
        RECT 73.700 183.060 73.840 187.930 ;
        RECT 75.080 183.060 75.220 190.650 ;
        RECT 75.480 190.560 75.740 190.650 ;
        RECT 76.000 190.200 76.140 193.280 ;
        RECT 76.460 191.220 76.600 196.680 ;
        RECT 77.380 195.980 77.520 198.380 ;
        RECT 77.840 197.000 77.980 198.720 ;
        RECT 80.080 198.040 80.340 198.360 ;
        RECT 80.140 197.340 80.280 198.040 ;
        RECT 80.080 197.020 80.340 197.340 ;
        RECT 77.780 196.680 78.040 197.000 ;
        RECT 77.840 196.320 77.980 196.680 ;
        RECT 77.780 196.000 78.040 196.320 ;
        RECT 77.320 195.660 77.580 195.980 ;
        RECT 83.820 194.620 83.960 199.060 ;
        RECT 83.760 194.300 84.020 194.620 ;
        RECT 77.320 193.620 77.580 193.940 ;
        RECT 84.680 193.620 84.940 193.940 ;
        RECT 86.520 193.620 86.780 193.940 ;
        RECT 77.380 191.220 77.520 193.620 ;
        RECT 76.400 190.900 76.660 191.220 ;
        RECT 77.320 190.900 77.580 191.220 ;
        RECT 75.940 189.880 76.200 190.200 ;
        RECT 75.480 183.080 75.740 183.400 ;
        RECT 73.640 182.740 73.900 183.060 ;
        RECT 75.020 182.740 75.280 183.060 ;
        RECT 71.340 182.060 71.600 182.380 ;
        RECT 70.480 180.110 71.080 180.250 ;
        RECT 68.120 179.000 68.380 179.320 ;
        RECT 68.180 177.620 68.320 179.000 ;
        RECT 68.120 177.300 68.380 177.620 ;
        RECT 68.640 167.080 68.780 179.680 ;
        RECT 69.100 179.600 69.700 179.740 ;
        RECT 69.960 179.680 70.220 180.000 ;
        RECT 69.030 177.445 69.310 177.815 ;
        RECT 69.040 177.300 69.300 177.445 ;
        RECT 69.040 176.620 69.300 176.940 ;
        RECT 69.100 175.660 69.240 176.620 ;
        RECT 69.560 176.340 69.700 179.600 ;
        RECT 70.020 177.815 70.160 179.680 ;
        RECT 69.950 177.445 70.230 177.815 ;
        RECT 69.560 176.200 70.160 176.340 ;
        RECT 69.100 175.520 69.700 175.660 ;
        RECT 69.040 173.900 69.300 174.220 ;
        RECT 69.100 172.180 69.240 173.900 ;
        RECT 69.040 171.860 69.300 172.180 ;
        RECT 68.580 166.760 68.840 167.080 ;
        RECT 67.660 166.080 67.920 166.400 ;
        RECT 67.720 161.640 67.860 166.080 ;
        RECT 69.100 165.720 69.240 171.860 ;
        RECT 69.560 166.060 69.700 175.520 ;
        RECT 70.020 175.240 70.160 176.200 ;
        RECT 69.960 174.920 70.220 175.240 ;
        RECT 69.960 166.420 70.220 166.740 ;
        RECT 69.500 165.740 69.760 166.060 ;
        RECT 69.040 165.400 69.300 165.720 ;
        RECT 67.660 161.320 67.920 161.640 ;
        RECT 65.360 159.960 65.620 160.280 ;
        RECT 66.280 159.960 66.540 160.280 ;
        RECT 65.420 158.580 65.560 159.960 ;
        RECT 65.360 158.260 65.620 158.580 ;
        RECT 66.340 153.820 66.480 159.960 ;
        RECT 66.740 155.375 67.000 155.520 ;
        RECT 66.730 155.005 67.010 155.375 ;
        RECT 67.200 154.520 67.460 154.840 ;
        RECT 66.280 153.500 66.540 153.820 ;
        RECT 65.820 152.820 66.080 153.140 ;
        RECT 65.880 151.100 66.020 152.820 ;
        RECT 65.820 150.780 66.080 151.100 ;
        RECT 65.360 149.420 65.620 149.740 ;
        RECT 65.420 147.700 65.560 149.420 ;
        RECT 67.260 148.380 67.400 154.520 ;
        RECT 67.660 153.160 67.920 153.480 ;
        RECT 67.720 150.420 67.860 153.160 ;
        RECT 68.120 151.800 68.380 152.120 ;
        RECT 67.660 150.100 67.920 150.420 ;
        RECT 67.200 148.060 67.460 148.380 ;
        RECT 65.360 147.380 65.620 147.700 ;
        RECT 65.420 144.640 65.560 147.380 ;
        RECT 65.360 144.320 65.620 144.640 ;
        RECT 64.960 140.160 66.020 140.300 ;
        RECT 64.960 139.880 65.100 140.160 ;
        RECT 64.440 139.560 64.700 139.880 ;
        RECT 64.900 139.560 65.160 139.880 ;
        RECT 64.500 138.520 64.640 139.560 ;
        RECT 65.360 139.220 65.620 139.540 ;
        RECT 64.900 138.880 65.160 139.200 ;
        RECT 64.440 138.200 64.700 138.520 ;
        RECT 63.980 136.840 64.240 137.160 ;
        RECT 63.980 136.160 64.240 136.480 ;
        RECT 62.600 124.940 62.860 125.260 ;
        RECT 62.660 122.540 62.800 124.940 ;
        RECT 63.520 124.830 63.780 124.920 ;
        RECT 64.040 124.830 64.180 136.160 ;
        RECT 64.960 136.140 65.100 138.880 ;
        RECT 65.420 138.860 65.560 139.220 ;
        RECT 65.360 138.540 65.620 138.860 ;
        RECT 65.420 137.500 65.560 138.540 ;
        RECT 65.360 137.180 65.620 137.500 ;
        RECT 64.900 135.820 65.160 136.140 ;
        RECT 64.960 134.010 65.100 135.820 ;
        RECT 65.420 134.780 65.560 137.180 ;
        RECT 65.880 137.160 66.020 140.160 ;
        RECT 67.260 139.540 67.400 148.060 ;
        RECT 68.180 139.880 68.320 151.800 ;
        RECT 68.580 149.080 68.840 149.400 ;
        RECT 68.640 148.380 68.780 149.080 ;
        RECT 68.580 148.060 68.840 148.380 ;
        RECT 68.640 147.360 68.780 148.060 ;
        RECT 68.580 147.040 68.840 147.360 ;
        RECT 69.100 145.060 69.240 165.400 ;
        RECT 70.020 161.300 70.160 166.420 ;
        RECT 69.960 160.980 70.220 161.300 ;
        RECT 69.500 159.960 69.760 160.280 ;
        RECT 69.560 156.200 69.700 159.960 ;
        RECT 69.500 155.880 69.760 156.200 ;
        RECT 69.560 153.820 69.700 155.880 ;
        RECT 69.500 153.500 69.760 153.820 ;
        RECT 70.480 152.460 70.620 180.110 ;
        RECT 70.870 179.485 71.150 179.855 ;
        RECT 70.880 179.340 71.140 179.485 ;
        RECT 71.400 178.300 71.540 182.060 ;
        RECT 72.720 181.720 72.980 182.040 ;
        RECT 73.180 181.720 73.440 182.040 ;
        RECT 72.260 180.020 72.520 180.340 ;
        RECT 71.800 179.340 72.060 179.660 ;
        RECT 71.340 177.980 71.600 178.300 ;
        RECT 70.880 177.640 71.140 177.960 ;
        RECT 70.940 174.900 71.080 177.640 ;
        RECT 71.340 177.300 71.600 177.620 ;
        RECT 70.880 174.580 71.140 174.900 ;
        RECT 71.400 174.560 71.540 177.300 ;
        RECT 71.340 174.240 71.600 174.560 ;
        RECT 71.400 169.120 71.540 174.240 ;
        RECT 71.340 168.800 71.600 169.120 ;
        RECT 71.400 160.700 71.540 168.800 ;
        RECT 70.940 160.560 71.540 160.700 ;
        RECT 70.940 158.240 71.080 160.560 ;
        RECT 70.880 157.920 71.140 158.240 ;
        RECT 70.940 153.480 71.080 157.920 ;
        RECT 70.880 153.160 71.140 153.480 ;
        RECT 71.860 152.800 72.000 179.340 ;
        RECT 72.320 178.300 72.460 180.020 ;
        RECT 72.260 177.980 72.520 178.300 ;
        RECT 72.250 177.445 72.530 177.815 ;
        RECT 72.260 177.300 72.520 177.445 ;
        RECT 72.260 168.460 72.520 168.780 ;
        RECT 72.320 165.720 72.460 168.460 ;
        RECT 72.260 165.400 72.520 165.720 ;
        RECT 72.320 163.680 72.460 165.400 ;
        RECT 72.260 163.360 72.520 163.680 ;
        RECT 72.260 160.300 72.520 160.620 ;
        RECT 72.320 159.260 72.460 160.300 ;
        RECT 72.260 158.940 72.520 159.260 ;
        RECT 72.260 157.240 72.520 157.560 ;
        RECT 72.320 154.840 72.460 157.240 ;
        RECT 72.260 154.520 72.520 154.840 ;
        RECT 71.800 152.480 72.060 152.800 ;
        RECT 70.420 152.140 70.680 152.460 ;
        RECT 70.480 150.420 70.620 152.140 ;
        RECT 70.420 150.100 70.680 150.420 ;
        RECT 70.480 147.700 70.620 150.100 ;
        RECT 70.880 149.080 71.140 149.400 ;
        RECT 70.420 147.380 70.680 147.700 ;
        RECT 69.100 144.920 69.700 145.060 ;
        RECT 69.040 144.320 69.300 144.640 ;
        RECT 68.580 141.600 68.840 141.920 ;
        RECT 68.120 139.560 68.380 139.880 ;
        RECT 66.280 139.220 66.540 139.540 ;
        RECT 67.200 139.220 67.460 139.540 ;
        RECT 65.820 136.840 66.080 137.160 ;
        RECT 65.880 136.480 66.020 136.840 ;
        RECT 65.820 136.160 66.080 136.480 ;
        RECT 65.880 134.780 66.020 136.160 ;
        RECT 65.360 134.460 65.620 134.780 ;
        RECT 65.820 134.460 66.080 134.780 ;
        RECT 65.360 134.010 65.620 134.100 ;
        RECT 64.960 133.870 65.620 134.010 ;
        RECT 65.360 133.780 65.620 133.870 ;
        RECT 65.820 133.780 66.080 134.100 ;
        RECT 65.880 130.700 66.020 133.780 ;
        RECT 64.900 130.380 65.160 130.700 ;
        RECT 65.820 130.380 66.080 130.700 ;
        RECT 64.440 125.620 64.700 125.940 ;
        RECT 63.520 124.690 64.180 124.830 ;
        RECT 63.520 124.600 63.780 124.690 ;
        RECT 64.040 123.900 64.180 124.690 ;
        RECT 63.980 123.580 64.240 123.900 ;
        RECT 62.600 122.220 62.860 122.540 ;
        RECT 64.040 121.180 64.180 123.580 ;
        RECT 64.500 122.880 64.640 125.620 ;
        RECT 64.960 122.880 65.100 130.380 ;
        RECT 66.340 130.360 66.480 139.220 ;
        RECT 68.640 139.200 68.780 141.600 ;
        RECT 68.580 138.880 68.840 139.200 ;
        RECT 68.640 133.760 68.780 138.880 ;
        RECT 69.100 136.480 69.240 144.320 ;
        RECT 69.560 141.580 69.700 144.920 ;
        RECT 69.960 143.640 70.220 143.960 ;
        RECT 70.020 141.920 70.160 143.640 ;
        RECT 69.960 141.600 70.220 141.920 ;
        RECT 69.500 141.260 69.760 141.580 ;
        RECT 70.420 141.260 70.680 141.580 ;
        RECT 69.500 138.880 69.760 139.200 ;
        RECT 69.560 137.500 69.700 138.880 ;
        RECT 69.500 137.180 69.760 137.500 ;
        RECT 69.040 136.160 69.300 136.480 ;
        RECT 68.580 133.440 68.840 133.760 ;
        RECT 66.280 130.040 66.540 130.360 ;
        RECT 66.340 129.340 66.480 130.040 ;
        RECT 66.280 129.020 66.540 129.340 ;
        RECT 68.640 128.320 68.780 133.440 ;
        RECT 69.100 131.380 69.240 136.160 ;
        RECT 69.040 131.060 69.300 131.380 ;
        RECT 69.960 130.040 70.220 130.360 ;
        RECT 69.500 128.680 69.760 129.000 ;
        RECT 68.580 128.000 68.840 128.320 ;
        RECT 64.440 122.560 64.700 122.880 ;
        RECT 64.900 122.560 65.160 122.880 ;
        RECT 63.980 120.860 64.240 121.180 ;
        RECT 62.140 119.500 62.400 119.820 ;
        RECT 62.200 118.460 62.340 119.500 ;
        RECT 64.960 118.460 65.100 122.560 ;
        RECT 68.120 121.880 68.380 122.200 ;
        RECT 62.140 118.140 62.400 118.460 ;
        RECT 64.900 118.140 65.160 118.460 ;
        RECT 66.280 117.800 66.540 118.120 ;
        RECT 63.980 117.460 64.240 117.780 ;
        RECT 64.040 115.060 64.180 117.460 ;
        RECT 66.340 115.740 66.480 117.800 ;
        RECT 66.280 115.420 66.540 115.740 ;
        RECT 63.980 114.740 64.240 115.060 ;
        RECT 68.180 114.720 68.320 121.880 ;
        RECT 68.640 119.480 68.780 128.000 ;
        RECT 69.560 126.620 69.700 128.680 ;
        RECT 69.500 126.300 69.760 126.620 ;
        RECT 70.020 125.600 70.160 130.040 ;
        RECT 69.960 125.280 70.220 125.600 ;
        RECT 70.480 125.260 70.620 141.260 ;
        RECT 70.940 140.220 71.080 149.080 ;
        RECT 71.860 147.360 72.000 152.480 ;
        RECT 71.800 147.040 72.060 147.360 ;
        RECT 72.260 140.920 72.520 141.240 ;
        RECT 70.880 139.900 71.140 140.220 ;
        RECT 70.940 139.200 71.080 139.900 ;
        RECT 72.320 139.880 72.460 140.920 ;
        RECT 72.260 139.560 72.520 139.880 ;
        RECT 70.880 138.880 71.140 139.200 ;
        RECT 70.880 138.200 71.140 138.520 ;
        RECT 70.940 136.820 71.080 138.200 ;
        RECT 70.880 136.500 71.140 136.820 ;
        RECT 72.780 131.040 72.920 181.720 ;
        RECT 73.240 180.340 73.380 181.720 ;
        RECT 73.700 181.020 73.840 182.740 ;
        RECT 73.640 180.700 73.900 181.020 ;
        RECT 73.180 180.020 73.440 180.340 ;
        RECT 73.700 179.660 73.840 180.700 ;
        RECT 75.020 180.360 75.280 180.680 ;
        RECT 74.560 179.680 74.820 180.000 ;
        RECT 73.640 179.340 73.900 179.660 ;
        RECT 73.700 177.960 73.840 179.340 ;
        RECT 74.100 177.980 74.360 178.300 ;
        RECT 73.640 177.640 73.900 177.960 ;
        RECT 73.640 176.960 73.900 177.280 ;
        RECT 74.160 177.135 74.300 177.980 ;
        RECT 73.180 176.620 73.440 176.940 ;
        RECT 73.240 174.560 73.380 176.620 ;
        RECT 73.700 175.580 73.840 176.960 ;
        RECT 74.090 176.765 74.370 177.135 ;
        RECT 74.620 176.940 74.760 179.680 ;
        RECT 75.080 177.815 75.220 180.360 ;
        RECT 75.010 177.445 75.290 177.815 ;
        RECT 75.540 177.620 75.680 183.080 ;
        RECT 76.000 180.680 76.140 189.880 ;
        RECT 76.460 183.820 76.600 190.900 ;
        RECT 84.740 190.200 84.880 193.620 ;
        RECT 85.140 193.280 85.400 193.600 ;
        RECT 78.240 189.880 78.500 190.200 ;
        RECT 84.680 189.880 84.940 190.200 ;
        RECT 76.460 183.740 77.060 183.820 ;
        RECT 76.400 183.680 77.060 183.740 ;
        RECT 76.400 183.420 76.660 183.680 ;
        RECT 76.400 182.740 76.660 183.060 ;
        RECT 75.940 180.360 76.200 180.680 ;
        RECT 75.480 177.300 75.740 177.620 ;
        RECT 75.940 177.300 76.200 177.620 ;
        RECT 74.160 175.580 74.300 176.765 ;
        RECT 74.560 176.620 74.820 176.940 ;
        RECT 75.540 175.580 75.680 177.300 ;
        RECT 73.640 175.260 73.900 175.580 ;
        RECT 74.100 175.260 74.360 175.580 ;
        RECT 75.480 175.260 75.740 175.580 ;
        RECT 73.180 174.240 73.440 174.560 ;
        RECT 75.540 174.220 75.680 175.260 ;
        RECT 76.000 175.240 76.140 177.300 ;
        RECT 76.460 177.280 76.600 182.740 ;
        RECT 76.920 180.340 77.060 183.680 ;
        RECT 77.780 182.740 78.040 183.060 ;
        RECT 77.320 182.060 77.580 182.380 ;
        RECT 76.860 180.020 77.120 180.340 ;
        RECT 76.920 179.320 77.060 180.020 ;
        RECT 77.380 179.660 77.520 182.060 ;
        RECT 77.320 179.340 77.580 179.660 ;
        RECT 76.860 179.000 77.120 179.320 ;
        RECT 77.840 177.620 77.980 182.740 ;
        RECT 77.780 177.300 78.040 177.620 ;
        RECT 76.400 176.960 76.660 177.280 ;
        RECT 77.320 177.020 77.580 177.280 ;
        RECT 77.320 176.960 77.980 177.020 ;
        RECT 77.380 176.880 77.980 176.960 ;
        RECT 77.840 176.600 77.980 176.880 ;
        RECT 77.320 176.280 77.580 176.600 ;
        RECT 77.780 176.280 78.040 176.600 ;
        RECT 75.940 174.920 76.200 175.240 ;
        RECT 76.000 174.220 76.140 174.920 ;
        RECT 75.480 173.900 75.740 174.220 ;
        RECT 75.940 173.900 76.200 174.220 ;
        RECT 73.180 169.140 73.440 169.460 ;
        RECT 73.240 166.740 73.380 169.140 ;
        RECT 76.400 168.120 76.660 168.440 ;
        RECT 73.640 166.760 73.900 167.080 ;
        RECT 73.180 166.420 73.440 166.740 ;
        RECT 73.180 165.400 73.440 165.720 ;
        RECT 73.240 163.680 73.380 165.400 ;
        RECT 73.180 163.360 73.440 163.680 ;
        RECT 73.240 158.240 73.380 163.360 ;
        RECT 73.180 157.920 73.440 158.240 ;
        RECT 73.180 146.360 73.440 146.680 ;
        RECT 73.240 145.660 73.380 146.360 ;
        RECT 73.180 145.340 73.440 145.660 ;
        RECT 72.720 130.720 72.980 131.040 ;
        RECT 73.180 130.040 73.440 130.360 ;
        RECT 71.800 128.570 72.060 128.660 ;
        RECT 70.940 128.430 72.060 128.570 ;
        RECT 70.940 126.620 71.080 128.430 ;
        RECT 71.800 128.340 72.060 128.430 ;
        RECT 70.880 126.300 71.140 126.620 ;
        RECT 73.240 125.260 73.380 130.040 ;
        RECT 70.420 124.940 70.680 125.260 ;
        RECT 73.180 124.940 73.440 125.260 ;
        RECT 69.960 124.600 70.220 124.920 ;
        RECT 70.020 120.160 70.160 124.600 ;
        RECT 69.960 119.840 70.220 120.160 ;
        RECT 68.580 119.160 68.840 119.480 ;
        RECT 68.640 117.440 68.780 119.160 ;
        RECT 68.580 117.120 68.840 117.440 ;
        RECT 70.480 115.060 70.620 124.940 ;
        RECT 73.240 122.540 73.380 124.940 ;
        RECT 73.700 123.220 73.840 166.760 ;
        RECT 74.560 165.740 74.820 166.060 ;
        RECT 74.100 159.960 74.360 160.280 ;
        RECT 74.160 158.920 74.300 159.960 ;
        RECT 74.100 158.600 74.360 158.920 ;
        RECT 74.160 158.240 74.300 158.600 ;
        RECT 74.100 157.920 74.360 158.240 ;
        RECT 74.620 153.220 74.760 165.740 ;
        RECT 75.020 157.580 75.280 157.900 ;
        RECT 75.080 156.200 75.220 157.580 ;
        RECT 75.940 157.240 76.200 157.560 ;
        RECT 75.020 155.880 75.280 156.200 ;
        RECT 74.160 153.080 74.760 153.220 ;
        RECT 74.160 152.800 74.300 153.080 ;
        RECT 74.100 152.480 74.360 152.800 ;
        RECT 74.160 136.140 74.300 152.480 ;
        RECT 75.020 151.800 75.280 152.120 ;
        RECT 75.080 150.760 75.220 151.800 ;
        RECT 76.000 150.760 76.140 157.240 ;
        RECT 76.460 155.860 76.600 168.120 ;
        RECT 76.860 157.240 77.120 157.560 ;
        RECT 76.400 155.540 76.660 155.860 ;
        RECT 75.020 150.440 75.280 150.760 ;
        RECT 75.940 150.440 76.200 150.760 ;
        RECT 76.400 149.080 76.660 149.400 ;
        RECT 75.940 143.980 76.200 144.300 ;
        RECT 74.100 135.820 74.360 136.140 ;
        RECT 74.160 131.380 74.300 135.820 ;
        RECT 74.100 131.060 74.360 131.380 ;
        RECT 73.640 122.900 73.900 123.220 ;
        RECT 73.180 122.220 73.440 122.540 ;
        RECT 73.700 120.160 73.840 122.900 ;
        RECT 73.640 119.840 73.900 120.160 ;
        RECT 70.880 117.460 71.140 117.780 ;
        RECT 70.940 115.740 71.080 117.460 ;
        RECT 73.640 117.120 73.900 117.440 ;
        RECT 70.880 115.420 71.140 115.740 ;
        RECT 70.420 114.740 70.680 115.060 ;
        RECT 68.120 114.400 68.380 114.720 ;
        RECT 70.480 112.680 70.620 114.740 ;
        RECT 70.420 112.360 70.680 112.680 ;
        RECT 73.180 109.640 73.440 109.960 ;
        RECT 61.680 108.620 61.940 108.940 ;
        RECT 61.740 107.580 61.880 108.620 ;
        RECT 70.880 108.280 71.140 108.600 ;
        RECT 61.680 107.260 61.940 107.580 ;
        RECT 61.220 106.580 61.480 106.900 ;
        RECT 50.640 105.900 50.900 106.220 ;
        RECT 60.820 106.160 61.420 106.300 ;
        RECT 50.180 104.540 50.440 104.860 ;
        RECT 50.700 103.840 50.840 105.900 ;
        RECT 56.620 105.560 56.880 105.880 ;
        RECT 50.640 103.520 50.900 103.840 ;
        RECT 56.680 103.500 56.820 105.560 ;
        RECT 61.280 104.180 61.420 106.160 ;
        RECT 64.440 105.900 64.700 106.220 ;
        RECT 63.980 105.560 64.240 105.880 ;
        RECT 61.220 103.860 61.480 104.180 ;
        RECT 56.620 103.180 56.880 103.500 ;
        RECT 54.320 102.840 54.580 103.160 ;
        RECT 61.680 102.840 61.940 103.160 ;
        RECT 54.380 101.800 54.520 102.840 ;
        RECT 61.740 101.800 61.880 102.840 ;
        RECT 64.040 101.800 64.180 105.560 ;
        RECT 64.500 103.500 64.640 105.900 ;
        RECT 70.940 103.500 71.080 108.280 ;
        RECT 64.440 103.180 64.700 103.500 ;
        RECT 70.880 103.180 71.140 103.500 ;
        RECT 73.240 102.220 73.380 109.640 ;
        RECT 73.700 106.900 73.840 117.120 ;
        RECT 74.160 110.300 74.300 131.060 ;
        RECT 75.020 130.040 75.280 130.360 ;
        RECT 75.080 129.340 75.220 130.040 ;
        RECT 75.020 129.020 75.280 129.340 ;
        RECT 75.080 128.660 75.220 129.020 ;
        RECT 75.020 128.340 75.280 128.660 ;
        RECT 75.480 119.160 75.740 119.480 ;
        RECT 75.540 118.120 75.680 119.160 ;
        RECT 75.480 117.800 75.740 118.120 ;
        RECT 74.100 109.980 74.360 110.300 ;
        RECT 75.480 108.960 75.740 109.280 ;
        RECT 74.100 108.620 74.360 108.940 ;
        RECT 73.640 106.580 73.900 106.900 ;
        RECT 73.700 104.180 73.840 106.580 ;
        RECT 74.160 104.860 74.300 108.620 ;
        RECT 74.100 104.540 74.360 104.860 ;
        RECT 73.640 103.860 73.900 104.180 ;
        RECT 73.240 102.080 74.300 102.220 ;
        RECT 54.320 101.480 54.580 101.800 ;
        RECT 61.680 101.480 61.940 101.800 ;
        RECT 63.980 101.480 64.240 101.800 ;
        RECT 54.780 100.120 55.040 100.440 ;
        RECT 60.760 100.120 61.020 100.440 ;
        RECT 68.120 100.120 68.380 100.440 ;
        RECT 50.170 90.660 50.450 91.170 ;
        RECT 48.860 90.520 50.450 90.660 ;
        RECT 54.840 90.660 54.980 100.120 ;
        RECT 56.150 90.660 56.430 91.170 ;
        RECT 54.840 90.520 56.430 90.660 ;
        RECT 60.820 90.660 60.960 100.120 ;
        RECT 68.180 91.170 68.320 100.120 ;
        RECT 74.160 91.170 74.300 102.080 ;
        RECT 75.540 101.460 75.680 108.960 ;
        RECT 76.000 106.810 76.140 143.980 ;
        RECT 76.460 129.340 76.600 149.080 ;
        RECT 76.920 136.480 77.060 157.240 ;
        RECT 77.380 150.080 77.520 176.280 ;
        RECT 77.840 174.560 77.980 176.280 ;
        RECT 78.300 174.560 78.440 189.880 ;
        RECT 85.200 185.860 85.340 193.280 ;
        RECT 85.600 188.070 85.860 188.160 ;
        RECT 86.580 188.070 86.720 193.620 ;
        RECT 87.500 191.220 87.640 201.190 ;
        RECT 107.680 196.000 107.940 196.320 ;
        RECT 121.020 196.000 121.280 196.320 ;
        RECT 107.740 194.280 107.880 196.000 ;
        RECT 116.420 195.660 116.680 195.980 ;
        RECT 109.060 195.320 109.320 195.640 ;
        RECT 107.680 193.960 107.940 194.280 ;
        RECT 90.200 193.620 90.460 193.940 ;
        RECT 87.440 190.900 87.700 191.220 ;
        RECT 87.500 188.160 87.640 190.900 ;
        RECT 90.260 188.500 90.400 193.620 ;
        RECT 109.120 193.600 109.260 195.320 ;
        RECT 115.960 193.620 116.220 193.940 ;
        RECT 104.920 193.280 105.180 193.600 ;
        RECT 107.220 193.280 107.480 193.600 ;
        RECT 109.060 193.280 109.320 193.600 ;
        RECT 110.900 193.280 111.160 193.600 ;
        RECT 111.820 193.280 112.080 193.600 ;
        RECT 90.660 192.600 90.920 192.920 ;
        RECT 93.880 192.600 94.140 192.920 ;
        RECT 97.560 192.600 97.820 192.920 ;
        RECT 90.720 190.540 90.860 192.600 ;
        RECT 93.940 191.220 94.080 192.600 ;
        RECT 93.880 190.900 94.140 191.220 ;
        RECT 90.660 190.220 90.920 190.540 ;
        RECT 90.200 188.180 90.460 188.500 ;
        RECT 91.120 188.180 91.380 188.500 ;
        RECT 85.600 187.930 86.720 188.070 ;
        RECT 85.600 187.840 85.860 187.930 ;
        RECT 85.200 185.780 85.800 185.860 ;
        RECT 86.580 185.780 86.720 187.930 ;
        RECT 87.440 187.840 87.700 188.160 ;
        RECT 85.200 185.720 85.860 185.780 ;
        RECT 85.600 185.460 85.860 185.720 ;
        RECT 86.520 185.460 86.780 185.780 ;
        RECT 79.620 185.120 79.880 185.440 ;
        RECT 79.680 182.720 79.820 185.120 ;
        RECT 81.000 184.440 81.260 184.760 ;
        RECT 84.680 184.440 84.940 184.760 ;
        RECT 79.620 182.400 79.880 182.720 ;
        RECT 79.160 181.720 79.420 182.040 ;
        RECT 78.700 175.260 78.960 175.580 ;
        RECT 78.760 174.560 78.900 175.260 ;
        RECT 77.780 174.240 78.040 174.560 ;
        RECT 78.240 174.240 78.500 174.560 ;
        RECT 78.700 174.240 78.960 174.560 ;
        RECT 78.240 173.560 78.500 173.880 ;
        RECT 78.300 170.140 78.440 173.560 ;
        RECT 78.240 169.820 78.500 170.140 ;
        RECT 78.700 169.140 78.960 169.460 ;
        RECT 78.240 168.120 78.500 168.440 ;
        RECT 78.300 163.680 78.440 168.120 ;
        RECT 78.760 164.020 78.900 169.140 ;
        RECT 78.700 163.700 78.960 164.020 ;
        RECT 78.240 163.360 78.500 163.680 ;
        RECT 78.760 161.640 78.900 163.700 ;
        RECT 78.700 161.320 78.960 161.640 ;
        RECT 78.240 157.920 78.500 158.240 ;
        RECT 78.700 157.920 78.960 158.240 ;
        RECT 78.300 155.860 78.440 157.920 ;
        RECT 78.760 156.200 78.900 157.920 ;
        RECT 78.700 155.880 78.960 156.200 ;
        RECT 78.240 155.540 78.500 155.860 ;
        RECT 78.700 154.860 78.960 155.180 ;
        RECT 77.780 150.100 78.040 150.420 ;
        RECT 77.320 149.760 77.580 150.080 ;
        RECT 77.840 148.380 77.980 150.100 ;
        RECT 77.780 148.060 78.040 148.380 ;
        RECT 78.240 147.040 78.500 147.360 ;
        RECT 78.300 146.680 78.440 147.040 ;
        RECT 78.240 146.360 78.500 146.680 ;
        RECT 78.760 144.980 78.900 154.860 ;
        RECT 78.700 144.660 78.960 144.980 ;
        RECT 78.700 137.180 78.960 137.500 ;
        RECT 76.860 136.160 77.120 136.480 ;
        RECT 77.780 135.480 78.040 135.800 ;
        RECT 76.400 129.020 76.660 129.340 ;
        RECT 76.860 128.680 77.120 129.000 ;
        RECT 76.920 128.320 77.060 128.680 ;
        RECT 76.860 128.000 77.120 128.320 ;
        RECT 76.920 126.620 77.060 128.000 ;
        RECT 76.860 126.300 77.120 126.620 ;
        RECT 77.840 109.960 77.980 135.480 ;
        RECT 78.760 132.060 78.900 137.180 ;
        RECT 79.220 136.820 79.360 181.720 ;
        RECT 81.060 180.340 81.200 184.440 ;
        RECT 84.740 183.400 84.880 184.440 ;
        RECT 84.680 183.080 84.940 183.400 ;
        RECT 83.300 181.720 83.560 182.040 ;
        RECT 83.360 181.020 83.500 181.720 ;
        RECT 83.300 180.700 83.560 181.020 ;
        RECT 85.660 180.680 85.800 185.460 ;
        RECT 85.600 180.360 85.860 180.680 ;
        RECT 81.000 180.020 81.260 180.340 ;
        RECT 83.760 179.340 84.020 179.660 ;
        RECT 81.460 179.000 81.720 179.320 ;
        RECT 83.820 179.175 83.960 179.340 ;
        RECT 81.520 175.580 81.660 179.000 ;
        RECT 83.750 178.805 84.030 179.175 ;
        RECT 83.820 177.815 83.960 178.805 ;
        RECT 83.750 177.445 84.030 177.815 ;
        RECT 84.220 176.280 84.480 176.600 ;
        RECT 81.460 175.260 81.720 175.580 ;
        RECT 82.840 174.920 83.100 175.240 ;
        RECT 82.900 174.560 83.040 174.920 ;
        RECT 84.280 174.560 84.420 176.280 ;
        RECT 85.660 175.580 85.800 180.360 ;
        RECT 86.580 177.960 86.720 185.460 ;
        RECT 87.500 183.400 87.640 187.840 ;
        RECT 90.260 185.440 90.400 188.180 ;
        RECT 91.180 186.120 91.320 188.180 ;
        RECT 97.620 188.160 97.760 192.600 ;
        RECT 104.980 191.900 105.120 193.280 ;
        RECT 105.840 192.600 106.100 192.920 ;
        RECT 104.920 191.580 105.180 191.900 ;
        RECT 105.900 191.220 106.040 192.600 ;
        RECT 98.480 190.900 98.740 191.220 ;
        RECT 105.840 190.900 106.100 191.220 ;
        RECT 98.020 190.560 98.280 190.880 ;
        RECT 98.080 189.180 98.220 190.560 ;
        RECT 98.020 188.860 98.280 189.180 ;
        RECT 97.560 187.840 97.820 188.160 ;
        RECT 96.640 187.160 96.900 187.480 ;
        RECT 91.120 185.800 91.380 186.120 ;
        RECT 96.700 185.780 96.840 187.160 ;
        RECT 98.540 186.460 98.680 190.900 ;
        RECT 102.620 188.520 102.880 188.840 ;
        RECT 102.160 187.160 102.420 187.480 ;
        RECT 102.220 186.460 102.360 187.160 ;
        RECT 102.680 186.460 102.820 188.520 ;
        RECT 98.480 186.140 98.740 186.460 ;
        RECT 102.160 186.140 102.420 186.460 ;
        RECT 102.620 186.140 102.880 186.460 ;
        RECT 105.900 186.120 106.040 190.900 ;
        RECT 107.280 188.160 107.420 193.280 ;
        RECT 107.680 192.600 107.940 192.920 ;
        RECT 107.740 191.220 107.880 192.600 ;
        RECT 107.680 190.900 107.940 191.220 ;
        RECT 109.980 189.880 110.240 190.200 ;
        RECT 110.440 189.880 110.700 190.200 ;
        RECT 110.040 188.500 110.180 189.880 ;
        RECT 109.980 188.180 110.240 188.500 ;
        RECT 107.220 187.840 107.480 188.160 ;
        RECT 107.680 187.500 107.940 187.820 ;
        RECT 105.840 185.800 106.100 186.120 ;
        RECT 96.640 185.460 96.900 185.780 ;
        RECT 90.200 185.120 90.460 185.440 ;
        RECT 91.580 184.780 91.840 185.100 ;
        RECT 91.640 183.740 91.780 184.780 ;
        RECT 96.700 183.740 96.840 185.460 ;
        RECT 99.400 185.120 99.660 185.440 ;
        RECT 97.100 184.440 97.360 184.760 ;
        RECT 98.940 184.500 99.200 184.760 ;
        RECT 98.540 184.440 99.200 184.500 ;
        RECT 90.660 183.420 90.920 183.740 ;
        RECT 91.580 183.420 91.840 183.740 ;
        RECT 96.640 183.420 96.900 183.740 ;
        RECT 87.440 183.080 87.700 183.400 ;
        RECT 87.500 181.020 87.640 183.080 ;
        RECT 87.440 180.700 87.700 181.020 ;
        RECT 86.520 177.640 86.780 177.960 ;
        RECT 87.500 177.620 87.640 180.700 ;
        RECT 87.440 177.300 87.700 177.620 ;
        RECT 85.600 175.260 85.860 175.580 ;
        RECT 82.840 174.240 83.100 174.560 ;
        RECT 84.220 174.240 84.480 174.560 ;
        RECT 80.080 173.900 80.340 174.220 ;
        RECT 81.920 174.130 82.180 174.220 ;
        RECT 81.920 173.990 82.580 174.130 ;
        RECT 81.920 173.900 82.180 173.990 ;
        RECT 79.620 146.360 79.880 146.680 ;
        RECT 79.680 145.320 79.820 146.360 ;
        RECT 79.620 145.000 79.880 145.320 ;
        RECT 80.140 144.640 80.280 173.900 ;
        RECT 80.540 162.680 80.800 163.000 ;
        RECT 80.600 161.980 80.740 162.680 ;
        RECT 80.540 161.660 80.800 161.980 ;
        RECT 80.600 158.580 80.740 161.660 ;
        RECT 81.000 159.960 81.260 160.280 ;
        RECT 80.540 158.260 80.800 158.580 ;
        RECT 81.060 157.900 81.200 159.960 ;
        RECT 81.000 157.580 81.260 157.900 ;
        RECT 81.460 147.040 81.720 147.360 ;
        RECT 81.920 147.040 82.180 147.360 ;
        RECT 80.080 144.320 80.340 144.640 ;
        RECT 80.080 143.640 80.340 143.960 ;
        RECT 79.620 138.200 79.880 138.520 ;
        RECT 79.160 136.500 79.420 136.820 ;
        RECT 79.680 136.480 79.820 138.200 ;
        RECT 79.620 136.160 79.880 136.480 ;
        RECT 79.160 135.480 79.420 135.800 ;
        RECT 79.220 134.440 79.360 135.480 ;
        RECT 79.160 134.120 79.420 134.440 ;
        RECT 78.700 131.740 78.960 132.060 ;
        RECT 79.160 131.290 79.420 131.380 ;
        RECT 79.160 131.150 79.820 131.290 ;
        RECT 79.160 131.060 79.420 131.150 ;
        RECT 78.700 130.380 78.960 130.700 ;
        RECT 78.240 128.340 78.500 128.660 ;
        RECT 78.300 127.640 78.440 128.340 ;
        RECT 78.240 127.320 78.500 127.640 ;
        RECT 78.300 119.480 78.440 127.320 ;
        RECT 78.760 120.160 78.900 130.380 ;
        RECT 79.680 128.320 79.820 131.150 ;
        RECT 80.140 129.340 80.280 143.640 ;
        RECT 81.520 139.540 81.660 147.040 ;
        RECT 81.980 139.540 82.120 147.040 ;
        RECT 81.460 139.220 81.720 139.540 ;
        RECT 81.920 139.220 82.180 139.540 ;
        RECT 81.520 136.480 81.660 139.220 ;
        RECT 81.980 136.480 82.120 139.220 ;
        RECT 81.460 136.160 81.720 136.480 ;
        RECT 81.920 136.160 82.180 136.480 ;
        RECT 82.440 133.760 82.580 173.990 ;
        RECT 87.500 171.840 87.640 177.300 ;
        RECT 90.720 174.900 90.860 183.420 ;
        RECT 96.180 183.080 96.440 183.400 ;
        RECT 91.120 182.740 91.380 183.060 ;
        RECT 91.180 182.040 91.320 182.740 ;
        RECT 91.120 181.720 91.380 182.040 ;
        RECT 94.800 181.720 95.060 182.040 ;
        RECT 94.860 180.340 95.000 181.720 ;
        RECT 94.800 180.020 95.060 180.340 ;
        RECT 95.720 179.680 95.980 180.000 ;
        RECT 95.780 178.300 95.920 179.680 ;
        RECT 96.240 178.300 96.380 183.080 ;
        RECT 95.720 177.980 95.980 178.300 ;
        RECT 96.180 177.980 96.440 178.300 ;
        RECT 97.160 177.620 97.300 184.440 ;
        RECT 98.540 184.360 99.140 184.440 ;
        RECT 98.540 180.340 98.680 184.360 ;
        RECT 99.460 181.020 99.600 185.120 ;
        RECT 101.240 183.420 101.500 183.740 ;
        RECT 99.860 183.080 100.120 183.400 ;
        RECT 99.920 181.020 100.060 183.080 ;
        RECT 99.400 180.700 99.660 181.020 ;
        RECT 99.860 180.700 100.120 181.020 ;
        RECT 98.480 180.020 98.740 180.340 ;
        RECT 100.780 179.680 101.040 180.000 ;
        RECT 100.840 177.620 100.980 179.680 ;
        RECT 101.300 177.635 101.440 183.420 ;
        RECT 105.900 182.720 106.040 185.800 ;
        RECT 105.840 182.400 106.100 182.720 ;
        RECT 105.900 180.680 106.040 182.400 ;
        RECT 105.840 180.360 106.100 180.680 ;
        RECT 105.840 179.680 106.100 180.000 ;
        RECT 107.220 179.680 107.480 180.000 ;
        RECT 103.080 179.000 103.340 179.320 ;
        RECT 101.700 177.980 101.960 178.300 ;
        RECT 97.100 177.300 97.360 177.620 ;
        RECT 100.780 177.300 101.040 177.620 ;
        RECT 101.240 177.315 101.500 177.635 ;
        RECT 101.760 177.620 101.900 177.980 ;
        RECT 101.700 177.300 101.960 177.620 ;
        RECT 102.150 177.445 102.430 177.815 ;
        RECT 90.660 174.580 90.920 174.900 ;
        RECT 97.160 172.860 97.300 177.300 ;
        RECT 99.860 176.280 100.120 176.600 ;
        RECT 97.100 172.540 97.360 172.860 ;
        RECT 98.480 172.200 98.740 172.520 ;
        RECT 87.440 171.520 87.700 171.840 ;
        RECT 90.200 171.520 90.460 171.840 ;
        RECT 90.260 169.460 90.400 171.520 ;
        RECT 90.660 170.840 90.920 171.160 ;
        RECT 90.720 169.800 90.860 170.840 ;
        RECT 98.540 170.140 98.680 172.200 ;
        RECT 92.040 169.820 92.300 170.140 ;
        RECT 93.880 169.820 94.140 170.140 ;
        RECT 98.480 169.820 98.740 170.140 ;
        RECT 90.660 169.480 90.920 169.800 ;
        RECT 92.100 169.460 92.240 169.820 ;
        RECT 90.200 169.140 90.460 169.460 ;
        RECT 92.040 169.140 92.300 169.460 ;
        RECT 87.440 168.800 87.700 169.120 ;
        RECT 84.220 168.460 84.480 168.780 ;
        RECT 83.300 168.120 83.560 168.440 ;
        RECT 82.840 166.080 83.100 166.400 ;
        RECT 82.900 164.700 83.040 166.080 ;
        RECT 82.840 164.380 83.100 164.700 ;
        RECT 83.360 163.680 83.500 168.120 ;
        RECT 84.280 167.080 84.420 168.460 ;
        RECT 84.220 166.760 84.480 167.080 ;
        RECT 87.500 164.700 87.640 168.800 ;
        RECT 90.260 166.400 90.400 169.140 ;
        RECT 90.200 166.080 90.460 166.400 ;
        RECT 87.440 164.380 87.700 164.700 ;
        RECT 83.300 163.360 83.560 163.680 ;
        RECT 90.260 160.960 90.400 166.080 ;
        RECT 93.940 164.020 94.080 169.820 ;
        RECT 95.720 166.420 95.980 166.740 ;
        RECT 93.880 163.700 94.140 164.020 ;
        RECT 90.660 162.680 90.920 163.000 ;
        RECT 90.720 161.980 90.860 162.680 ;
        RECT 90.660 161.660 90.920 161.980 ;
        RECT 93.880 161.320 94.140 161.640 ;
        RECT 83.300 160.640 83.560 160.960 ;
        RECT 90.200 160.640 90.460 160.960 ;
        RECT 83.360 155.860 83.500 160.640 ;
        RECT 87.900 159.960 88.160 160.280 ;
        RECT 87.960 158.580 88.100 159.960 ;
        RECT 87.900 158.260 88.160 158.580 ;
        RECT 90.260 158.240 90.400 160.640 ;
        RECT 93.940 159.260 94.080 161.320 ;
        RECT 95.780 160.280 95.920 166.420 ;
        RECT 97.100 162.680 97.360 163.000 ;
        RECT 96.640 160.980 96.900 161.300 ;
        RECT 95.720 159.960 95.980 160.280 ;
        RECT 93.880 158.940 94.140 159.260 ;
        RECT 95.780 158.240 95.920 159.960 ;
        RECT 96.700 159.260 96.840 160.980 ;
        RECT 96.640 158.940 96.900 159.260 ;
        RECT 97.160 158.240 97.300 162.680 ;
        RECT 98.940 158.600 99.200 158.920 ;
        RECT 83.760 157.920 84.020 158.240 ;
        RECT 90.200 157.920 90.460 158.240 ;
        RECT 93.880 157.920 94.140 158.240 ;
        RECT 95.720 157.920 95.980 158.240 ;
        RECT 97.100 157.920 97.360 158.240 ;
        RECT 83.820 155.860 83.960 157.920 ;
        RECT 83.300 155.540 83.560 155.860 ;
        RECT 83.760 155.540 84.020 155.860 ;
        RECT 82.840 154.860 83.100 155.180 ;
        RECT 82.900 134.100 83.040 154.860 ;
        RECT 86.520 152.480 86.780 152.800 ;
        RECT 85.600 150.780 85.860 151.100 ;
        RECT 85.140 149.760 85.400 150.080 ;
        RECT 85.200 148.380 85.340 149.760 ;
        RECT 85.140 148.060 85.400 148.380 ;
        RECT 83.300 147.720 83.560 148.040 ;
        RECT 83.360 147.360 83.500 147.720 ;
        RECT 83.300 147.040 83.560 147.360 ;
        RECT 83.360 139.540 83.500 147.040 ;
        RECT 85.200 144.640 85.340 148.060 ;
        RECT 85.660 147.700 85.800 150.780 ;
        RECT 86.060 150.100 86.320 150.420 ;
        RECT 85.600 147.380 85.860 147.700 ;
        RECT 86.120 146.680 86.260 150.100 ;
        RECT 86.580 147.360 86.720 152.480 ;
        RECT 90.260 150.080 90.400 157.920 ;
        RECT 93.940 153.480 94.080 157.920 ;
        RECT 99.000 155.860 99.140 158.600 ;
        RECT 98.940 155.540 99.200 155.860 ;
        RECT 99.400 155.540 99.660 155.860 ;
        RECT 97.560 154.520 97.820 154.840 ;
        RECT 93.880 153.160 94.140 153.480 ;
        RECT 95.720 153.160 95.980 153.480 ;
        RECT 92.960 151.800 93.220 152.120 ;
        RECT 93.020 150.760 93.160 151.800 ;
        RECT 92.960 150.440 93.220 150.760 ;
        RECT 90.200 149.760 90.460 150.080 ;
        RECT 91.120 149.760 91.380 150.080 ;
        RECT 86.980 149.080 87.240 149.400 ;
        RECT 90.660 149.080 90.920 149.400 ;
        RECT 86.520 147.040 86.780 147.360 ;
        RECT 86.060 146.360 86.320 146.680 ;
        RECT 86.120 145.660 86.260 146.360 ;
        RECT 86.060 145.340 86.320 145.660 ;
        RECT 86.060 144.660 86.320 144.980 ;
        RECT 85.140 144.320 85.400 144.640 ;
        RECT 83.300 139.220 83.560 139.540 ;
        RECT 83.360 136.480 83.500 139.220 ;
        RECT 85.200 139.200 85.340 144.320 ;
        RECT 86.120 140.220 86.260 144.660 ;
        RECT 86.060 139.900 86.320 140.220 ;
        RECT 85.140 138.880 85.400 139.200 ;
        RECT 85.200 136.820 85.340 138.880 ;
        RECT 86.120 137.500 86.260 139.900 ;
        RECT 86.060 137.180 86.320 137.500 ;
        RECT 85.140 136.500 85.400 136.820 ;
        RECT 83.300 136.160 83.560 136.480 ;
        RECT 82.840 133.780 83.100 134.100 ;
        RECT 82.380 133.440 82.640 133.760 ;
        RECT 83.300 133.100 83.560 133.420 ;
        RECT 81.460 132.760 81.720 133.080 ;
        RECT 81.000 130.040 81.260 130.360 ;
        RECT 81.060 129.340 81.200 130.040 ;
        RECT 80.080 129.020 80.340 129.340 ;
        RECT 81.000 129.020 81.260 129.340 ;
        RECT 79.620 128.000 79.880 128.320 ;
        RECT 79.680 126.280 79.820 128.000 ;
        RECT 79.620 125.960 79.880 126.280 ;
        RECT 79.680 120.500 79.820 125.960 ;
        RECT 79.620 120.180 79.880 120.500 ;
        RECT 78.700 119.840 78.960 120.160 ;
        RECT 78.240 119.160 78.500 119.480 ;
        RECT 78.300 118.460 78.440 119.160 ;
        RECT 78.240 118.140 78.500 118.460 ;
        RECT 78.760 117.440 78.900 119.840 ;
        RECT 81.000 119.160 81.260 119.480 ;
        RECT 81.060 117.780 81.200 119.160 ;
        RECT 81.000 117.460 81.260 117.780 ;
        RECT 78.700 117.120 78.960 117.440 ;
        RECT 78.760 115.740 78.900 117.120 ;
        RECT 78.700 115.420 78.960 115.740 ;
        RECT 79.220 112.340 80.280 112.420 ;
        RECT 79.160 112.280 80.280 112.340 ;
        RECT 79.160 112.020 79.420 112.280 ;
        RECT 80.140 112.000 80.280 112.280 ;
        RECT 79.620 111.680 79.880 112.000 ;
        RECT 80.080 111.680 80.340 112.000 ;
        RECT 77.780 109.640 78.040 109.960 ;
        RECT 79.680 106.900 79.820 111.680 ;
        RECT 76.400 106.810 76.660 106.900 ;
        RECT 76.000 106.670 76.660 106.810 ;
        RECT 76.400 106.580 76.660 106.670 ;
        RECT 79.620 106.580 79.880 106.900 ;
        RECT 78.240 105.900 78.500 106.220 ;
        RECT 77.320 105.560 77.580 105.880 ;
        RECT 77.780 105.560 78.040 105.880 ;
        RECT 77.380 104.180 77.520 105.560 ;
        RECT 77.320 103.860 77.580 104.180 ;
        RECT 77.840 101.800 77.980 105.560 ;
        RECT 78.300 103.840 78.440 105.900 ;
        RECT 81.520 105.790 81.660 132.760 ;
        RECT 83.360 129.340 83.500 133.100 ;
        RECT 83.300 129.020 83.560 129.340 ;
        RECT 85.140 128.000 85.400 128.320 ;
        RECT 83.300 127.320 83.560 127.640 ;
        RECT 81.920 124.940 82.180 125.260 ;
        RECT 81.980 123.900 82.120 124.940 ;
        RECT 81.920 123.580 82.180 123.900 ;
        RECT 83.360 123.220 83.500 127.320 ;
        RECT 83.760 125.280 84.020 125.600 ;
        RECT 83.820 123.900 83.960 125.280 ;
        RECT 83.760 123.580 84.020 123.900 ;
        RECT 82.380 122.900 82.640 123.220 ;
        RECT 83.300 122.900 83.560 123.220 ;
        RECT 82.440 120.160 82.580 122.900 ;
        RECT 83.760 120.180 84.020 120.500 ;
        RECT 82.380 119.840 82.640 120.160 ;
        RECT 82.840 119.160 83.100 119.480 ;
        RECT 82.900 114.380 83.040 119.160 ;
        RECT 83.820 117.440 83.960 120.180 ;
        RECT 84.220 119.840 84.480 120.160 ;
        RECT 84.280 118.460 84.420 119.840 ;
        RECT 84.680 119.160 84.940 119.480 ;
        RECT 84.220 118.140 84.480 118.460 ;
        RECT 83.760 117.120 84.020 117.440 ;
        RECT 83.820 115.740 83.960 117.120 ;
        RECT 83.760 115.420 84.020 115.740 ;
        RECT 84.740 115.060 84.880 119.160 ;
        RECT 85.200 118.460 85.340 128.000 ;
        RECT 85.140 118.140 85.400 118.460 ;
        RECT 85.140 117.460 85.400 117.780 ;
        RECT 85.200 115.060 85.340 117.460 ;
        RECT 84.680 114.740 84.940 115.060 ;
        RECT 85.140 114.740 85.400 115.060 ;
        RECT 82.840 114.060 83.100 114.380 ;
        RECT 81.920 111.680 82.180 112.000 ;
        RECT 81.980 109.280 82.120 111.680 ;
        RECT 81.920 108.960 82.180 109.280 ;
        RECT 81.980 106.560 82.120 108.960 ;
        RECT 85.200 106.560 85.340 114.740 ;
        RECT 85.600 108.620 85.860 108.940 ;
        RECT 81.920 106.240 82.180 106.560 ;
        RECT 85.140 106.240 85.400 106.560 ;
        RECT 81.520 105.650 82.120 105.790 ;
        RECT 78.240 103.520 78.500 103.840 ;
        RECT 81.980 103.160 82.120 105.650 ;
        RECT 85.200 104.180 85.340 106.240 ;
        RECT 85.660 104.860 85.800 108.620 ;
        RECT 86.060 108.280 86.320 108.600 ;
        RECT 85.600 104.540 85.860 104.860 ;
        RECT 85.140 103.860 85.400 104.180 ;
        RECT 81.920 102.840 82.180 103.160 ;
        RECT 77.780 101.480 78.040 101.800 ;
        RECT 75.480 101.140 75.740 101.460 ;
        RECT 80.080 100.120 80.340 100.440 ;
        RECT 80.140 91.170 80.280 100.120 ;
        RECT 86.120 91.170 86.260 108.280 ;
        RECT 87.040 106.900 87.180 149.080 ;
        RECT 90.200 147.380 90.460 147.700 ;
        RECT 90.260 145.660 90.400 147.380 ;
        RECT 90.200 145.340 90.460 145.660 ;
        RECT 90.720 144.980 90.860 149.080 ;
        RECT 91.180 145.570 91.320 149.760 ;
        RECT 95.780 147.360 95.920 153.160 ;
        RECT 93.880 147.040 94.140 147.360 ;
        RECT 95.720 147.040 95.980 147.360 ;
        RECT 96.180 147.040 96.440 147.360 ;
        RECT 91.580 145.570 91.840 145.660 ;
        RECT 91.180 145.430 91.840 145.570 ;
        RECT 91.580 145.340 91.840 145.430 ;
        RECT 90.660 144.660 90.920 144.980 ;
        RECT 90.660 138.880 90.920 139.200 ;
        RECT 87.440 135.820 87.700 136.140 ;
        RECT 87.500 134.780 87.640 135.820 ;
        RECT 90.720 135.800 90.860 138.880 ;
        RECT 91.120 138.200 91.380 138.520 ;
        RECT 91.180 136.820 91.320 138.200 ;
        RECT 93.940 136.820 94.080 147.040 ;
        RECT 96.240 145.660 96.380 147.040 ;
        RECT 97.100 146.360 97.360 146.680 ;
        RECT 96.180 145.340 96.440 145.660 ;
        RECT 97.160 145.320 97.300 146.360 ;
        RECT 97.100 145.000 97.360 145.320 ;
        RECT 94.340 138.200 94.600 138.520 ;
        RECT 91.120 136.500 91.380 136.820 ;
        RECT 93.880 136.500 94.140 136.820 ;
        RECT 90.660 135.480 90.920 135.800 ;
        RECT 90.720 134.860 90.860 135.480 ;
        RECT 90.260 134.780 90.860 134.860 ;
        RECT 87.440 134.460 87.700 134.780 ;
        RECT 90.200 134.720 90.860 134.780 ;
        RECT 90.200 134.460 90.460 134.720 ;
        RECT 92.040 134.460 92.300 134.780 ;
        RECT 90.660 134.120 90.920 134.440 ;
        RECT 87.900 133.780 88.160 134.100 ;
        RECT 87.960 131.040 88.100 133.780 ;
        RECT 90.720 132.060 90.860 134.120 ;
        RECT 92.100 134.100 92.240 134.460 ;
        RECT 92.040 133.780 92.300 134.100 ;
        RECT 93.940 133.760 94.080 136.500 ;
        RECT 94.400 134.780 94.540 138.200 ;
        RECT 95.260 135.480 95.520 135.800 ;
        RECT 94.340 134.460 94.600 134.780 ;
        RECT 93.880 133.440 94.140 133.760 ;
        RECT 90.660 131.740 90.920 132.060 ;
        RECT 95.320 131.040 95.460 135.480 ;
        RECT 96.640 133.780 96.900 134.100 ;
        RECT 96.700 132.060 96.840 133.780 ;
        RECT 96.640 131.740 96.900 132.060 ;
        RECT 97.620 131.040 97.760 154.520 ;
        RECT 99.460 153.820 99.600 155.540 ;
        RECT 99.400 153.500 99.660 153.820 ;
        RECT 98.940 150.780 99.200 151.100 ;
        RECT 99.000 147.360 99.140 150.780 ;
        RECT 98.940 147.040 99.200 147.360 ;
        RECT 99.400 139.900 99.660 140.220 ;
        RECT 98.020 137.180 98.280 137.500 ;
        RECT 98.080 136.480 98.220 137.180 ;
        RECT 99.460 136.480 99.600 139.900 ;
        RECT 98.020 136.160 98.280 136.480 ;
        RECT 99.400 136.160 99.660 136.480 ;
        RECT 98.480 135.820 98.740 136.140 ;
        RECT 98.540 133.080 98.680 135.820 ;
        RECT 98.940 133.440 99.200 133.760 ;
        RECT 98.480 132.760 98.740 133.080 ;
        RECT 87.900 130.720 88.160 131.040 ;
        RECT 95.260 130.720 95.520 131.040 ;
        RECT 97.560 130.720 97.820 131.040 ;
        RECT 91.580 130.040 91.840 130.360 ;
        RECT 97.100 130.040 97.360 130.360 ;
        RECT 98.020 130.040 98.280 130.360 ;
        RECT 91.120 128.680 91.380 129.000 ;
        RECT 89.280 123.415 89.540 123.560 ;
        RECT 89.270 123.045 89.550 123.415 ;
        RECT 91.180 121.180 91.320 128.680 ;
        RECT 91.640 127.640 91.780 130.040 ;
        RECT 97.160 128.660 97.300 130.040 ;
        RECT 97.100 128.340 97.360 128.660 ;
        RECT 97.560 128.000 97.820 128.320 ;
        RECT 91.580 127.320 91.840 127.640 ;
        RECT 91.120 120.860 91.380 121.180 ;
        RECT 97.620 120.500 97.760 128.000 ;
        RECT 97.560 120.180 97.820 120.500 ;
        RECT 87.440 119.500 87.700 119.820 ;
        RECT 87.500 117.780 87.640 119.500 ;
        RECT 89.740 118.140 90.000 118.460 ;
        RECT 87.440 117.460 87.700 117.780 ;
        RECT 89.800 114.720 89.940 118.140 ;
        RECT 97.620 114.720 97.760 120.180 ;
        RECT 89.740 114.400 90.000 114.720 ;
        RECT 97.560 114.400 97.820 114.720 ;
        RECT 94.340 112.020 94.600 112.340 ;
        RECT 93.880 111.680 94.140 112.000 ;
        RECT 87.440 108.280 87.700 108.600 ;
        RECT 90.660 108.280 90.920 108.600 ;
        RECT 86.980 106.580 87.240 106.900 ;
        RECT 87.500 103.840 87.640 108.280 ;
        RECT 90.200 105.560 90.460 105.880 ;
        RECT 87.440 103.520 87.700 103.840 ;
        RECT 90.260 101.800 90.400 105.560 ;
        RECT 90.720 104.180 90.860 108.280 ;
        RECT 93.940 107.240 94.080 111.680 ;
        RECT 94.400 109.280 94.540 112.020 ;
        RECT 98.080 109.960 98.220 130.040 ;
        RECT 99.000 128.660 99.140 133.440 ;
        RECT 99.400 131.400 99.660 131.720 ;
        RECT 99.460 129.000 99.600 131.400 ;
        RECT 99.920 131.380 100.060 176.280 ;
        RECT 101.760 173.880 101.900 177.300 ;
        RECT 102.220 174.560 102.360 177.445 ;
        RECT 102.160 174.240 102.420 174.560 ;
        RECT 101.700 173.560 101.960 173.880 ;
        RECT 102.620 168.120 102.880 168.440 ;
        RECT 101.700 166.760 101.960 167.080 ;
        RECT 100.780 166.080 101.040 166.400 ;
        RECT 100.320 165.400 100.580 165.720 ;
        RECT 100.380 163.000 100.520 165.400 ;
        RECT 100.320 162.680 100.580 163.000 ;
        RECT 100.380 155.860 100.520 162.680 ;
        RECT 100.840 161.980 100.980 166.080 ;
        RECT 101.240 162.680 101.500 163.000 ;
        RECT 100.780 161.660 101.040 161.980 ;
        RECT 101.300 161.300 101.440 162.680 ;
        RECT 101.760 161.980 101.900 166.760 ;
        RECT 102.680 164.020 102.820 168.120 ;
        RECT 102.620 163.700 102.880 164.020 ;
        RECT 101.700 161.660 101.960 161.980 ;
        RECT 101.240 160.980 101.500 161.300 ;
        RECT 100.320 155.540 100.580 155.860 ;
        RECT 101.240 152.480 101.500 152.800 ;
        RECT 100.320 139.560 100.580 139.880 ;
        RECT 100.380 138.860 100.520 139.560 ;
        RECT 101.300 139.540 101.440 152.480 ;
        RECT 101.240 139.220 101.500 139.540 ;
        RECT 101.700 139.220 101.960 139.540 ;
        RECT 100.320 138.540 100.580 138.860 ;
        RECT 100.380 136.480 100.520 138.540 ;
        RECT 100.320 136.160 100.580 136.480 ;
        RECT 101.240 135.480 101.500 135.800 ;
        RECT 100.320 131.740 100.580 132.060 ;
        RECT 99.860 131.060 100.120 131.380 ;
        RECT 100.380 129.340 100.520 131.740 ;
        RECT 101.300 131.040 101.440 135.480 ;
        RECT 101.760 134.440 101.900 139.220 ;
        RECT 101.700 134.120 101.960 134.440 ;
        RECT 103.140 131.380 103.280 179.000 ;
        RECT 105.900 177.280 106.040 179.680 ;
        RECT 106.760 179.000 107.020 179.320 ;
        RECT 106.820 177.620 106.960 179.000 ;
        RECT 107.280 178.300 107.420 179.680 ;
        RECT 107.220 177.980 107.480 178.300 ;
        RECT 107.740 177.620 107.880 187.500 ;
        RECT 110.500 185.440 110.640 189.880 ;
        RECT 110.440 185.120 110.700 185.440 ;
        RECT 109.520 183.420 109.780 183.740 ;
        RECT 109.060 181.720 109.320 182.040 ;
        RECT 109.120 180.340 109.260 181.720 ;
        RECT 109.060 180.020 109.320 180.340 ;
        RECT 109.580 179.740 109.720 183.420 ;
        RECT 109.980 182.400 110.240 182.720 ;
        RECT 109.120 179.600 109.720 179.740 ;
        RECT 110.040 179.660 110.180 182.400 ;
        RECT 109.120 179.320 109.260 179.600 ;
        RECT 109.980 179.340 110.240 179.660 ;
        RECT 109.060 179.000 109.320 179.320 ;
        RECT 109.120 178.300 109.260 179.000 ;
        RECT 109.060 177.980 109.320 178.300 ;
        RECT 106.760 177.300 107.020 177.620 ;
        RECT 107.680 177.300 107.940 177.620 ;
        RECT 108.600 177.300 108.860 177.620 ;
        RECT 105.840 176.960 106.100 177.280 ;
        RECT 106.820 176.940 106.960 177.300 ;
        RECT 106.760 176.620 107.020 176.940 ;
        RECT 104.920 176.280 105.180 176.600 ;
        RECT 104.460 168.800 104.720 169.120 ;
        RECT 104.520 164.700 104.660 168.800 ;
        RECT 104.460 164.380 104.720 164.700 ;
        RECT 104.460 163.700 104.720 164.020 ;
        RECT 104.520 155.860 104.660 163.700 ;
        RECT 104.460 155.540 104.720 155.860 ;
        RECT 104.460 154.520 104.720 154.840 ;
        RECT 104.000 152.140 104.260 152.460 ;
        RECT 104.060 151.100 104.200 152.140 ;
        RECT 104.000 150.780 104.260 151.100 ;
        RECT 104.520 147.100 104.660 154.520 ;
        RECT 104.980 148.040 105.120 176.280 ;
        RECT 106.760 174.580 107.020 174.900 ;
        RECT 106.300 171.520 106.560 171.840 ;
        RECT 106.360 166.740 106.500 171.520 ;
        RECT 106.300 166.420 106.560 166.740 ;
        RECT 106.820 166.140 106.960 174.580 ;
        RECT 108.140 172.540 108.400 172.860 ;
        RECT 107.680 170.840 107.940 171.160 ;
        RECT 106.360 166.000 106.960 166.140 ;
        RECT 105.380 159.960 105.640 160.280 ;
        RECT 105.440 158.240 105.580 159.960 ;
        RECT 105.840 158.600 106.100 158.920 ;
        RECT 105.380 157.920 105.640 158.240 ;
        RECT 105.900 155.860 106.040 158.600 ;
        RECT 105.840 155.540 106.100 155.860 ;
        RECT 105.900 152.800 106.040 155.540 ;
        RECT 105.840 152.480 106.100 152.800 ;
        RECT 105.380 151.800 105.640 152.120 ;
        RECT 104.920 147.720 105.180 148.040 ;
        RECT 105.440 147.360 105.580 151.800 ;
        RECT 106.360 150.080 106.500 166.000 ;
        RECT 106.760 162.680 107.020 163.000 ;
        RECT 106.820 161.300 106.960 162.680 ;
        RECT 106.760 160.980 107.020 161.300 ;
        RECT 106.760 155.880 107.020 156.200 ;
        RECT 106.820 154.580 106.960 155.880 ;
        RECT 106.820 154.440 107.420 154.580 ;
        RECT 107.280 152.800 107.420 154.440 ;
        RECT 107.740 152.800 107.880 170.840 ;
        RECT 108.200 163.680 108.340 172.540 ;
        RECT 108.660 172.520 108.800 177.300 ;
        RECT 109.980 176.960 110.240 177.280 ;
        RECT 109.520 176.620 109.780 176.940 ;
        RECT 109.580 173.880 109.720 176.620 ;
        RECT 110.040 175.240 110.180 176.960 ;
        RECT 109.980 174.920 110.240 175.240 ;
        RECT 109.520 173.560 109.780 173.880 ;
        RECT 108.600 172.200 108.860 172.520 ;
        RECT 109.580 172.180 109.720 173.560 ;
        RECT 110.040 172.180 110.180 174.920 ;
        RECT 110.500 172.180 110.640 185.120 ;
        RECT 110.960 176.600 111.100 193.280 ;
        RECT 111.880 186.460 112.020 193.280 ;
        RECT 114.120 192.600 114.380 192.920 ;
        RECT 115.500 192.600 115.760 192.920 ;
        RECT 114.180 188.500 114.320 192.600 ;
        RECT 115.560 190.540 115.700 192.600 ;
        RECT 115.500 190.220 115.760 190.540 ;
        RECT 114.120 188.180 114.380 188.500 ;
        RECT 111.820 186.140 112.080 186.460 ;
        RECT 111.880 183.060 112.020 186.140 ;
        RECT 111.820 182.740 112.080 183.060 ;
        RECT 112.740 182.060 113.000 182.380 ;
        RECT 112.800 177.620 112.940 182.060 ;
        RECT 113.660 179.680 113.920 180.000 ;
        RECT 113.720 178.300 113.860 179.680 ;
        RECT 113.660 177.980 113.920 178.300 ;
        RECT 116.020 177.620 116.160 193.620 ;
        RECT 116.480 189.180 116.620 195.660 ;
        RECT 121.080 190.880 121.220 196.000 ;
        RECT 121.020 190.560 121.280 190.880 ;
        RECT 117.800 190.220 118.060 190.540 ;
        RECT 117.860 189.180 118.000 190.220 ;
        RECT 116.420 188.860 116.680 189.180 ;
        RECT 117.800 188.860 118.060 189.180 ;
        RECT 121.080 188.160 121.220 190.560 ;
        RECT 121.020 187.840 121.280 188.160 ;
        RECT 117.340 182.740 117.600 183.060 ;
        RECT 117.400 178.300 117.540 182.740 ;
        RECT 121.080 182.720 121.220 187.840 ;
        RECT 124.240 183.080 124.500 183.400 ;
        RECT 121.020 182.400 121.280 182.720 ;
        RECT 119.180 181.720 119.440 182.040 ;
        RECT 119.240 179.740 119.380 181.720 ;
        RECT 121.080 180.340 121.220 182.400 ;
        RECT 124.300 181.020 124.440 183.080 ;
        RECT 124.700 182.400 124.960 182.720 ;
        RECT 124.240 180.700 124.500 181.020 ;
        RECT 121.020 180.020 121.280 180.340 ;
        RECT 119.240 179.660 119.840 179.740 ;
        RECT 119.240 179.600 119.900 179.660 ;
        RECT 119.640 179.340 119.900 179.600 ;
        RECT 117.340 177.980 117.600 178.300 ;
        RECT 112.740 177.300 113.000 177.620 ;
        RECT 115.960 177.300 116.220 177.620 ;
        RECT 115.500 176.960 115.760 177.280 ;
        RECT 110.900 176.280 111.160 176.600 ;
        RECT 113.660 176.280 113.920 176.600 ;
        RECT 112.280 175.260 112.540 175.580 ;
        RECT 111.360 173.900 111.620 174.220 ;
        RECT 109.520 171.860 109.780 172.180 ;
        RECT 109.980 171.860 110.240 172.180 ;
        RECT 110.440 171.860 110.700 172.180 ;
        RECT 110.900 171.750 111.160 171.840 ;
        RECT 111.420 171.750 111.560 173.900 ;
        RECT 112.340 173.620 112.480 175.260 ;
        RECT 113.720 174.560 113.860 176.280 ;
        RECT 115.560 174.560 115.700 176.960 ;
        RECT 113.660 174.240 113.920 174.560 ;
        RECT 114.580 174.240 114.840 174.560 ;
        RECT 115.500 174.240 115.760 174.560 ;
        RECT 110.900 171.610 111.560 171.750 ;
        RECT 110.900 171.520 111.160 171.610 ;
        RECT 109.060 170.840 109.320 171.160 ;
        RECT 108.140 163.360 108.400 163.680 ;
        RECT 108.600 162.680 108.860 163.000 ;
        RECT 108.660 161.980 108.800 162.680 ;
        RECT 108.600 161.660 108.860 161.980 ;
        RECT 108.140 160.980 108.400 161.300 ;
        RECT 108.200 155.860 108.340 160.980 ;
        RECT 108.140 155.540 108.400 155.860 ;
        RECT 108.600 154.860 108.860 155.180 ;
        RECT 108.660 152.800 108.800 154.860 ;
        RECT 107.220 152.480 107.480 152.800 ;
        RECT 107.680 152.480 107.940 152.800 ;
        RECT 108.600 152.480 108.860 152.800 ;
        RECT 108.140 151.800 108.400 152.120 ;
        RECT 108.200 150.420 108.340 151.800 ;
        RECT 108.600 150.780 108.860 151.100 ;
        RECT 108.140 150.100 108.400 150.420 ;
        RECT 106.300 149.760 106.560 150.080 ;
        RECT 107.680 149.760 107.940 150.080 ;
        RECT 106.760 148.060 107.020 148.380 ;
        RECT 104.520 146.960 105.120 147.100 ;
        RECT 105.380 147.040 105.640 147.360 ;
        RECT 104.000 146.360 104.260 146.680 ;
        RECT 104.460 146.360 104.720 146.680 ;
        RECT 104.060 145.320 104.200 146.360 ;
        RECT 104.520 145.660 104.660 146.360 ;
        RECT 104.460 145.340 104.720 145.660 ;
        RECT 104.000 145.000 104.260 145.320 ;
        RECT 103.530 136.645 103.810 137.015 ;
        RECT 103.540 136.500 103.800 136.645 ;
        RECT 104.460 131.740 104.720 132.060 ;
        RECT 103.080 131.060 103.340 131.380 ;
        RECT 101.240 130.720 101.500 131.040 ;
        RECT 104.520 129.340 104.660 131.740 ;
        RECT 104.980 131.040 105.120 146.960 ;
        RECT 105.380 144.320 105.640 144.640 ;
        RECT 105.440 133.760 105.580 144.320 ;
        RECT 105.840 139.560 106.100 139.880 ;
        RECT 105.380 133.440 105.640 133.760 ;
        RECT 104.920 130.720 105.180 131.040 ;
        RECT 105.900 130.700 106.040 139.560 ;
        RECT 106.300 135.480 106.560 135.800 ;
        RECT 106.360 134.100 106.500 135.480 ;
        RECT 106.300 133.780 106.560 134.100 ;
        RECT 105.840 130.380 106.100 130.700 ;
        RECT 106.820 129.340 106.960 148.060 ;
        RECT 107.740 147.270 107.880 149.760 ;
        RECT 108.660 147.360 108.800 150.780 ;
        RECT 108.140 147.270 108.400 147.360 ;
        RECT 107.740 147.130 108.400 147.270 ;
        RECT 108.140 147.040 108.400 147.130 ;
        RECT 108.600 147.040 108.860 147.360 ;
        RECT 108.200 145.660 108.340 147.040 ;
        RECT 108.140 145.340 108.400 145.660 ;
        RECT 107.680 144.660 107.940 144.980 ;
        RECT 107.740 137.500 107.880 144.660 ;
        RECT 108.660 144.640 108.800 147.040 ;
        RECT 108.600 144.320 108.860 144.640 ;
        RECT 108.600 143.640 108.860 143.960 ;
        RECT 108.660 141.920 108.800 143.640 ;
        RECT 109.120 142.260 109.260 170.840 ;
        RECT 111.420 169.460 111.560 171.610 ;
        RECT 111.880 173.480 112.480 173.620 ;
        RECT 111.360 169.140 111.620 169.460 ;
        RECT 109.980 168.460 110.240 168.780 ;
        RECT 110.440 168.460 110.700 168.780 ;
        RECT 109.520 162.680 109.780 163.000 ;
        RECT 109.580 161.300 109.720 162.680 ;
        RECT 109.520 160.980 109.780 161.300 ;
        RECT 110.040 159.260 110.180 168.460 ;
        RECT 110.500 167.420 110.640 168.460 ;
        RECT 110.440 167.100 110.700 167.420 ;
        RECT 110.900 165.400 111.160 165.720 ;
        RECT 110.960 161.300 111.100 165.400 ;
        RECT 110.900 160.980 111.160 161.300 ;
        RECT 111.880 160.140 112.020 173.480 ;
        RECT 112.280 172.540 112.540 172.860 ;
        RECT 112.340 172.180 112.480 172.540 ;
        RECT 114.640 172.520 114.780 174.240 ;
        RECT 117.800 173.900 118.060 174.220 ;
        RECT 117.340 173.560 117.600 173.880 ;
        RECT 114.580 172.200 114.840 172.520 ;
        RECT 112.280 171.860 112.540 172.180 ;
        RECT 117.400 171.840 117.540 173.560 ;
        RECT 117.860 172.180 118.000 173.900 ;
        RECT 124.760 172.180 124.900 182.400 ;
        RECT 117.800 171.860 118.060 172.180 ;
        RECT 124.700 171.860 124.960 172.180 ;
        RECT 117.340 171.520 117.600 171.840 ;
        RECT 120.560 171.520 120.820 171.840 ;
        RECT 112.280 171.180 112.540 171.500 ;
        RECT 112.340 169.120 112.480 171.180 ;
        RECT 113.660 170.840 113.920 171.160 ;
        RECT 115.500 170.840 115.760 171.160 ;
        RECT 112.740 169.140 113.000 169.460 ;
        RECT 112.280 168.800 112.540 169.120 ;
        RECT 112.280 168.120 112.540 168.440 ;
        RECT 112.340 166.740 112.480 168.120 ;
        RECT 112.280 166.420 112.540 166.740 ;
        RECT 112.800 164.020 112.940 169.140 ;
        RECT 113.200 166.080 113.460 166.400 ;
        RECT 112.740 163.700 113.000 164.020 ;
        RECT 112.800 160.960 112.940 163.700 ;
        RECT 112.740 160.640 113.000 160.960 ;
        RECT 110.500 160.000 112.020 160.140 ;
        RECT 109.980 158.940 110.240 159.260 ;
        RECT 110.500 155.260 110.640 160.000 ;
        RECT 113.260 155.860 113.400 166.080 ;
        RECT 113.720 163.340 113.860 170.840 ;
        RECT 115.560 169.540 115.700 170.840 ;
        RECT 115.560 169.460 116.620 169.540 ;
        RECT 115.560 169.400 116.680 169.460 ;
        RECT 113.660 163.020 113.920 163.340 ;
        RECT 115.560 161.980 115.700 169.400 ;
        RECT 116.420 169.140 116.680 169.400 ;
        RECT 120.620 169.120 120.760 171.520 ;
        RECT 124.240 170.840 124.500 171.160 ;
        RECT 124.300 170.140 124.440 170.840 ;
        RECT 124.240 169.820 124.500 170.140 ;
        RECT 124.760 169.800 124.900 171.860 ;
        RECT 124.700 169.480 124.960 169.800 ;
        RECT 120.560 168.800 120.820 169.120 ;
        RECT 121.480 168.460 121.740 168.780 ;
        RECT 121.020 168.120 121.280 168.440 ;
        RECT 121.080 167.080 121.220 168.120 ;
        RECT 121.020 166.760 121.280 167.080 ;
        RECT 115.500 161.660 115.760 161.980 ;
        RECT 111.360 155.540 111.620 155.860 ;
        RECT 113.200 155.540 113.460 155.860 ;
        RECT 109.580 155.120 110.640 155.260 ;
        RECT 109.060 141.940 109.320 142.260 ;
        RECT 108.600 141.600 108.860 141.920 ;
        RECT 108.600 139.220 108.860 139.540 ;
        RECT 109.060 139.220 109.320 139.540 ;
        RECT 107.680 137.180 107.940 137.500 ;
        RECT 108.660 136.140 108.800 139.220 ;
        RECT 109.120 137.500 109.260 139.220 ;
        RECT 109.060 137.180 109.320 137.500 ;
        RECT 109.050 136.645 109.330 137.015 ;
        RECT 109.060 136.500 109.320 136.645 ;
        RECT 108.600 135.820 108.860 136.140 ;
        RECT 109.580 134.100 109.720 155.120 ;
        RECT 110.440 154.520 110.700 154.840 ;
        RECT 110.900 154.520 111.160 154.840 ;
        RECT 109.980 150.100 110.240 150.420 ;
        RECT 110.040 147.360 110.180 150.100 ;
        RECT 109.980 147.040 110.240 147.360 ;
        RECT 110.040 144.980 110.180 147.040 ;
        RECT 109.980 144.660 110.240 144.980 ;
        RECT 109.980 142.620 110.240 142.940 ;
        RECT 109.520 133.780 109.780 134.100 ;
        RECT 109.060 132.760 109.320 133.080 ;
        RECT 107.220 130.040 107.480 130.360 ;
        RECT 100.320 129.020 100.580 129.340 ;
        RECT 104.460 129.020 104.720 129.340 ;
        RECT 106.760 129.020 107.020 129.340 ;
        RECT 99.400 128.680 99.660 129.000 ;
        RECT 98.940 128.340 99.200 128.660 ;
        RECT 99.000 125.640 99.140 128.340 ;
        RECT 104.920 128.000 105.180 128.320 ;
        RECT 98.540 125.600 99.140 125.640 ;
        RECT 98.480 125.500 99.140 125.600 ;
        RECT 98.480 125.280 98.740 125.500 ;
        RECT 98.540 122.880 98.680 125.280 ;
        RECT 98.480 122.560 98.740 122.880 ;
        RECT 98.540 120.070 98.680 122.560 ;
        RECT 104.980 120.160 105.120 128.000 ;
        RECT 105.840 125.620 106.100 125.940 ;
        RECT 105.380 123.415 105.640 123.560 ;
        RECT 105.370 123.045 105.650 123.415 ;
        RECT 105.900 120.500 106.040 125.620 ;
        RECT 105.840 120.180 106.100 120.500 ;
        RECT 98.940 120.070 99.200 120.160 ;
        RECT 98.540 119.930 99.200 120.070 ;
        RECT 98.540 117.780 98.680 119.930 ;
        RECT 98.940 119.840 99.200 119.930 ;
        RECT 103.080 119.840 103.340 120.160 ;
        RECT 104.920 119.840 105.180 120.160 ;
        RECT 98.940 118.140 99.200 118.460 ;
        RECT 98.480 117.460 98.740 117.780 ;
        RECT 98.020 109.640 98.280 109.960 ;
        RECT 94.340 108.960 94.600 109.280 ;
        RECT 98.020 108.280 98.280 108.600 ;
        RECT 93.880 106.920 94.140 107.240 ;
        RECT 97.560 106.240 97.820 106.560 ;
        RECT 97.620 104.860 97.760 106.240 ;
        RECT 97.560 104.540 97.820 104.860 ;
        RECT 90.660 103.860 90.920 104.180 ;
        RECT 90.200 101.480 90.460 101.800 ;
        RECT 93.880 100.120 94.140 100.440 ;
        RECT 62.130 90.660 62.410 91.170 ;
        RECT 60.820 90.520 62.410 90.660 ;
        RECT 37.750 88.780 38.970 89.290 ;
        RECT 37.680 86.810 39.070 88.780 ;
        RECT 43.810 88.630 45.030 89.530 ;
        RECT 50.170 89.040 50.450 90.520 ;
        RECT 56.150 89.190 56.430 90.520 ;
        RECT 49.740 88.640 50.960 89.040 ;
        RECT 37.750 85.420 38.970 86.810 ;
        RECT 43.810 86.720 45.140 88.630 ;
        RECT 49.740 86.920 51.010 88.640 ;
        RECT 43.810 85.660 45.030 86.720 ;
        RECT 49.740 85.170 50.960 86.920 ;
        RECT 55.530 85.320 56.750 89.190 ;
        RECT 62.130 88.870 62.410 90.520 ;
        RECT 68.110 89.840 68.390 91.170 ;
        RECT 67.730 89.640 68.670 89.840 ;
        RECT 61.720 88.640 62.940 88.870 ;
        RECT 61.720 86.600 63.130 88.640 ;
        RECT 61.720 85.000 62.940 86.600 ;
        RECT 67.580 85.770 68.800 89.640 ;
        RECT 74.090 88.160 74.370 91.170 ;
        RECT 80.070 88.180 80.350 91.170 ;
        RECT 73.850 84.290 75.070 88.160 ;
        RECT 79.730 84.310 80.950 88.180 ;
        RECT 86.050 87.970 86.330 91.170 ;
        RECT 92.030 90.660 92.310 91.170 ;
        RECT 93.940 90.660 94.080 100.120 ;
        RECT 98.080 91.170 98.220 108.280 ;
        RECT 98.540 106.470 98.680 117.460 ;
        RECT 99.000 115.060 99.140 118.140 ;
        RECT 99.860 117.460 100.120 117.780 ;
        RECT 99.920 115.740 100.060 117.460 ;
        RECT 103.140 115.740 103.280 119.840 ;
        RECT 104.000 119.160 104.260 119.480 ;
        RECT 104.060 118.120 104.200 119.160 ;
        RECT 104.980 118.460 105.120 119.840 ;
        RECT 104.920 118.140 105.180 118.460 ;
        RECT 104.000 117.800 104.260 118.120 ;
        RECT 99.860 115.420 100.120 115.740 ;
        RECT 103.080 115.420 103.340 115.740 ;
        RECT 105.900 115.400 106.040 120.180 ;
        RECT 106.300 119.160 106.560 119.480 ;
        RECT 105.840 115.080 106.100 115.400 ;
        RECT 98.940 114.740 99.200 115.060 ;
        RECT 106.360 114.720 106.500 119.160 ;
        RECT 106.300 114.400 106.560 114.720 ;
        RECT 106.300 112.700 106.560 113.020 ;
        RECT 99.860 109.300 100.120 109.620 ;
        RECT 99.400 108.620 99.660 108.940 ;
        RECT 99.460 107.580 99.600 108.620 ;
        RECT 99.400 107.260 99.660 107.580 ;
        RECT 99.920 107.240 100.060 109.300 ;
        RECT 99.860 106.920 100.120 107.240 ;
        RECT 98.940 106.470 99.200 106.560 ;
        RECT 98.540 106.330 99.200 106.470 ;
        RECT 98.940 106.240 99.200 106.330 ;
        RECT 99.000 104.520 99.140 106.240 ;
        RECT 98.940 104.200 99.200 104.520 ;
        RECT 106.360 104.180 106.500 112.700 ;
        RECT 107.280 112.340 107.420 130.040 ;
        RECT 109.120 129.340 109.260 132.760 ;
        RECT 110.040 132.060 110.180 142.620 ;
        RECT 110.500 134.100 110.640 154.520 ;
        RECT 110.960 141.920 111.100 154.520 ;
        RECT 111.420 153.480 111.560 155.540 ;
        RECT 112.280 154.860 112.540 155.180 ;
        RECT 111.360 153.160 111.620 153.480 ;
        RECT 112.340 152.800 112.480 154.860 ;
        RECT 115.560 153.140 115.700 161.660 ;
        RECT 121.540 158.240 121.680 168.460 ;
        RECT 124.760 166.740 124.900 169.480 ;
        RECT 124.700 166.420 124.960 166.740 ;
        RECT 124.240 165.400 124.500 165.720 ;
        RECT 123.320 163.360 123.580 163.680 ;
        RECT 123.380 161.640 123.520 163.360 ;
        RECT 124.300 161.980 124.440 165.400 ;
        RECT 124.760 164.020 124.900 166.420 ;
        RECT 124.700 163.700 124.960 164.020 ;
        RECT 124.240 161.660 124.500 161.980 ;
        RECT 123.320 161.320 123.580 161.640 ;
        RECT 121.480 157.920 121.740 158.240 ;
        RECT 120.560 157.580 120.820 157.900 ;
        RECT 116.880 155.200 117.140 155.520 ;
        RECT 115.500 152.820 115.760 153.140 ;
        RECT 112.280 152.480 112.540 152.800 ;
        RECT 115.960 152.140 116.220 152.460 ;
        RECT 114.580 149.420 114.840 149.740 ;
        RECT 113.660 149.080 113.920 149.400 ;
        RECT 114.120 149.080 114.380 149.400 ;
        RECT 112.740 147.380 113.000 147.700 ;
        RECT 111.360 145.340 111.620 145.660 ;
        RECT 111.420 144.890 111.560 145.340 ;
        RECT 111.820 144.890 112.080 144.980 ;
        RECT 111.420 144.750 112.080 144.890 ;
        RECT 110.900 141.600 111.160 141.920 ;
        RECT 111.420 140.220 111.560 144.750 ;
        RECT 111.820 144.660 112.080 144.750 ;
        RECT 112.800 144.640 112.940 147.380 ;
        RECT 113.720 145.740 113.860 149.080 ;
        RECT 114.180 146.680 114.320 149.080 ;
        RECT 114.120 146.360 114.380 146.680 ;
        RECT 113.720 145.600 114.320 145.740 ;
        RECT 112.740 144.320 113.000 144.640 ;
        RECT 111.820 143.980 112.080 144.300 ;
        RECT 110.900 139.900 111.160 140.220 ;
        RECT 111.360 139.900 111.620 140.220 ;
        RECT 110.960 139.620 111.100 139.900 ;
        RECT 111.880 139.620 112.020 143.980 ;
        RECT 112.800 142.260 112.940 144.320 ;
        RECT 112.740 141.940 113.000 142.260 ;
        RECT 110.960 139.480 112.020 139.620 ;
        RECT 112.280 139.560 112.540 139.880 ;
        RECT 111.360 139.220 111.620 139.480 ;
        RECT 111.360 138.540 111.620 138.860 ;
        RECT 111.420 136.480 111.560 138.540 ;
        RECT 111.360 136.160 111.620 136.480 ;
        RECT 111.820 136.160 112.080 136.480 ;
        RECT 110.440 133.780 110.700 134.100 ;
        RECT 111.880 133.760 112.020 136.160 ;
        RECT 112.340 134.440 112.480 139.560 ;
        RECT 112.800 136.820 112.940 141.940 ;
        RECT 113.660 140.920 113.920 141.240 ;
        RECT 113.200 136.840 113.460 137.160 ;
        RECT 112.740 136.500 113.000 136.820 ;
        RECT 112.280 134.120 112.540 134.440 ;
        RECT 113.260 134.100 113.400 136.840 ;
        RECT 113.200 133.780 113.460 134.100 ;
        RECT 111.820 133.440 112.080 133.760 ;
        RECT 113.720 133.500 113.860 140.920 ;
        RECT 110.900 132.760 111.160 133.080 ;
        RECT 109.980 131.740 110.240 132.060 ;
        RECT 109.980 130.720 110.240 131.040 ;
        RECT 109.060 129.020 109.320 129.340 ;
        RECT 110.040 128.660 110.180 130.720 ;
        RECT 109.980 128.340 110.240 128.660 ;
        RECT 110.440 128.340 110.700 128.660 ;
        RECT 109.060 128.000 109.320 128.320 ;
        RECT 109.120 125.600 109.260 128.000 ;
        RECT 109.060 125.280 109.320 125.600 ;
        RECT 109.060 124.600 109.320 124.920 ;
        RECT 109.120 122.200 109.260 124.600 ;
        RECT 109.060 121.880 109.320 122.200 ;
        RECT 110.500 119.820 110.640 128.340 ;
        RECT 110.440 119.500 110.700 119.820 ;
        RECT 109.980 119.160 110.240 119.480 ;
        RECT 110.040 118.120 110.180 119.160 ;
        RECT 109.980 117.800 110.240 118.120 ;
        RECT 107.220 112.020 107.480 112.340 ;
        RECT 110.960 111.840 111.100 132.760 ;
        RECT 111.880 129.000 112.020 133.440 ;
        RECT 113.260 133.360 113.860 133.500 ;
        RECT 112.280 130.720 112.540 131.040 ;
        RECT 111.820 128.680 112.080 129.000 ;
        RECT 111.880 123.900 112.020 128.680 ;
        RECT 112.340 123.980 112.480 130.720 ;
        RECT 111.820 123.580 112.080 123.900 ;
        RECT 112.340 123.840 112.940 123.980 ;
        RECT 111.880 122.880 112.020 123.580 ;
        RECT 111.820 122.560 112.080 122.880 ;
        RECT 111.360 117.690 111.620 117.780 ;
        RECT 111.880 117.690 112.020 122.560 ;
        RECT 112.800 122.200 112.940 123.840 ;
        RECT 112.740 121.880 113.000 122.200 ;
        RECT 111.360 117.550 112.020 117.690 ;
        RECT 111.360 117.460 111.620 117.550 ;
        RECT 111.880 115.400 112.020 117.550 ;
        RECT 111.820 115.080 112.080 115.400 ;
        RECT 111.880 111.840 112.020 115.080 ;
        RECT 112.800 115.060 112.940 121.880 ;
        RECT 112.740 114.740 113.000 115.060 ;
        RECT 110.960 111.700 111.560 111.840 ;
        RECT 111.880 111.700 112.480 111.840 ;
        RECT 109.980 109.640 110.240 109.960 ;
        RECT 106.760 108.280 107.020 108.600 ;
        RECT 106.820 107.240 106.960 108.280 ;
        RECT 106.760 106.920 107.020 107.240 ;
        RECT 106.760 106.240 107.020 106.560 ;
        RECT 106.820 104.860 106.960 106.240 ;
        RECT 109.060 105.560 109.320 105.880 ;
        RECT 106.760 104.540 107.020 104.860 ;
        RECT 106.300 103.860 106.560 104.180 ;
        RECT 109.120 103.840 109.260 105.560 ;
        RECT 109.060 103.520 109.320 103.840 ;
        RECT 104.000 100.120 104.260 100.440 ;
        RECT 104.060 91.170 104.200 100.120 ;
        RECT 110.040 91.170 110.180 109.640 ;
        RECT 111.420 109.280 111.560 111.700 ;
        RECT 111.360 108.960 111.620 109.280 ;
        RECT 110.900 108.620 111.160 108.940 ;
        RECT 110.440 105.560 110.700 105.880 ;
        RECT 110.500 103.500 110.640 105.560 ;
        RECT 110.960 104.860 111.100 108.620 ;
        RECT 111.820 108.280 112.080 108.600 ;
        RECT 110.900 104.540 111.160 104.860 ;
        RECT 111.880 104.180 112.020 108.280 ;
        RECT 112.340 106.560 112.480 111.700 ;
        RECT 113.260 109.280 113.400 133.360 ;
        RECT 114.180 129.340 114.320 145.600 ;
        RECT 114.120 129.020 114.380 129.340 ;
        RECT 113.660 119.500 113.920 119.820 ;
        RECT 113.720 118.460 113.860 119.500 ;
        RECT 113.660 118.140 113.920 118.460 ;
        RECT 114.640 109.280 114.780 149.420 ;
        RECT 116.020 148.380 116.160 152.140 ;
        RECT 115.960 148.060 116.220 148.380 ;
        RECT 115.960 139.220 116.220 139.540 ;
        RECT 116.020 136.140 116.160 139.220 ;
        RECT 116.420 138.430 116.680 138.520 ;
        RECT 116.940 138.430 117.080 155.200 ;
        RECT 120.620 153.820 120.760 157.580 ;
        RECT 121.540 155.860 121.680 157.920 ;
        RECT 121.480 155.540 121.740 155.860 ;
        RECT 120.560 153.500 120.820 153.820 ;
        RECT 117.800 151.800 118.060 152.120 ;
        RECT 117.860 150.420 118.000 151.800 ;
        RECT 117.800 150.100 118.060 150.420 ;
        RECT 117.800 146.700 118.060 147.020 ;
        RECT 117.340 146.360 117.600 146.680 ;
        RECT 117.400 145.660 117.540 146.360 ;
        RECT 117.340 145.340 117.600 145.660 ;
        RECT 117.860 144.640 118.000 146.700 ;
        RECT 120.620 144.980 120.760 153.500 ;
        RECT 123.320 151.800 123.580 152.120 ;
        RECT 123.380 150.760 123.520 151.800 ;
        RECT 123.320 150.440 123.580 150.760 ;
        RECT 126.080 149.760 126.340 150.080 ;
        RECT 126.140 147.360 126.280 149.760 ;
        RECT 123.780 147.040 124.040 147.360 ;
        RECT 125.160 147.040 125.420 147.360 ;
        RECT 126.080 147.040 126.340 147.360 ;
        RECT 121.020 146.700 121.280 147.020 ;
        RECT 121.080 145.660 121.220 146.700 ;
        RECT 123.840 145.660 123.980 147.040 ;
        RECT 121.020 145.340 121.280 145.660 ;
        RECT 123.780 145.340 124.040 145.660 ;
        RECT 120.560 144.660 120.820 144.980 ;
        RECT 117.800 144.320 118.060 144.640 ;
        RECT 117.860 141.920 118.000 144.320 ;
        RECT 120.620 141.920 120.760 144.660 ;
        RECT 124.700 142.280 124.960 142.600 ;
        RECT 117.800 141.600 118.060 141.920 ;
        RECT 120.560 141.660 120.820 141.920 ;
        RECT 120.560 141.600 121.220 141.660 ;
        RECT 120.620 141.520 121.220 141.600 ;
        RECT 117.340 140.920 117.600 141.240 ;
        RECT 120.560 140.920 120.820 141.240 ;
        RECT 117.400 138.860 117.540 140.920 ;
        RECT 120.620 139.880 120.760 140.920 ;
        RECT 121.080 140.220 121.220 141.520 ;
        RECT 121.020 139.900 121.280 140.220 ;
        RECT 120.560 139.560 120.820 139.880 ;
        RECT 124.240 138.880 124.500 139.200 ;
        RECT 117.340 138.540 117.600 138.860 ;
        RECT 116.420 138.290 117.080 138.430 ;
        RECT 116.420 138.200 116.680 138.290 ;
        RECT 115.960 135.820 116.220 136.140 ;
        RECT 116.940 128.660 117.080 138.290 ;
        RECT 124.300 137.500 124.440 138.880 ;
        RECT 124.240 137.180 124.500 137.500 ;
        RECT 124.760 136.480 124.900 142.280 ;
        RECT 121.020 136.160 121.280 136.480 ;
        RECT 124.700 136.160 124.960 136.480 ;
        RECT 121.080 134.780 121.220 136.160 ;
        RECT 121.020 134.460 121.280 134.780 ;
        RECT 116.420 128.340 116.680 128.660 ;
        RECT 116.880 128.340 117.140 128.660 ;
        RECT 115.040 128.000 115.300 128.320 ;
        RECT 115.100 126.620 115.240 128.000 ;
        RECT 115.040 126.300 115.300 126.620 ;
        RECT 116.480 125.260 116.620 128.340 ;
        RECT 116.420 124.940 116.680 125.260 ;
        RECT 116.940 120.160 117.080 128.340 ;
        RECT 118.720 127.320 118.980 127.640 ;
        RECT 121.020 127.320 121.280 127.640 ;
        RECT 118.780 125.260 118.920 127.320 ;
        RECT 121.080 125.940 121.220 127.320 ;
        RECT 121.020 125.620 121.280 125.940 ;
        RECT 124.700 125.280 124.960 125.600 ;
        RECT 118.720 124.940 118.980 125.260 ;
        RECT 120.560 124.600 120.820 124.920 ;
        RECT 119.180 123.240 119.440 123.560 ;
        RECT 118.260 122.560 118.520 122.880 ;
        RECT 118.320 120.500 118.460 122.560 ;
        RECT 119.240 121.180 119.380 123.240 ;
        RECT 119.180 120.860 119.440 121.180 ;
        RECT 118.260 120.180 118.520 120.500 ;
        RECT 120.620 120.160 120.760 124.600 ;
        RECT 124.240 122.900 124.500 123.220 ;
        RECT 124.300 121.180 124.440 122.900 ;
        RECT 124.760 122.880 124.900 125.280 ;
        RECT 124.700 122.560 124.960 122.880 ;
        RECT 124.240 120.860 124.500 121.180 ;
        RECT 116.420 119.840 116.680 120.160 ;
        RECT 116.880 119.840 117.140 120.160 ;
        RECT 120.560 119.840 120.820 120.160 ;
        RECT 116.480 118.460 116.620 119.840 ;
        RECT 116.420 118.140 116.680 118.460 ;
        RECT 116.940 118.120 117.080 119.840 ;
        RECT 116.880 117.800 117.140 118.120 ;
        RECT 115.500 117.460 115.760 117.780 ;
        RECT 117.340 117.460 117.600 117.780 ;
        RECT 115.560 115.740 115.700 117.460 ;
        RECT 115.500 115.420 115.760 115.740 ;
        RECT 115.500 114.060 115.760 114.380 ;
        RECT 115.560 110.300 115.700 114.060 ;
        RECT 117.400 110.300 117.540 117.460 ;
        RECT 124.240 114.400 124.500 114.720 ;
        RECT 120.560 111.000 120.820 111.320 ;
        RECT 115.500 109.980 115.760 110.300 ;
        RECT 117.340 109.980 117.600 110.300 ;
        RECT 113.200 108.960 113.460 109.280 ;
        RECT 114.580 108.960 114.840 109.280 ;
        RECT 115.960 108.960 116.220 109.280 ;
        RECT 116.020 107.580 116.160 108.960 ;
        RECT 115.960 107.260 116.220 107.580 ;
        RECT 112.280 106.240 112.540 106.560 ;
        RECT 120.100 106.240 120.360 106.560 ;
        RECT 115.040 105.560 115.300 105.880 ;
        RECT 111.820 103.860 112.080 104.180 ;
        RECT 110.440 103.180 110.700 103.500 ;
        RECT 110.900 102.840 111.160 103.160 ;
        RECT 110.960 101.800 111.100 102.840 ;
        RECT 115.100 101.800 115.240 105.560 ;
        RECT 120.160 104.180 120.300 106.240 ;
        RECT 120.100 103.860 120.360 104.180 ;
        RECT 110.900 101.480 111.160 101.800 ;
        RECT 115.040 101.480 115.300 101.800 ;
        RECT 115.960 100.120 116.220 100.440 ;
        RECT 116.020 91.170 116.160 100.120 ;
        RECT 92.030 90.520 94.080 90.660 ;
        RECT 92.030 88.370 92.310 90.520 ;
        RECT 98.010 88.500 98.290 91.170 ;
        RECT 103.990 88.610 104.270 91.170 ;
        RECT 109.970 89.290 110.250 91.170 ;
        RECT 115.950 89.570 116.230 91.170 ;
        RECT 120.620 90.660 120.760 111.000 ;
        RECT 121.020 108.280 121.280 108.600 ;
        RECT 121.080 107.240 121.220 108.280 ;
        RECT 124.300 107.580 124.440 114.400 ;
        RECT 125.220 112.340 125.360 147.040 ;
        RECT 126.140 139.200 126.280 147.040 ;
        RECT 126.080 138.880 126.340 139.200 ;
        RECT 126.140 136.820 126.280 138.880 ;
        RECT 126.080 136.500 126.340 136.820 ;
        RECT 127.920 117.120 128.180 117.440 ;
        RECT 126.080 113.720 126.340 114.040 ;
        RECT 126.140 112.680 126.280 113.720 ;
        RECT 126.080 112.360 126.340 112.680 ;
        RECT 125.160 112.020 125.420 112.340 ;
        RECT 124.700 111.000 124.960 111.320 ;
        RECT 124.760 109.620 124.900 111.000 ;
        RECT 124.700 109.300 124.960 109.620 ;
        RECT 126.080 108.960 126.340 109.280 ;
        RECT 124.240 107.260 124.500 107.580 ;
        RECT 121.020 106.920 121.280 107.240 ;
        RECT 126.140 106.560 126.280 108.960 ;
        RECT 126.080 106.240 126.340 106.560 ;
        RECT 125.160 102.840 125.420 103.160 ;
        RECT 125.220 101.460 125.360 102.840 ;
        RECT 125.160 101.140 125.420 101.460 ;
        RECT 127.980 91.170 128.120 117.120 ;
        RECT 121.930 90.660 122.210 91.170 ;
        RECT 120.620 90.520 122.210 90.660 ;
        RECT 121.930 89.570 122.210 90.520 ;
        RECT 74.090 80.440 74.370 84.290 ;
        RECT 20.140 80.160 74.370 80.440 ;
        RECT 20.140 75.650 20.420 80.160 ;
        RECT 80.070 79.800 80.350 84.310 ;
        RECT 85.470 84.100 86.690 87.970 ;
        RECT 91.460 84.500 92.680 88.370 ;
        RECT 97.600 84.630 98.820 88.500 ;
        RECT 103.650 84.740 104.870 88.610 ;
        RECT 109.620 85.420 110.840 89.290 ;
        RECT 115.740 85.700 116.960 89.570 ;
        RECT 121.520 85.700 122.740 89.570 ;
        RECT 127.910 89.380 128.190 91.170 ;
        RECT 31.380 79.520 80.350 79.800 ;
        RECT 31.380 75.850 31.660 79.520 ;
        RECT 86.050 79.170 86.330 84.100 ;
        RECT 42.510 78.890 86.330 79.170 ;
        RECT 19.330 73.120 21.890 75.650 ;
        RECT 28.185 73.180 30.255 74.460 ;
        RECT 30.670 73.320 33.230 75.850 ;
        RECT 42.510 75.750 42.790 78.890 ;
        RECT 92.030 78.570 92.310 84.500 ;
        RECT 53.830 78.290 92.310 78.570 ;
        RECT 53.830 75.820 54.110 78.290 ;
        RECT 98.010 77.990 98.290 84.630 ;
        RECT 64.900 77.710 98.290 77.990 ;
        RECT 20.145 70.600 20.555 73.120 ;
        RECT 31.345 70.610 31.755 73.320 ;
        RECT 39.475 73.150 41.545 74.430 ;
        RECT 41.910 73.220 44.470 75.750 ;
        RECT 20.165 49.090 20.555 70.600 ;
        RECT 26.485 63.200 26.755 65.240 ;
        RECT 27.615 63.200 27.885 65.200 ;
        RECT 26.485 56.510 27.885 63.200 ;
        RECT 26.485 55.190 26.755 56.510 ;
        RECT 27.615 55.150 27.885 56.510 ;
        RECT 28.885 55.260 29.205 65.190 ;
        RECT 28.885 55.200 29.215 55.260 ;
        RECT 26.405 54.290 27.535 54.300 ;
        RECT 28.895 54.290 29.215 55.200 ;
        RECT 25.765 53.490 26.125 54.110 ;
        RECT 25.845 52.610 26.105 53.490 ;
        RECT 26.385 53.240 29.215 54.290 ;
        RECT 25.675 52.230 26.205 52.610 ;
        RECT 26.405 52.020 27.535 53.240 ;
        RECT 28.895 53.220 29.215 53.240 ;
        RECT 22.205 50.990 22.475 51.940 ;
        RECT 22.205 50.840 22.675 50.990 ;
        RECT 22.205 50.160 22.765 50.840 ;
        RECT 22.285 50.150 22.765 50.160 ;
        RECT 21.575 49.620 22.195 49.980 ;
        RECT 21.615 49.090 22.045 49.620 ;
        RECT 20.165 48.670 22.045 49.090 ;
        RECT 22.535 48.960 22.765 50.150 ;
        RECT 21.615 47.800 22.045 48.670 ;
        RECT 22.455 48.360 22.835 48.960 ;
        RECT 21.435 47.440 22.055 47.800 ;
        RECT 22.055 46.990 22.325 47.240 ;
        RECT 22.535 46.990 22.765 48.360 ;
        RECT 22.055 46.880 22.765 46.990 ;
        RECT 26.235 47.780 27.615 52.020 ;
        RECT 31.365 49.100 31.755 70.610 ;
        RECT 42.565 70.580 42.975 73.220 ;
        RECT 50.055 73.090 52.125 74.370 ;
        RECT 53.150 73.290 55.710 75.820 ;
        RECT 64.900 75.810 65.180 77.710 ;
        RECT 103.990 77.230 104.270 84.740 ;
        RECT 76.140 76.950 104.270 77.230 ;
        RECT 37.685 63.210 37.955 65.250 ;
        RECT 38.815 63.210 39.085 65.210 ;
        RECT 37.685 56.520 39.085 63.210 ;
        RECT 37.685 55.200 37.955 56.520 ;
        RECT 38.815 55.160 39.085 56.520 ;
        RECT 40.085 55.270 40.405 65.200 ;
        RECT 40.085 55.210 40.415 55.270 ;
        RECT 37.605 54.300 38.735 54.310 ;
        RECT 40.095 54.300 40.415 55.210 ;
        RECT 36.965 53.500 37.325 54.120 ;
        RECT 37.045 52.620 37.305 53.500 ;
        RECT 37.585 53.250 40.415 54.300 ;
        RECT 36.875 52.240 37.405 52.620 ;
        RECT 37.605 52.030 38.735 53.250 ;
        RECT 40.095 53.230 40.415 53.250 ;
        RECT 33.405 51.000 33.675 51.950 ;
        RECT 33.405 50.850 33.875 51.000 ;
        RECT 33.405 50.170 33.965 50.850 ;
        RECT 33.485 50.160 33.965 50.170 ;
        RECT 32.775 49.630 33.395 49.990 ;
        RECT 32.815 49.100 33.245 49.630 ;
        RECT 31.365 48.680 33.245 49.100 ;
        RECT 33.735 48.970 33.965 50.160 ;
        RECT 32.815 47.810 33.245 48.680 ;
        RECT 33.655 48.370 34.035 48.970 ;
        RECT 26.235 46.920 26.535 47.780 ;
        RECT 27.315 46.920 27.615 47.780 ;
        RECT 32.635 47.450 33.255 47.810 ;
        RECT 33.255 47.000 33.525 47.250 ;
        RECT 33.735 47.000 33.965 48.370 ;
        RECT 33.255 46.890 33.965 47.000 ;
        RECT 37.435 47.790 38.815 52.030 ;
        RECT 42.585 49.070 42.975 70.580 ;
        RECT 53.815 70.560 54.225 73.290 ;
        RECT 61.475 73.120 63.545 74.400 ;
        RECT 64.400 73.280 66.960 75.810 ;
        RECT 76.140 75.740 76.420 76.950 ;
        RECT 109.970 76.610 110.250 85.420 ;
        RECT 87.580 76.330 110.250 76.610 ;
        RECT 87.580 75.760 87.860 76.330 ;
        RECT 115.950 76.030 116.230 85.700 ;
        RECT 98.850 75.840 116.230 76.030 ;
        RECT 48.905 63.180 49.175 65.220 ;
        RECT 50.035 63.180 50.305 65.180 ;
        RECT 48.905 56.490 50.305 63.180 ;
        RECT 48.905 55.170 49.175 56.490 ;
        RECT 50.035 55.130 50.305 56.490 ;
        RECT 51.305 55.240 51.625 65.170 ;
        RECT 51.305 55.180 51.635 55.240 ;
        RECT 48.825 54.270 49.955 54.280 ;
        RECT 51.315 54.270 51.635 55.180 ;
        RECT 48.185 53.470 48.545 54.090 ;
        RECT 48.265 52.590 48.525 53.470 ;
        RECT 48.805 53.220 51.635 54.270 ;
        RECT 48.095 52.210 48.625 52.590 ;
        RECT 48.825 52.000 49.955 53.220 ;
        RECT 51.315 53.200 51.635 53.220 ;
        RECT 44.625 50.970 44.895 51.920 ;
        RECT 44.625 50.820 45.095 50.970 ;
        RECT 44.625 50.140 45.185 50.820 ;
        RECT 44.705 50.130 45.185 50.140 ;
        RECT 43.995 49.600 44.615 49.960 ;
        RECT 44.035 49.070 44.465 49.600 ;
        RECT 42.585 48.650 44.465 49.070 ;
        RECT 44.955 48.940 45.185 50.130 ;
        RECT 37.435 46.930 37.735 47.790 ;
        RECT 38.515 46.930 38.815 47.790 ;
        RECT 44.035 47.780 44.465 48.650 ;
        RECT 44.875 48.340 45.255 48.940 ;
        RECT 43.855 47.420 44.475 47.780 ;
        RECT 44.475 46.970 44.745 47.220 ;
        RECT 44.955 46.970 45.185 48.340 ;
        RECT 22.055 46.570 22.715 46.880 ;
        RECT 22.055 46.400 22.325 46.570 ;
        RECT 27.565 46.380 28.045 46.760 ;
        RECT 33.255 46.580 33.915 46.890 ;
        RECT 44.475 46.860 45.185 46.970 ;
        RECT 48.655 47.760 50.035 52.000 ;
        RECT 53.835 49.050 54.225 70.560 ;
        RECT 65.035 70.550 65.445 73.280 ;
        RECT 72.585 73.130 74.655 74.410 ;
        RECT 75.550 73.210 78.110 75.740 ;
        RECT 60.155 63.160 60.425 65.200 ;
        RECT 61.285 63.160 61.555 65.160 ;
        RECT 60.155 56.470 61.555 63.160 ;
        RECT 60.155 55.150 60.425 56.470 ;
        RECT 61.285 55.110 61.555 56.470 ;
        RECT 62.555 55.220 62.875 65.150 ;
        RECT 62.555 55.160 62.885 55.220 ;
        RECT 60.075 54.250 61.205 54.260 ;
        RECT 62.565 54.250 62.885 55.160 ;
        RECT 59.435 53.450 59.795 54.070 ;
        RECT 59.515 52.570 59.775 53.450 ;
        RECT 60.055 53.200 62.885 54.250 ;
        RECT 59.345 52.190 59.875 52.570 ;
        RECT 60.075 51.980 61.205 53.200 ;
        RECT 62.565 53.180 62.885 53.200 ;
        RECT 55.875 50.950 56.145 51.900 ;
        RECT 55.875 50.800 56.345 50.950 ;
        RECT 55.875 50.120 56.435 50.800 ;
        RECT 55.955 50.110 56.435 50.120 ;
        RECT 55.245 49.580 55.865 49.940 ;
        RECT 55.285 49.050 55.715 49.580 ;
        RECT 53.835 48.630 55.715 49.050 ;
        RECT 56.205 48.920 56.435 50.110 ;
        RECT 55.285 47.760 55.715 48.630 ;
        RECT 56.125 48.320 56.505 48.920 ;
        RECT 48.655 46.900 48.955 47.760 ;
        RECT 49.735 46.900 50.035 47.760 ;
        RECT 55.105 47.400 55.725 47.760 ;
        RECT 55.725 46.950 55.995 47.200 ;
        RECT 56.205 46.950 56.435 48.320 ;
        RECT 33.255 46.410 33.525 46.580 ;
        RECT 38.765 46.390 39.245 46.770 ;
        RECT 44.475 46.550 45.135 46.860 ;
        RECT 55.725 46.840 56.435 46.950 ;
        RECT 59.905 47.740 61.285 51.980 ;
        RECT 65.055 49.040 65.445 70.550 ;
        RECT 76.275 70.540 76.685 73.210 ;
        RECT 83.855 73.120 85.925 74.400 ;
        RECT 86.850 73.230 89.410 75.760 ;
        RECT 98.150 75.750 116.230 75.840 ;
        RECT 87.525 70.550 87.935 73.230 ;
        RECT 95.045 73.060 97.115 74.340 ;
        RECT 98.150 73.310 100.710 75.750 ;
        RECT 109.390 75.480 111.950 75.560 ;
        RECT 121.930 75.480 122.210 85.700 ;
        RECT 127.550 85.510 128.770 89.380 ;
        RECT 127.910 76.040 128.190 85.510 ;
        RECT 109.390 75.200 122.210 75.480 ;
        RECT 71.375 63.150 71.645 65.190 ;
        RECT 72.505 63.150 72.775 65.150 ;
        RECT 71.375 56.460 72.775 63.150 ;
        RECT 71.375 55.140 71.645 56.460 ;
        RECT 72.505 55.100 72.775 56.460 ;
        RECT 73.775 55.210 74.095 65.140 ;
        RECT 73.775 55.150 74.105 55.210 ;
        RECT 71.295 54.240 72.425 54.250 ;
        RECT 73.785 54.240 74.105 55.150 ;
        RECT 70.655 53.440 71.015 54.060 ;
        RECT 70.735 52.560 70.995 53.440 ;
        RECT 71.275 53.190 74.105 54.240 ;
        RECT 70.565 52.180 71.095 52.560 ;
        RECT 71.295 51.970 72.425 53.190 ;
        RECT 73.785 53.170 74.105 53.190 ;
        RECT 67.095 50.940 67.365 51.890 ;
        RECT 67.095 50.790 67.565 50.940 ;
        RECT 67.095 50.110 67.655 50.790 ;
        RECT 67.175 50.100 67.655 50.110 ;
        RECT 66.465 49.570 67.085 49.930 ;
        RECT 66.505 49.040 66.935 49.570 ;
        RECT 65.055 48.620 66.935 49.040 ;
        RECT 67.425 48.910 67.655 50.100 ;
        RECT 66.505 47.750 66.935 48.620 ;
        RECT 67.345 48.310 67.725 48.910 ;
        RECT 59.905 46.880 60.205 47.740 ;
        RECT 60.985 46.880 61.285 47.740 ;
        RECT 66.325 47.390 66.945 47.750 ;
        RECT 66.945 46.940 67.215 47.190 ;
        RECT 67.425 46.940 67.655 48.310 ;
        RECT 27.665 45.760 27.915 46.380 ;
        RECT 38.865 45.770 39.115 46.390 ;
        RECT 44.475 46.380 44.745 46.550 ;
        RECT 49.985 46.360 50.465 46.740 ;
        RECT 55.725 46.530 56.385 46.840 ;
        RECT 66.945 46.830 67.655 46.940 ;
        RECT 71.125 47.730 72.505 51.970 ;
        RECT 76.295 49.030 76.685 70.540 ;
        RECT 82.615 63.140 82.885 65.180 ;
        RECT 83.745 63.140 84.015 65.140 ;
        RECT 82.615 56.450 84.015 63.140 ;
        RECT 82.615 55.130 82.885 56.450 ;
        RECT 83.745 55.090 84.015 56.450 ;
        RECT 85.015 55.200 85.335 65.130 ;
        RECT 85.015 55.140 85.345 55.200 ;
        RECT 82.535 54.230 83.665 54.240 ;
        RECT 85.025 54.230 85.345 55.140 ;
        RECT 81.895 53.430 82.255 54.050 ;
        RECT 81.975 52.550 82.235 53.430 ;
        RECT 82.515 53.180 85.345 54.230 ;
        RECT 81.805 52.170 82.335 52.550 ;
        RECT 82.535 51.960 83.665 53.180 ;
        RECT 85.025 53.160 85.345 53.180 ;
        RECT 78.335 50.930 78.605 51.880 ;
        RECT 78.335 50.780 78.805 50.930 ;
        RECT 78.335 50.100 78.895 50.780 ;
        RECT 78.415 50.090 78.895 50.100 ;
        RECT 77.705 49.560 78.325 49.920 ;
        RECT 77.745 49.030 78.175 49.560 ;
        RECT 76.295 48.610 78.175 49.030 ;
        RECT 78.665 48.900 78.895 50.090 ;
        RECT 77.745 47.740 78.175 48.610 ;
        RECT 78.585 48.300 78.965 48.900 ;
        RECT 71.125 46.870 71.425 47.730 ;
        RECT 72.205 46.870 72.505 47.730 ;
        RECT 77.565 47.380 78.185 47.740 ;
        RECT 78.185 46.930 78.455 47.180 ;
        RECT 78.665 46.930 78.895 48.300 ;
        RECT 55.725 46.360 55.995 46.530 ;
        RECT 27.565 45.160 27.945 45.760 ;
        RECT 38.765 45.170 39.145 45.770 ;
        RECT 50.085 45.740 50.335 46.360 ;
        RECT 61.235 46.340 61.715 46.720 ;
        RECT 66.945 46.520 67.605 46.830 ;
        RECT 78.185 46.820 78.895 46.930 ;
        RECT 82.365 47.720 83.745 51.960 ;
        RECT 87.545 49.040 87.935 70.550 ;
        RECT 98.805 70.540 99.215 73.310 ;
        RECT 106.455 73.110 108.525 74.390 ;
        RECT 109.390 73.030 111.950 75.200 ;
        RECT 125.760 74.810 128.190 76.040 ;
        RECT 121.290 74.790 128.190 74.810 ;
        RECT 120.600 74.530 128.190 74.790 ;
        RECT 117.655 73.110 119.725 74.390 ;
        RECT 120.600 73.180 128.160 74.530 ;
        RECT 129.505 73.190 131.575 74.470 ;
        RECT 120.600 73.110 126.160 73.180 ;
        RECT 110.075 70.540 110.485 73.030 ;
        RECT 121.325 70.540 121.735 73.110 ;
        RECT 93.865 63.150 94.135 65.190 ;
        RECT 94.995 63.150 95.265 65.150 ;
        RECT 93.865 56.460 95.265 63.150 ;
        RECT 93.865 55.140 94.135 56.460 ;
        RECT 94.995 55.100 95.265 56.460 ;
        RECT 96.265 55.210 96.585 65.140 ;
        RECT 96.265 55.150 96.595 55.210 ;
        RECT 93.785 54.240 94.915 54.250 ;
        RECT 96.275 54.240 96.595 55.150 ;
        RECT 93.145 53.440 93.505 54.060 ;
        RECT 93.225 52.560 93.485 53.440 ;
        RECT 93.765 53.190 96.595 54.240 ;
        RECT 93.055 52.180 93.585 52.560 ;
        RECT 93.785 51.970 94.915 53.190 ;
        RECT 96.275 53.170 96.595 53.190 ;
        RECT 89.585 50.940 89.855 51.890 ;
        RECT 89.585 50.790 90.055 50.940 ;
        RECT 89.585 50.110 90.145 50.790 ;
        RECT 89.665 50.100 90.145 50.110 ;
        RECT 88.955 49.570 89.575 49.930 ;
        RECT 88.995 49.040 89.425 49.570 ;
        RECT 87.545 48.620 89.425 49.040 ;
        RECT 89.915 48.910 90.145 50.100 ;
        RECT 88.995 47.750 89.425 48.620 ;
        RECT 89.835 48.310 90.215 48.910 ;
        RECT 82.365 46.860 82.665 47.720 ;
        RECT 83.445 46.860 83.745 47.720 ;
        RECT 88.815 47.390 89.435 47.750 ;
        RECT 89.435 46.940 89.705 47.190 ;
        RECT 89.915 46.940 90.145 48.310 ;
        RECT 89.435 46.830 90.145 46.940 ;
        RECT 93.615 47.730 94.995 51.970 ;
        RECT 98.825 49.030 99.215 70.540 ;
        RECT 105.145 63.140 105.415 65.180 ;
        RECT 106.275 63.140 106.545 65.140 ;
        RECT 105.145 56.450 106.545 63.140 ;
        RECT 105.145 55.130 105.415 56.450 ;
        RECT 106.275 55.090 106.545 56.450 ;
        RECT 107.545 55.200 107.865 65.130 ;
        RECT 107.545 55.140 107.875 55.200 ;
        RECT 105.065 54.230 106.195 54.240 ;
        RECT 107.555 54.230 107.875 55.140 ;
        RECT 104.425 53.430 104.785 54.050 ;
        RECT 104.505 52.550 104.765 53.430 ;
        RECT 105.045 53.180 107.875 54.230 ;
        RECT 104.335 52.170 104.865 52.550 ;
        RECT 105.065 51.960 106.195 53.180 ;
        RECT 107.555 53.160 107.875 53.180 ;
        RECT 100.865 50.930 101.135 51.880 ;
        RECT 100.865 50.780 101.335 50.930 ;
        RECT 100.865 50.100 101.425 50.780 ;
        RECT 100.945 50.090 101.425 50.100 ;
        RECT 100.235 49.560 100.855 49.920 ;
        RECT 100.275 49.030 100.705 49.560 ;
        RECT 98.825 48.610 100.705 49.030 ;
        RECT 101.195 48.900 101.425 50.090 ;
        RECT 100.275 47.740 100.705 48.610 ;
        RECT 101.115 48.300 101.495 48.900 ;
        RECT 93.615 46.870 93.915 47.730 ;
        RECT 94.695 46.870 94.995 47.730 ;
        RECT 100.095 47.380 100.715 47.740 ;
        RECT 100.715 46.930 100.985 47.180 ;
        RECT 101.195 46.930 101.425 48.300 ;
        RECT 66.945 46.350 67.215 46.520 ;
        RECT 49.985 45.140 50.365 45.740 ;
        RECT 61.335 45.720 61.585 46.340 ;
        RECT 72.455 46.330 72.935 46.710 ;
        RECT 78.185 46.510 78.845 46.820 ;
        RECT 78.185 46.340 78.455 46.510 ;
        RECT 61.235 45.120 61.615 45.720 ;
        RECT 72.555 45.710 72.805 46.330 ;
        RECT 83.695 46.320 84.175 46.700 ;
        RECT 89.435 46.520 90.095 46.830 ;
        RECT 100.715 46.820 101.425 46.930 ;
        RECT 104.895 47.720 106.275 51.960 ;
        RECT 110.095 49.030 110.485 70.540 ;
        RECT 116.415 63.140 116.685 65.180 ;
        RECT 117.545 63.140 117.815 65.140 ;
        RECT 116.415 56.450 117.815 63.140 ;
        RECT 116.415 55.130 116.685 56.450 ;
        RECT 117.545 55.090 117.815 56.450 ;
        RECT 118.815 55.200 119.135 65.130 ;
        RECT 118.815 55.140 119.145 55.200 ;
        RECT 116.335 54.230 117.465 54.240 ;
        RECT 118.825 54.230 119.145 55.140 ;
        RECT 115.695 53.430 116.055 54.050 ;
        RECT 115.775 52.550 116.035 53.430 ;
        RECT 116.315 53.180 119.145 54.230 ;
        RECT 115.605 52.170 116.135 52.550 ;
        RECT 116.335 51.960 117.465 53.180 ;
        RECT 118.825 53.160 119.145 53.180 ;
        RECT 112.135 50.930 112.405 51.880 ;
        RECT 112.135 50.780 112.605 50.930 ;
        RECT 112.135 50.100 112.695 50.780 ;
        RECT 112.215 50.090 112.695 50.100 ;
        RECT 111.505 49.560 112.125 49.920 ;
        RECT 111.545 49.030 111.975 49.560 ;
        RECT 110.095 48.610 111.975 49.030 ;
        RECT 112.465 48.900 112.695 50.090 ;
        RECT 111.545 47.740 111.975 48.610 ;
        RECT 112.385 48.300 112.765 48.900 ;
        RECT 104.895 46.860 105.195 47.720 ;
        RECT 105.975 46.860 106.275 47.720 ;
        RECT 111.365 47.380 111.985 47.740 ;
        RECT 111.985 46.930 112.255 47.180 ;
        RECT 112.465 46.930 112.695 48.300 ;
        RECT 111.985 46.820 112.695 46.930 ;
        RECT 116.165 47.720 117.545 51.960 ;
        RECT 121.345 49.030 121.735 70.540 ;
        RECT 127.665 63.140 127.935 65.180 ;
        RECT 128.795 63.140 129.065 65.140 ;
        RECT 127.665 56.450 129.065 63.140 ;
        RECT 127.665 55.130 127.935 56.450 ;
        RECT 128.795 55.090 129.065 56.450 ;
        RECT 130.065 55.200 130.385 65.130 ;
        RECT 130.065 55.140 130.395 55.200 ;
        RECT 127.585 54.230 128.715 54.240 ;
        RECT 130.075 54.230 130.395 55.140 ;
        RECT 126.945 53.430 127.305 54.050 ;
        RECT 127.025 52.550 127.285 53.430 ;
        RECT 127.565 53.180 130.395 54.230 ;
        RECT 126.855 52.170 127.385 52.550 ;
        RECT 127.585 51.960 128.715 53.180 ;
        RECT 130.075 53.160 130.395 53.180 ;
        RECT 123.385 50.930 123.655 51.880 ;
        RECT 123.385 50.780 123.855 50.930 ;
        RECT 123.385 50.100 123.945 50.780 ;
        RECT 123.465 50.090 123.945 50.100 ;
        RECT 122.755 49.560 123.375 49.920 ;
        RECT 122.795 49.030 123.225 49.560 ;
        RECT 121.345 48.610 123.225 49.030 ;
        RECT 123.715 48.900 123.945 50.090 ;
        RECT 122.795 47.740 123.225 48.610 ;
        RECT 123.635 48.300 124.015 48.900 ;
        RECT 116.165 46.860 116.465 47.720 ;
        RECT 117.245 46.860 117.545 47.720 ;
        RECT 122.615 47.380 123.235 47.740 ;
        RECT 123.235 46.930 123.505 47.180 ;
        RECT 123.715 46.930 123.945 48.300 ;
        RECT 123.235 46.820 123.945 46.930 ;
        RECT 127.415 47.720 128.795 51.960 ;
        RECT 127.415 46.860 127.715 47.720 ;
        RECT 128.495 46.860 128.795 47.720 ;
        RECT 89.435 46.350 89.705 46.520 ;
        RECT 94.945 46.330 95.425 46.710 ;
        RECT 100.715 46.510 101.375 46.820 ;
        RECT 100.715 46.340 100.985 46.510 ;
        RECT 72.455 45.110 72.835 45.710 ;
        RECT 83.795 45.700 84.045 46.320 ;
        RECT 95.045 45.710 95.295 46.330 ;
        RECT 106.225 46.320 106.705 46.700 ;
        RECT 111.985 46.510 112.645 46.820 ;
        RECT 111.985 46.340 112.255 46.510 ;
        RECT 117.495 46.320 117.975 46.700 ;
        RECT 123.235 46.510 123.895 46.820 ;
        RECT 123.235 46.340 123.505 46.510 ;
        RECT 128.745 46.320 129.225 46.700 ;
        RECT 83.695 45.100 84.075 45.700 ;
        RECT 94.945 45.110 95.325 45.710 ;
        RECT 106.325 45.700 106.575 46.320 ;
        RECT 117.595 45.700 117.845 46.320 ;
        RECT 128.845 45.700 129.095 46.320 ;
        RECT 106.225 45.100 106.605 45.700 ;
        RECT 117.495 45.100 117.875 45.700 ;
        RECT 128.745 45.100 129.125 45.700 ;
        RECT 20.795 39.650 21.175 40.250 ;
        RECT 32.075 39.650 32.455 40.250 ;
        RECT 20.825 39.030 21.075 39.650 ;
        RECT 32.105 39.030 32.355 39.650 ;
        RECT 43.365 39.630 43.745 40.230 ;
        RECT 54.585 39.630 54.965 40.230 ;
        RECT 65.785 39.630 66.165 40.230 ;
        RECT 20.695 38.650 21.175 39.030 ;
        RECT 26.415 38.840 26.685 39.010 ;
        RECT 26.025 38.530 26.685 38.840 ;
        RECT 31.975 38.650 32.455 39.030 ;
        RECT 43.395 39.010 43.645 39.630 ;
        RECT 54.615 39.010 54.865 39.630 ;
        RECT 65.815 39.010 66.065 39.630 ;
        RECT 77.075 39.620 77.455 40.220 ;
        RECT 88.315 39.640 88.695 40.240 ;
        RECT 99.525 39.660 99.905 40.260 ;
        RECT 110.725 39.700 111.105 40.300 ;
        RECT 121.935 39.720 122.315 40.320 ;
        RECT 37.695 38.840 37.965 39.010 ;
        RECT 37.305 38.530 37.965 38.840 ;
        RECT 43.265 38.630 43.745 39.010 ;
        RECT 48.985 38.820 49.255 38.990 ;
        RECT 21.125 37.630 21.425 38.490 ;
        RECT 22.205 37.630 22.505 38.490 ;
        RECT 21.125 33.390 22.505 37.630 ;
        RECT 25.975 38.420 26.685 38.530 ;
        RECT 25.975 37.050 26.205 38.420 ;
        RECT 26.415 38.170 26.685 38.420 ;
        RECT 26.685 37.610 27.305 37.970 ;
        RECT 32.405 37.630 32.705 38.490 ;
        RECT 33.485 37.630 33.785 38.490 ;
        RECT 25.905 36.450 26.285 37.050 ;
        RECT 26.695 36.740 27.125 37.610 ;
        RECT 25.975 35.260 26.205 36.450 ;
        RECT 26.695 36.320 28.575 36.740 ;
        RECT 26.695 35.790 27.125 36.320 ;
        RECT 26.545 35.430 27.165 35.790 ;
        RECT 25.975 35.250 26.455 35.260 ;
        RECT 25.975 34.570 26.535 35.250 ;
        RECT 26.065 34.420 26.535 34.570 ;
        RECT 26.265 33.470 26.535 34.420 ;
        RECT 19.525 32.170 19.845 32.190 ;
        RECT 21.205 32.170 22.335 33.390 ;
        RECT 22.535 32.800 23.065 33.180 ;
        RECT 19.525 31.120 22.355 32.170 ;
        RECT 22.635 31.920 22.895 32.800 ;
        RECT 22.615 31.300 22.975 31.920 ;
        RECT 19.525 30.210 19.845 31.120 ;
        RECT 21.205 31.110 22.335 31.120 ;
        RECT 19.525 30.150 19.855 30.210 ;
        RECT 19.535 20.220 19.855 30.150 ;
        RECT 20.855 28.900 21.125 30.260 ;
        RECT 21.985 28.900 22.255 30.220 ;
        RECT 20.855 22.210 22.255 28.900 ;
        RECT 20.855 20.210 21.125 22.210 ;
        RECT 21.985 20.170 22.255 22.210 ;
        RECT 28.185 14.810 28.575 36.320 ;
        RECT 32.405 33.390 33.785 37.630 ;
        RECT 37.255 38.420 37.965 38.530 ;
        RECT 48.595 38.510 49.255 38.820 ;
        RECT 54.485 38.630 54.965 39.010 ;
        RECT 60.205 38.820 60.475 38.990 ;
        RECT 59.815 38.510 60.475 38.820 ;
        RECT 65.685 38.630 66.165 39.010 ;
        RECT 77.105 39.000 77.355 39.620 ;
        RECT 88.345 39.020 88.595 39.640 ;
        RECT 99.555 39.040 99.805 39.660 ;
        RECT 110.755 39.080 111.005 39.700 ;
        RECT 121.965 39.100 122.215 39.720 ;
        RECT 71.405 38.820 71.675 38.990 ;
        RECT 71.015 38.510 71.675 38.820 ;
        RECT 76.975 38.620 77.455 39.000 ;
        RECT 82.695 38.810 82.965 38.980 ;
        RECT 37.255 37.050 37.485 38.420 ;
        RECT 37.695 38.170 37.965 38.420 ;
        RECT 37.965 37.610 38.585 37.970 ;
        RECT 43.695 37.610 43.995 38.470 ;
        RECT 44.775 37.610 45.075 38.470 ;
        RECT 37.185 36.450 37.565 37.050 ;
        RECT 37.975 36.740 38.405 37.610 ;
        RECT 37.255 35.260 37.485 36.450 ;
        RECT 37.975 36.320 39.855 36.740 ;
        RECT 37.975 35.790 38.405 36.320 ;
        RECT 37.825 35.430 38.445 35.790 ;
        RECT 37.255 35.250 37.735 35.260 ;
        RECT 37.255 34.570 37.815 35.250 ;
        RECT 37.345 34.420 37.815 34.570 ;
        RECT 37.545 33.470 37.815 34.420 ;
        RECT 30.805 32.170 31.125 32.190 ;
        RECT 32.485 32.170 33.615 33.390 ;
        RECT 33.815 32.800 34.345 33.180 ;
        RECT 30.805 31.120 33.635 32.170 ;
        RECT 33.915 31.920 34.175 32.800 ;
        RECT 33.895 31.300 34.255 31.920 ;
        RECT 30.805 30.210 31.125 31.120 ;
        RECT 32.485 31.110 33.615 31.120 ;
        RECT 30.805 30.150 31.135 30.210 ;
        RECT 30.815 20.220 31.135 30.150 ;
        RECT 32.135 28.900 32.405 30.260 ;
        RECT 33.265 28.900 33.535 30.220 ;
        RECT 32.135 22.210 33.535 28.900 ;
        RECT 32.135 20.210 32.405 22.210 ;
        RECT 33.265 20.170 33.535 22.210 ;
        RECT 39.465 14.810 39.855 36.320 ;
        RECT 43.695 33.370 45.075 37.610 ;
        RECT 48.545 38.400 49.255 38.510 ;
        RECT 48.545 37.030 48.775 38.400 ;
        RECT 48.985 38.150 49.255 38.400 ;
        RECT 49.255 37.590 49.875 37.950 ;
        RECT 54.915 37.610 55.215 38.470 ;
        RECT 55.995 37.610 56.295 38.470 ;
        RECT 48.475 36.430 48.855 37.030 ;
        RECT 49.265 36.720 49.695 37.590 ;
        RECT 48.545 35.240 48.775 36.430 ;
        RECT 49.265 36.300 51.145 36.720 ;
        RECT 49.265 35.770 49.695 36.300 ;
        RECT 49.115 35.410 49.735 35.770 ;
        RECT 48.545 35.230 49.025 35.240 ;
        RECT 48.545 34.550 49.105 35.230 ;
        RECT 48.635 34.400 49.105 34.550 ;
        RECT 48.835 33.450 49.105 34.400 ;
        RECT 42.095 32.150 42.415 32.170 ;
        RECT 43.775 32.150 44.905 33.370 ;
        RECT 45.105 32.780 45.635 33.160 ;
        RECT 42.095 31.100 44.925 32.150 ;
        RECT 45.205 31.900 45.465 32.780 ;
        RECT 45.185 31.280 45.545 31.900 ;
        RECT 42.095 30.190 42.415 31.100 ;
        RECT 43.775 31.090 44.905 31.100 ;
        RECT 42.095 30.130 42.425 30.190 ;
        RECT 42.105 20.200 42.425 30.130 ;
        RECT 43.425 28.880 43.695 30.240 ;
        RECT 44.555 28.880 44.825 30.200 ;
        RECT 43.425 22.190 44.825 28.880 ;
        RECT 43.425 20.190 43.695 22.190 ;
        RECT 44.555 20.150 44.825 22.190 ;
        RECT 28.185 12.290 28.595 14.810 ;
        RECT 28.185 11.950 30.415 12.290 ;
        RECT 39.465 11.990 39.875 14.810 ;
        RECT 50.755 14.790 51.145 36.300 ;
        RECT 54.915 33.370 56.295 37.610 ;
        RECT 59.765 38.400 60.475 38.510 ;
        RECT 59.765 37.030 59.995 38.400 ;
        RECT 60.205 38.150 60.475 38.400 ;
        RECT 60.475 37.590 61.095 37.950 ;
        RECT 66.115 37.610 66.415 38.470 ;
        RECT 67.195 37.610 67.495 38.470 ;
        RECT 59.695 36.430 60.075 37.030 ;
        RECT 60.485 36.720 60.915 37.590 ;
        RECT 59.765 35.240 59.995 36.430 ;
        RECT 60.485 36.300 62.365 36.720 ;
        RECT 60.485 35.770 60.915 36.300 ;
        RECT 60.335 35.410 60.955 35.770 ;
        RECT 59.765 35.230 60.245 35.240 ;
        RECT 59.765 34.550 60.325 35.230 ;
        RECT 59.855 34.400 60.325 34.550 ;
        RECT 60.055 33.450 60.325 34.400 ;
        RECT 53.315 32.150 53.635 32.170 ;
        RECT 54.995 32.150 56.125 33.370 ;
        RECT 56.325 32.780 56.855 33.160 ;
        RECT 53.315 31.100 56.145 32.150 ;
        RECT 56.425 31.900 56.685 32.780 ;
        RECT 56.405 31.280 56.765 31.900 ;
        RECT 53.315 30.190 53.635 31.100 ;
        RECT 54.995 31.090 56.125 31.100 ;
        RECT 53.315 30.130 53.645 30.190 ;
        RECT 53.325 20.200 53.645 30.130 ;
        RECT 54.645 28.880 54.915 30.240 ;
        RECT 55.775 28.880 56.045 30.200 ;
        RECT 54.645 22.190 56.045 28.880 ;
        RECT 54.645 20.190 54.915 22.190 ;
        RECT 55.775 20.150 56.045 22.190 ;
        RECT 61.975 14.790 62.365 36.300 ;
        RECT 66.115 33.370 67.495 37.610 ;
        RECT 70.965 38.400 71.675 38.510 ;
        RECT 82.305 38.500 82.965 38.810 ;
        RECT 88.215 38.640 88.695 39.020 ;
        RECT 93.935 38.830 94.205 39.000 ;
        RECT 93.545 38.520 94.205 38.830 ;
        RECT 99.425 38.660 99.905 39.040 ;
        RECT 105.145 38.850 105.415 39.020 ;
        RECT 104.755 38.540 105.415 38.850 ;
        RECT 110.625 38.700 111.105 39.080 ;
        RECT 116.345 38.890 116.615 39.060 ;
        RECT 115.955 38.580 116.615 38.890 ;
        RECT 121.835 38.720 122.315 39.100 ;
        RECT 127.555 38.910 127.825 39.080 ;
        RECT 127.165 38.600 127.825 38.910 ;
        RECT 70.965 37.030 71.195 38.400 ;
        RECT 71.405 38.150 71.675 38.400 ;
        RECT 71.675 37.590 72.295 37.950 ;
        RECT 77.405 37.600 77.705 38.460 ;
        RECT 78.485 37.600 78.785 38.460 ;
        RECT 70.895 36.430 71.275 37.030 ;
        RECT 71.685 36.720 72.115 37.590 ;
        RECT 70.965 35.240 71.195 36.430 ;
        RECT 71.685 36.300 73.565 36.720 ;
        RECT 71.685 35.770 72.115 36.300 ;
        RECT 71.535 35.410 72.155 35.770 ;
        RECT 70.965 35.230 71.445 35.240 ;
        RECT 70.965 34.550 71.525 35.230 ;
        RECT 71.055 34.400 71.525 34.550 ;
        RECT 71.255 33.450 71.525 34.400 ;
        RECT 64.515 32.150 64.835 32.170 ;
        RECT 66.195 32.150 67.325 33.370 ;
        RECT 67.525 32.780 68.055 33.160 ;
        RECT 64.515 31.100 67.345 32.150 ;
        RECT 67.625 31.900 67.885 32.780 ;
        RECT 67.605 31.280 67.965 31.900 ;
        RECT 64.515 30.190 64.835 31.100 ;
        RECT 66.195 31.090 67.325 31.100 ;
        RECT 64.515 30.130 64.845 30.190 ;
        RECT 64.525 20.200 64.845 30.130 ;
        RECT 65.845 28.880 66.115 30.240 ;
        RECT 66.975 28.880 67.245 30.200 ;
        RECT 65.845 22.190 67.245 28.880 ;
        RECT 65.845 20.190 66.115 22.190 ;
        RECT 66.975 20.150 67.245 22.190 ;
        RECT 73.175 14.790 73.565 36.300 ;
        RECT 77.405 33.360 78.785 37.600 ;
        RECT 82.255 38.390 82.965 38.500 ;
        RECT 82.255 37.020 82.485 38.390 ;
        RECT 82.695 38.140 82.965 38.390 ;
        RECT 82.965 37.580 83.585 37.940 ;
        RECT 88.645 37.620 88.945 38.480 ;
        RECT 89.725 37.620 90.025 38.480 ;
        RECT 82.185 36.420 82.565 37.020 ;
        RECT 82.975 36.710 83.405 37.580 ;
        RECT 82.255 35.230 82.485 36.420 ;
        RECT 82.975 36.290 84.855 36.710 ;
        RECT 82.975 35.760 83.405 36.290 ;
        RECT 82.825 35.400 83.445 35.760 ;
        RECT 82.255 35.220 82.735 35.230 ;
        RECT 82.255 34.540 82.815 35.220 ;
        RECT 82.345 34.390 82.815 34.540 ;
        RECT 82.545 33.440 82.815 34.390 ;
        RECT 75.805 32.140 76.125 32.160 ;
        RECT 77.485 32.140 78.615 33.360 ;
        RECT 78.815 32.770 79.345 33.150 ;
        RECT 75.805 31.090 78.635 32.140 ;
        RECT 78.915 31.890 79.175 32.770 ;
        RECT 78.895 31.270 79.255 31.890 ;
        RECT 75.805 30.180 76.125 31.090 ;
        RECT 77.485 31.080 78.615 31.090 ;
        RECT 75.805 30.120 76.135 30.180 ;
        RECT 75.815 20.190 76.135 30.120 ;
        RECT 77.135 28.870 77.405 30.230 ;
        RECT 78.265 28.870 78.535 30.190 ;
        RECT 77.135 22.180 78.535 28.870 ;
        RECT 77.135 20.180 77.405 22.180 ;
        RECT 78.265 20.140 78.535 22.180 ;
        RECT 50.755 12.170 51.165 14.790 ;
        RECT 27.865 11.130 30.415 11.950 ;
        RECT 28.395 11.090 30.415 11.130 ;
        RECT 39.115 10.980 41.565 11.990 ;
        RECT 50.335 10.970 52.355 12.170 ;
        RECT 61.975 12.160 62.385 14.790 ;
        RECT 73.175 12.190 73.585 14.790 ;
        RECT 84.465 14.780 84.855 36.290 ;
        RECT 88.645 33.380 90.025 37.620 ;
        RECT 93.495 38.410 94.205 38.520 ;
        RECT 93.495 37.040 93.725 38.410 ;
        RECT 93.935 38.160 94.205 38.410 ;
        RECT 94.205 37.600 94.825 37.960 ;
        RECT 99.855 37.640 100.155 38.500 ;
        RECT 100.935 37.640 101.235 38.500 ;
        RECT 93.425 36.440 93.805 37.040 ;
        RECT 94.215 36.730 94.645 37.600 ;
        RECT 93.495 35.250 93.725 36.440 ;
        RECT 94.215 36.310 96.095 36.730 ;
        RECT 94.215 35.780 94.645 36.310 ;
        RECT 94.065 35.420 94.685 35.780 ;
        RECT 93.495 35.240 93.975 35.250 ;
        RECT 93.495 34.560 94.055 35.240 ;
        RECT 93.585 34.410 94.055 34.560 ;
        RECT 93.785 33.460 94.055 34.410 ;
        RECT 87.045 32.160 87.365 32.180 ;
        RECT 88.725 32.160 89.855 33.380 ;
        RECT 90.055 32.790 90.585 33.170 ;
        RECT 87.045 31.110 89.875 32.160 ;
        RECT 90.155 31.910 90.415 32.790 ;
        RECT 90.135 31.290 90.495 31.910 ;
        RECT 87.045 30.200 87.365 31.110 ;
        RECT 88.725 31.100 89.855 31.110 ;
        RECT 87.045 30.140 87.375 30.200 ;
        RECT 87.055 20.210 87.375 30.140 ;
        RECT 88.375 28.890 88.645 30.250 ;
        RECT 89.505 28.890 89.775 30.210 ;
        RECT 88.375 22.200 89.775 28.890 ;
        RECT 88.375 20.200 88.645 22.200 ;
        RECT 89.505 20.160 89.775 22.200 ;
        RECT 95.705 14.800 96.095 36.310 ;
        RECT 99.855 33.400 101.235 37.640 ;
        RECT 104.705 38.430 105.415 38.540 ;
        RECT 104.705 37.060 104.935 38.430 ;
        RECT 105.145 38.180 105.415 38.430 ;
        RECT 105.415 37.620 106.035 37.980 ;
        RECT 111.055 37.680 111.355 38.540 ;
        RECT 112.135 37.680 112.435 38.540 ;
        RECT 104.635 36.460 105.015 37.060 ;
        RECT 105.425 36.750 105.855 37.620 ;
        RECT 104.705 35.270 104.935 36.460 ;
        RECT 105.425 36.330 107.305 36.750 ;
        RECT 105.425 35.800 105.855 36.330 ;
        RECT 105.275 35.440 105.895 35.800 ;
        RECT 104.705 35.260 105.185 35.270 ;
        RECT 104.705 34.580 105.265 35.260 ;
        RECT 104.795 34.430 105.265 34.580 ;
        RECT 104.995 33.480 105.265 34.430 ;
        RECT 98.255 32.180 98.575 32.200 ;
        RECT 99.935 32.180 101.065 33.400 ;
        RECT 101.265 32.810 101.795 33.190 ;
        RECT 98.255 31.130 101.085 32.180 ;
        RECT 101.365 31.930 101.625 32.810 ;
        RECT 101.345 31.310 101.705 31.930 ;
        RECT 98.255 30.220 98.575 31.130 ;
        RECT 99.935 31.120 101.065 31.130 ;
        RECT 98.255 30.160 98.585 30.220 ;
        RECT 98.265 20.230 98.585 30.160 ;
        RECT 99.585 28.910 99.855 30.270 ;
        RECT 100.715 28.910 100.985 30.230 ;
        RECT 99.585 22.220 100.985 28.910 ;
        RECT 99.585 20.220 99.855 22.220 ;
        RECT 100.715 20.180 100.985 22.220 ;
        RECT 106.915 14.820 107.305 36.330 ;
        RECT 111.055 33.440 112.435 37.680 ;
        RECT 115.905 38.470 116.615 38.580 ;
        RECT 115.905 37.100 116.135 38.470 ;
        RECT 116.345 38.220 116.615 38.470 ;
        RECT 116.615 37.660 117.235 38.020 ;
        RECT 122.265 37.700 122.565 38.560 ;
        RECT 123.345 37.700 123.645 38.560 ;
        RECT 115.835 36.500 116.215 37.100 ;
        RECT 116.625 36.790 117.055 37.660 ;
        RECT 115.905 35.310 116.135 36.500 ;
        RECT 116.625 36.370 118.505 36.790 ;
        RECT 116.625 35.840 117.055 36.370 ;
        RECT 116.475 35.480 117.095 35.840 ;
        RECT 115.905 35.300 116.385 35.310 ;
        RECT 115.905 34.620 116.465 35.300 ;
        RECT 115.995 34.470 116.465 34.620 ;
        RECT 116.195 33.520 116.465 34.470 ;
        RECT 109.455 32.220 109.775 32.240 ;
        RECT 111.135 32.220 112.265 33.440 ;
        RECT 112.465 32.850 112.995 33.230 ;
        RECT 109.455 31.170 112.285 32.220 ;
        RECT 112.565 31.970 112.825 32.850 ;
        RECT 112.545 31.350 112.905 31.970 ;
        RECT 109.455 30.260 109.775 31.170 ;
        RECT 111.135 31.160 112.265 31.170 ;
        RECT 109.455 30.200 109.785 30.260 ;
        RECT 109.465 20.270 109.785 30.200 ;
        RECT 110.785 28.950 111.055 30.310 ;
        RECT 111.915 28.950 112.185 30.270 ;
        RECT 110.785 22.260 112.185 28.950 ;
        RECT 110.785 20.260 111.055 22.260 ;
        RECT 111.915 20.220 112.185 22.260 ;
        RECT 118.115 14.860 118.505 36.370 ;
        RECT 122.265 33.460 123.645 37.700 ;
        RECT 127.115 38.490 127.825 38.600 ;
        RECT 127.115 37.120 127.345 38.490 ;
        RECT 127.555 38.240 127.825 38.490 ;
        RECT 127.825 37.680 128.445 38.040 ;
        RECT 127.045 36.520 127.425 37.120 ;
        RECT 127.835 36.810 128.265 37.680 ;
        RECT 127.115 35.330 127.345 36.520 ;
        RECT 127.835 36.390 129.715 36.810 ;
        RECT 127.835 35.860 128.265 36.390 ;
        RECT 127.685 35.500 128.305 35.860 ;
        RECT 127.115 35.320 127.595 35.330 ;
        RECT 127.115 34.640 127.675 35.320 ;
        RECT 127.205 34.490 127.675 34.640 ;
        RECT 127.405 33.540 127.675 34.490 ;
        RECT 120.665 32.240 120.985 32.260 ;
        RECT 122.345 32.240 123.475 33.460 ;
        RECT 123.675 32.870 124.205 33.250 ;
        RECT 120.665 31.190 123.495 32.240 ;
        RECT 123.775 31.990 124.035 32.870 ;
        RECT 123.755 31.370 124.115 31.990 ;
        RECT 120.665 30.280 120.985 31.190 ;
        RECT 122.345 31.180 123.475 31.190 ;
        RECT 120.665 30.220 120.995 30.280 ;
        RECT 120.675 20.290 120.995 30.220 ;
        RECT 121.995 28.970 122.265 30.330 ;
        RECT 123.125 28.970 123.395 30.290 ;
        RECT 121.995 22.280 123.395 28.970 ;
        RECT 121.995 20.280 122.265 22.280 ;
        RECT 123.125 20.240 123.395 22.280 ;
        RECT 129.325 14.880 129.715 36.390 ;
        RECT 61.415 10.960 63.435 12.160 ;
        RECT 72.725 10.990 74.745 12.190 ;
        RECT 84.465 12.180 84.875 14.780 ;
        RECT 95.705 12.180 96.115 14.800 ;
        RECT 106.915 12.230 107.325 14.820 ;
        RECT 118.115 12.230 118.525 14.860 ;
        RECT 129.325 12.260 129.735 14.880 ;
        RECT 83.845 10.980 85.865 12.180 ;
        RECT 95.145 10.980 97.165 12.180 ;
        RECT 106.335 11.030 108.355 12.230 ;
        RECT 117.565 11.030 119.585 12.230 ;
        RECT 128.865 11.060 130.885 12.260 ;
      LAYER met3 ;
        RECT 66.245 179.820 66.575 179.835 ;
        RECT 70.845 179.820 71.175 179.835 ;
        RECT 66.245 179.520 71.175 179.820 ;
        RECT 66.245 179.505 66.575 179.520 ;
        RECT 70.845 179.505 71.175 179.520 ;
        RECT 70.130 179.140 70.510 179.150 ;
        RECT 83.725 179.140 84.055 179.155 ;
        RECT 70.130 178.840 84.055 179.140 ;
        RECT 70.130 178.830 70.510 178.840 ;
        RECT 83.725 178.825 84.055 178.840 ;
        RECT 65.325 177.780 65.655 177.795 ;
        RECT 69.005 177.780 69.335 177.795 ;
        RECT 65.325 177.480 69.335 177.780 ;
        RECT 65.325 177.465 65.655 177.480 ;
        RECT 69.005 177.465 69.335 177.480 ;
        RECT 69.925 177.780 70.255 177.795 ;
        RECT 72.225 177.780 72.555 177.795 ;
        RECT 74.985 177.780 75.315 177.795 ;
        RECT 69.925 177.480 75.315 177.780 ;
        RECT 69.925 177.465 70.255 177.480 ;
        RECT 72.225 177.465 72.555 177.480 ;
        RECT 74.985 177.465 75.315 177.480 ;
        RECT 83.725 177.780 84.055 177.795 ;
        RECT 102.125 177.780 102.455 177.795 ;
        RECT 83.725 177.480 102.455 177.780 ;
        RECT 83.725 177.465 84.055 177.480 ;
        RECT 102.125 177.465 102.455 177.480 ;
        RECT 57.505 177.100 57.835 177.115 ;
        RECT 74.065 177.100 74.395 177.115 ;
        RECT 57.505 176.800 74.395 177.100 ;
        RECT 57.505 176.785 57.835 176.800 ;
        RECT 74.065 176.785 74.395 176.800 ;
        RECT 50.810 171.660 51.190 171.670 ;
        RECT 53.365 171.660 53.695 171.675 ;
        RECT 50.810 171.360 53.695 171.660 ;
        RECT 50.810 171.350 51.190 171.360 ;
        RECT 53.365 171.345 53.695 171.360 ;
        RECT 36.345 166.900 36.675 166.915 ;
        RECT 50.810 166.900 51.190 166.910 ;
        RECT 36.345 166.600 51.190 166.900 ;
        RECT 36.345 166.585 36.675 166.600 ;
        RECT 50.810 166.590 51.190 166.600 ;
        RECT 50.810 155.340 51.190 155.350 ;
        RECT 57.250 155.340 57.630 155.350 ;
        RECT 66.705 155.340 67.035 155.355 ;
        RECT 70.130 155.340 70.510 155.350 ;
        RECT 50.810 155.040 70.510 155.340 ;
        RECT 50.810 155.030 51.190 155.040 ;
        RECT 57.250 155.030 57.630 155.040 ;
        RECT 66.705 155.025 67.035 155.040 ;
        RECT 70.130 155.030 70.510 155.040 ;
        RECT 54.745 147.180 55.075 147.195 ;
        RECT 58.885 147.180 59.215 147.195 ;
        RECT 54.745 146.880 59.215 147.180 ;
        RECT 54.745 146.865 55.075 146.880 ;
        RECT 58.885 146.865 59.215 146.880 ;
        RECT 103.505 136.980 103.835 136.995 ;
        RECT 109.025 136.980 109.355 136.995 ;
        RECT 103.505 136.680 109.355 136.980 ;
        RECT 103.505 136.665 103.835 136.680 ;
        RECT 109.025 136.665 109.355 136.680 ;
        RECT 36.805 124.740 37.135 124.755 ;
        RECT 51.065 124.740 51.395 124.755 ;
        RECT 57.250 124.740 57.630 124.750 ;
        RECT 36.805 124.440 57.630 124.740 ;
        RECT 36.805 124.425 37.135 124.440 ;
        RECT 51.065 124.425 51.395 124.440 ;
        RECT 57.250 124.430 57.630 124.440 ;
        RECT 57.290 123.380 57.590 124.430 ;
        RECT 89.245 123.380 89.575 123.395 ;
        RECT 105.345 123.380 105.675 123.395 ;
        RECT 57.290 123.080 105.675 123.380 ;
        RECT 89.245 123.065 89.575 123.080 ;
        RECT 105.345 123.065 105.675 123.080 ;
        RECT 13.950 87.980 14.980 88.515 ;
        RECT 13.950 87.500 14.990 87.980 ;
        RECT 13.950 87.175 14.980 87.500 ;
        RECT 14.070 86.570 14.810 87.175 ;
        RECT 20.050 87.105 20.920 88.515 ;
        RECT 14.070 75.715 14.700 86.570 ;
        RECT 20.170 77.115 20.800 87.105 ;
        RECT 25.910 87.055 26.860 88.515 ;
        RECT 26.070 78.385 26.700 87.055 ;
        RECT 31.730 86.965 32.910 88.585 ;
        RECT 32.005 79.615 32.635 86.965 ;
        RECT 37.630 86.835 39.120 88.755 ;
        RECT 38.060 81.125 38.690 86.835 ;
        RECT 43.790 86.745 45.190 88.605 ;
        RECT 49.710 86.945 51.060 88.615 ;
        RECT 44.175 82.625 44.805 86.745 ;
        RECT 50.070 83.875 50.700 86.945 ;
        RECT 55.530 86.785 56.750 88.545 ;
        RECT 55.825 85.115 56.455 86.785 ;
        RECT 61.670 86.625 63.180 88.615 ;
        RECT 67.680 88.305 68.720 89.815 ;
        RECT 67.885 87.225 68.515 88.305 ;
        RECT 62.110 86.175 62.740 86.625 ;
        RECT 67.885 86.595 130.605 87.225 ;
        RECT 62.110 85.545 118.855 86.175 ;
        RECT 55.825 84.485 107.605 85.115 ;
        RECT 50.070 83.245 96.285 83.875 ;
        RECT 44.175 81.995 85.055 82.625 ;
        RECT 38.060 80.495 73.765 81.125 ;
        RECT 32.005 78.985 62.635 79.615 ;
        RECT 26.070 77.755 51.245 78.385 ;
        RECT 20.170 76.485 40.645 77.115 ;
        RECT 14.070 75.660 29.295 75.715 ;
        RECT 40.015 75.710 40.645 76.485 ;
        RECT 14.070 75.085 30.410 75.660 ;
        RECT 27.850 74.670 30.410 75.085 ;
        RECT 27.850 73.120 30.450 74.670 ;
        RECT 39.060 74.510 41.620 75.710 ;
        RECT 50.615 75.580 51.245 77.755 ;
        RECT 62.005 75.690 62.635 78.985 ;
        RECT 49.930 74.650 52.490 75.580 ;
        RECT 20.145 54.060 20.605 54.135 ;
        RECT 25.715 54.060 26.175 54.085 ;
        RECT 20.145 53.620 26.175 54.060 ;
        RECT 20.145 53.565 20.605 53.620 ;
        RECT 25.715 53.515 26.175 53.620 ;
        RECT 22.405 48.870 22.885 48.935 ;
        RECT 22.405 48.550 24.205 48.870 ;
        RECT 22.405 48.385 22.885 48.550 ;
        RECT 23.635 45.710 24.195 48.550 ;
        RECT 27.515 45.710 27.995 45.735 ;
        RECT 23.635 45.290 27.995 45.710 ;
        RECT 23.635 45.280 24.195 45.290 ;
        RECT 27.515 45.185 27.995 45.290 ;
        RECT 20.745 40.120 21.225 40.225 ;
        RECT 24.545 40.120 25.105 40.130 ;
        RECT 20.745 39.700 25.105 40.120 ;
        RECT 20.745 39.675 21.225 39.700 ;
        RECT 24.545 36.860 25.105 39.700 ;
        RECT 25.855 36.860 26.335 37.025 ;
        RECT 24.535 36.540 26.335 36.860 ;
        RECT 25.855 36.475 26.335 36.540 ;
        RECT 22.565 31.790 23.025 31.895 ;
        RECT 28.135 31.790 28.595 31.845 ;
        RECT 22.565 31.350 28.595 31.790 ;
        RECT 22.565 31.325 23.025 31.350 ;
        RECT 28.135 31.275 28.595 31.350 ;
        RECT 29.765 12.265 30.255 73.120 ;
        RECT 38.960 73.080 41.730 74.510 ;
        RECT 31.345 54.070 31.805 54.145 ;
        RECT 36.915 54.070 37.375 54.095 ;
        RECT 31.345 53.630 37.375 54.070 ;
        RECT 31.345 53.575 31.805 53.630 ;
        RECT 36.915 53.525 37.375 53.630 ;
        RECT 33.605 48.880 34.085 48.945 ;
        RECT 33.605 48.560 35.405 48.880 ;
        RECT 33.605 48.395 34.085 48.560 ;
        RECT 34.835 45.720 35.395 48.560 ;
        RECT 38.715 45.720 39.195 45.745 ;
        RECT 34.835 45.300 39.195 45.720 ;
        RECT 34.835 45.290 35.395 45.300 ;
        RECT 38.715 45.195 39.195 45.300 ;
        RECT 32.025 40.120 32.505 40.225 ;
        RECT 35.825 40.120 36.385 40.130 ;
        RECT 32.025 39.700 36.385 40.120 ;
        RECT 32.025 39.675 32.505 39.700 ;
        RECT 35.825 36.860 36.385 39.700 ;
        RECT 37.135 36.860 37.615 37.025 ;
        RECT 35.815 36.540 37.615 36.860 ;
        RECT 37.135 36.475 37.615 36.540 ;
        RECT 33.845 31.790 34.305 31.895 ;
        RECT 39.415 31.790 39.875 31.845 ;
        RECT 33.845 31.350 39.875 31.790 ;
        RECT 33.845 31.325 34.305 31.350 ;
        RECT 39.415 31.275 39.875 31.350 ;
        RECT 41.055 12.360 41.545 73.080 ;
        RECT 49.930 73.030 52.530 74.650 ;
        RECT 61.330 74.530 63.890 75.690 ;
        RECT 73.135 75.580 73.765 80.495 ;
        RECT 84.425 75.690 85.055 81.995 ;
        RECT 72.340 74.980 74.900 75.580 ;
        RECT 42.565 54.040 43.025 54.115 ;
        RECT 48.135 54.040 48.595 54.065 ;
        RECT 42.565 53.600 48.595 54.040 ;
        RECT 42.565 53.545 43.025 53.600 ;
        RECT 48.135 53.495 48.595 53.600 ;
        RECT 44.825 48.850 45.305 48.915 ;
        RECT 44.825 48.530 46.625 48.850 ;
        RECT 44.825 48.365 45.305 48.530 ;
        RECT 46.055 45.690 46.615 48.530 ;
        RECT 49.935 45.690 50.415 45.715 ;
        RECT 46.055 45.270 50.415 45.690 ;
        RECT 46.055 45.260 46.615 45.270 ;
        RECT 49.935 45.165 50.415 45.270 ;
        RECT 43.315 40.100 43.795 40.205 ;
        RECT 47.115 40.100 47.675 40.110 ;
        RECT 43.315 39.680 47.675 40.100 ;
        RECT 43.315 39.655 43.795 39.680 ;
        RECT 47.115 36.840 47.675 39.680 ;
        RECT 48.425 36.840 48.905 37.005 ;
        RECT 47.105 36.520 48.905 36.840 ;
        RECT 48.425 36.455 48.905 36.520 ;
        RECT 45.135 31.770 45.595 31.875 ;
        RECT 50.705 31.770 51.165 31.825 ;
        RECT 45.135 31.330 51.165 31.770 ;
        RECT 45.135 31.305 45.595 31.330 ;
        RECT 50.705 31.255 51.165 31.330 ;
        RECT 41.055 12.350 41.555 12.360 ;
        RECT 28.345 11.115 30.465 12.265 ;
        RECT 41.065 11.965 41.555 12.350 ;
        RECT 51.635 12.145 52.125 73.030 ;
        RECT 61.260 73.010 64.060 74.530 ;
        RECT 72.340 73.050 75.020 74.980 ;
        RECT 83.730 74.540 86.290 75.690 ;
        RECT 95.655 75.580 96.285 83.245 ;
        RECT 106.975 75.640 107.605 84.485 ;
        RECT 118.225 75.650 118.855 85.545 ;
        RECT 129.975 75.650 130.605 86.595 ;
        RECT 53.815 54.020 54.275 54.095 ;
        RECT 59.385 54.020 59.845 54.045 ;
        RECT 53.815 53.580 59.845 54.020 ;
        RECT 53.815 53.525 54.275 53.580 ;
        RECT 59.385 53.475 59.845 53.580 ;
        RECT 56.075 48.830 56.555 48.895 ;
        RECT 56.075 48.510 57.875 48.830 ;
        RECT 56.075 48.345 56.555 48.510 ;
        RECT 57.305 45.670 57.865 48.510 ;
        RECT 61.185 45.670 61.665 45.695 ;
        RECT 57.305 45.250 61.665 45.670 ;
        RECT 57.305 45.240 57.865 45.250 ;
        RECT 61.185 45.145 61.665 45.250 ;
        RECT 54.535 40.100 55.015 40.205 ;
        RECT 58.335 40.100 58.895 40.110 ;
        RECT 54.535 39.680 58.895 40.100 ;
        RECT 54.535 39.655 55.015 39.680 ;
        RECT 58.335 36.840 58.895 39.680 ;
        RECT 59.645 36.840 60.125 37.005 ;
        RECT 58.325 36.520 60.125 36.840 ;
        RECT 59.645 36.455 60.125 36.520 ;
        RECT 56.355 31.770 56.815 31.875 ;
        RECT 61.925 31.770 62.385 31.825 ;
        RECT 56.355 31.330 62.385 31.770 ;
        RECT 56.355 31.305 56.815 31.330 ;
        RECT 61.925 31.255 62.385 31.330 ;
        RECT 29.765 11.100 30.255 11.115 ;
        RECT 39.065 11.005 41.615 11.965 ;
        RECT 50.285 10.995 52.405 12.145 ;
        RECT 62.915 12.135 63.405 73.010 ;
        RECT 65.035 54.010 65.495 54.085 ;
        RECT 70.605 54.010 71.065 54.035 ;
        RECT 65.035 53.570 71.065 54.010 ;
        RECT 65.035 53.515 65.495 53.570 ;
        RECT 70.605 53.465 71.065 53.570 ;
        RECT 67.295 48.820 67.775 48.885 ;
        RECT 67.295 48.500 69.095 48.820 ;
        RECT 67.295 48.335 67.775 48.500 ;
        RECT 68.525 45.660 69.085 48.500 ;
        RECT 72.405 45.660 72.885 45.685 ;
        RECT 68.525 45.240 72.885 45.660 ;
        RECT 68.525 45.230 69.085 45.240 ;
        RECT 72.405 45.135 72.885 45.240 ;
        RECT 65.735 40.100 66.215 40.205 ;
        RECT 69.535 40.100 70.095 40.110 ;
        RECT 65.735 39.680 70.095 40.100 ;
        RECT 65.735 39.655 66.215 39.680 ;
        RECT 69.535 36.840 70.095 39.680 ;
        RECT 70.845 36.840 71.325 37.005 ;
        RECT 69.525 36.520 71.325 36.840 ;
        RECT 70.845 36.455 71.325 36.520 ;
        RECT 67.555 31.770 68.015 31.875 ;
        RECT 73.125 31.770 73.585 31.825 ;
        RECT 67.555 31.330 73.585 31.770 ;
        RECT 67.555 31.305 68.015 31.330 ;
        RECT 73.125 31.255 73.585 31.330 ;
        RECT 74.055 12.165 74.545 73.050 ;
        RECT 83.690 73.000 86.290 74.540 ;
        RECT 94.960 74.710 97.520 75.580 ;
        RECT 94.960 73.020 97.570 74.710 ;
        RECT 106.340 74.460 108.900 75.640 ;
        RECT 117.470 74.720 120.030 75.650 ;
        RECT 76.275 54.000 76.735 54.075 ;
        RECT 81.845 54.000 82.305 54.025 ;
        RECT 76.275 53.560 82.305 54.000 ;
        RECT 76.275 53.505 76.735 53.560 ;
        RECT 81.845 53.455 82.305 53.560 ;
        RECT 78.535 48.810 79.015 48.875 ;
        RECT 78.535 48.490 80.335 48.810 ;
        RECT 78.535 48.325 79.015 48.490 ;
        RECT 79.765 45.650 80.325 48.490 ;
        RECT 83.645 45.650 84.125 45.675 ;
        RECT 79.765 45.230 84.125 45.650 ;
        RECT 79.765 45.220 80.325 45.230 ;
        RECT 83.645 45.125 84.125 45.230 ;
        RECT 77.025 40.090 77.505 40.195 ;
        RECT 80.825 40.090 81.385 40.100 ;
        RECT 77.025 39.670 81.385 40.090 ;
        RECT 77.025 39.645 77.505 39.670 ;
        RECT 80.825 36.830 81.385 39.670 ;
        RECT 82.135 36.830 82.615 36.995 ;
        RECT 80.815 36.510 82.615 36.830 ;
        RECT 82.135 36.445 82.615 36.510 ;
        RECT 78.845 31.760 79.305 31.865 ;
        RECT 84.415 31.760 84.875 31.815 ;
        RECT 78.845 31.320 84.875 31.760 ;
        RECT 78.845 31.295 79.305 31.320 ;
        RECT 84.415 31.245 84.875 31.320 ;
        RECT 61.365 10.985 63.485 12.135 ;
        RECT 72.675 11.015 74.795 12.165 ;
        RECT 85.375 12.155 85.865 73.000 ;
        RECT 87.525 54.010 87.985 54.085 ;
        RECT 93.095 54.010 93.555 54.035 ;
        RECT 87.525 53.570 93.555 54.010 ;
        RECT 87.525 53.515 87.985 53.570 ;
        RECT 93.095 53.465 93.555 53.570 ;
        RECT 89.785 48.820 90.265 48.885 ;
        RECT 89.785 48.500 91.585 48.820 ;
        RECT 89.785 48.335 90.265 48.500 ;
        RECT 91.015 45.660 91.575 48.500 ;
        RECT 94.895 45.660 95.375 45.685 ;
        RECT 91.015 45.240 95.375 45.660 ;
        RECT 91.015 45.230 91.575 45.240 ;
        RECT 94.895 45.135 95.375 45.240 ;
        RECT 88.265 40.110 88.745 40.215 ;
        RECT 92.065 40.110 92.625 40.120 ;
        RECT 88.265 39.690 92.625 40.110 ;
        RECT 88.265 39.665 88.745 39.690 ;
        RECT 92.065 36.850 92.625 39.690 ;
        RECT 93.375 36.850 93.855 37.015 ;
        RECT 92.055 36.530 93.855 36.850 ;
        RECT 93.375 36.465 93.855 36.530 ;
        RECT 90.085 31.780 90.545 31.885 ;
        RECT 95.655 31.780 96.115 31.835 ;
        RECT 90.085 31.340 96.115 31.780 ;
        RECT 90.085 31.315 90.545 31.340 ;
        RECT 95.655 31.265 96.115 31.340 ;
        RECT 96.605 12.155 97.095 73.020 ;
        RECT 106.150 73.000 109.060 74.460 ;
        RECT 117.470 73.070 120.000 74.720 ;
        RECT 129.290 74.650 131.850 75.650 ;
        RECT 129.300 73.140 131.820 74.650 ;
        RECT 98.805 54.000 99.265 54.075 ;
        RECT 104.375 54.000 104.835 54.025 ;
        RECT 98.805 53.560 104.835 54.000 ;
        RECT 98.805 53.505 99.265 53.560 ;
        RECT 104.375 53.455 104.835 53.560 ;
        RECT 101.065 48.810 101.545 48.875 ;
        RECT 101.065 48.490 102.865 48.810 ;
        RECT 101.065 48.325 101.545 48.490 ;
        RECT 102.295 45.650 102.855 48.490 ;
        RECT 106.175 45.650 106.655 45.675 ;
        RECT 102.295 45.230 106.655 45.650 ;
        RECT 102.295 45.220 102.855 45.230 ;
        RECT 106.175 45.125 106.655 45.230 ;
        RECT 99.475 40.130 99.955 40.235 ;
        RECT 103.275 40.130 103.835 40.140 ;
        RECT 99.475 39.710 103.835 40.130 ;
        RECT 99.475 39.685 99.955 39.710 ;
        RECT 103.275 36.870 103.835 39.710 ;
        RECT 104.585 36.870 105.065 37.035 ;
        RECT 103.265 36.550 105.065 36.870 ;
        RECT 104.585 36.485 105.065 36.550 ;
        RECT 101.295 31.800 101.755 31.905 ;
        RECT 106.865 31.800 107.325 31.855 ;
        RECT 101.295 31.360 107.325 31.800 ;
        RECT 101.295 31.335 101.755 31.360 ;
        RECT 106.865 31.285 107.325 31.360 ;
        RECT 107.865 12.205 108.355 73.000 ;
        RECT 110.075 54.000 110.535 54.075 ;
        RECT 115.645 54.000 116.105 54.025 ;
        RECT 110.075 53.560 116.105 54.000 ;
        RECT 110.075 53.505 110.535 53.560 ;
        RECT 115.645 53.455 116.105 53.560 ;
        RECT 112.335 48.810 112.815 48.875 ;
        RECT 112.335 48.490 114.135 48.810 ;
        RECT 112.335 48.325 112.815 48.490 ;
        RECT 113.565 45.650 114.125 48.490 ;
        RECT 117.445 45.650 117.925 45.675 ;
        RECT 113.565 45.230 117.925 45.650 ;
        RECT 113.565 45.220 114.125 45.230 ;
        RECT 117.445 45.125 117.925 45.230 ;
        RECT 110.675 40.170 111.155 40.275 ;
        RECT 114.475 40.170 115.035 40.180 ;
        RECT 110.675 39.750 115.035 40.170 ;
        RECT 110.675 39.725 111.155 39.750 ;
        RECT 114.475 36.910 115.035 39.750 ;
        RECT 115.785 36.910 116.265 37.075 ;
        RECT 114.465 36.590 116.265 36.910 ;
        RECT 115.785 36.525 116.265 36.590 ;
        RECT 112.495 31.840 112.955 31.945 ;
        RECT 118.065 31.840 118.525 31.895 ;
        RECT 112.495 31.400 118.525 31.840 ;
        RECT 112.495 31.375 112.955 31.400 ;
        RECT 118.065 31.325 118.525 31.400 ;
        RECT 119.085 12.205 119.575 73.070 ;
        RECT 121.325 54.000 121.785 54.075 ;
        RECT 126.895 54.000 127.355 54.025 ;
        RECT 121.325 53.560 127.355 54.000 ;
        RECT 121.325 53.505 121.785 53.560 ;
        RECT 126.895 53.455 127.355 53.560 ;
        RECT 123.585 48.810 124.065 48.875 ;
        RECT 123.585 48.490 125.385 48.810 ;
        RECT 123.585 48.325 124.065 48.490 ;
        RECT 124.815 45.650 125.375 48.490 ;
        RECT 128.695 45.650 129.175 45.675 ;
        RECT 124.815 45.230 129.175 45.650 ;
        RECT 124.815 45.220 125.375 45.230 ;
        RECT 128.695 45.125 129.175 45.230 ;
        RECT 121.885 40.190 122.365 40.295 ;
        RECT 125.685 40.190 126.245 40.200 ;
        RECT 121.885 39.770 126.245 40.190 ;
        RECT 121.885 39.745 122.365 39.770 ;
        RECT 125.685 36.930 126.245 39.770 ;
        RECT 126.995 36.930 127.475 37.095 ;
        RECT 125.675 36.610 127.475 36.930 ;
        RECT 126.995 36.545 127.475 36.610 ;
        RECT 123.705 31.860 124.165 31.965 ;
        RECT 129.275 31.860 129.735 31.915 ;
        RECT 123.705 31.420 129.735 31.860 ;
        RECT 123.705 31.395 124.165 31.420 ;
        RECT 129.275 31.345 129.735 31.420 ;
        RECT 130.335 12.235 130.825 73.140 ;
        RECT 74.055 11.010 74.545 11.015 ;
        RECT 83.795 11.005 85.915 12.155 ;
        RECT 95.095 11.005 97.215 12.155 ;
        RECT 106.285 11.055 108.405 12.205 ;
        RECT 117.515 11.055 119.635 12.205 ;
        RECT 128.815 11.085 130.935 12.235 ;
        RECT 107.865 11.010 108.355 11.055 ;
        RECT 119.085 11.050 119.575 11.055 ;
        RECT 85.375 11.000 85.865 11.005 ;
        RECT 96.605 10.980 97.095 11.005 ;
      LAYER met4 ;
        RECT 70.155 178.825 70.485 179.155 ;
        RECT 50.835 171.345 51.165 171.675 ;
        RECT 50.850 166.915 51.150 171.345 ;
        RECT 50.835 166.585 51.165 166.915 ;
        RECT 50.850 155.355 51.150 166.585 ;
        RECT 70.170 155.355 70.470 178.825 ;
        RECT 50.835 155.025 51.165 155.355 ;
        RECT 57.275 155.025 57.605 155.355 ;
        RECT 70.155 155.025 70.485 155.355 ;
        RECT 57.290 124.755 57.590 155.025 ;
        RECT 57.275 124.425 57.605 124.755 ;
  END
END tt_um_08_sws
END LIBRARY

